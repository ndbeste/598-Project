module accbin2
    #( parameter bW = 8 )
    (
    input  logic [0:18*12*12*bW-1] i_accbin_in,
    input  logic [bW-1:0]          kernel_offset,
    output logic [0:8*8-1]         o_accbin_out
    );

logic [bW-1:0] sum_out         [0:11][0:11];
logic [bW-1:0] accbin_in  [0:4][0:11][0:11];
logic          accbin_out      [0: 7][0: 7];

genvar i,j,k;
for (i=0; i<12; i=i+1) begin
    for (j=0; j<12; j=j+1) begin
        for (k=0; k<18; k=k+1) begin
            assign accbin_in[i][j][k][l] = i_accbin_in[ 12*18*bW*i + 18*bW*j + bW*k : 12*18*bW*i + 18*bW*j + bW*k + 7];
        end
    end
end

for (i=0; i<12; i=i+1) begin
    for (j=0; j<12; j=j+1) begin
        assign o_accbin_out[ i*12 + j ] = accbin_out[i][j];
    end
end
assign sum_out[0][0][bW-1:0] = accbin_in[0][0][0][bW-1:0] + accbin_in[1][0][0][bW-1:0] + accbin_in[2][0][0][bW-1:0] + accbin_in[3][0][0][bW-1:0] + accbin_in[4][0][0][bW-1:0] + accbin_in[5][0][0][bW-1:0] + accbin_in[6][0][0][bW-1:0] + accbin_in[7][0][0][bW-1:0] + accbin_in[8][0][0][bW-1:0] + accbin_in[9][0][0][bW-1:0] + accbin_in[10][0][0][bW-1:0] + accbin_in[11][0][0][bW-1:0] + accbin_in[12][0][0][bW-1:0] + accbin_in[13][0][0][bW-1:0] + accbin_in[14][0][0][bW-1:0] + accbin_in[15][0][0][bW-1:0] + accbin_in[16][0][0][bW-1:0] + accbin_in[17][0][0][bW-1:0];
assign sum_out[0][1][bW-1:0] = accbin_in[0][0][1][bW-1:0] + accbin_in[1][0][1][bW-1:0] + accbin_in[2][0][1][bW-1:0] + accbin_in[3][0][1][bW-1:0] + accbin_in[4][0][1][bW-1:0] + accbin_in[5][0][1][bW-1:0] + accbin_in[6][0][1][bW-1:0] + accbin_in[7][0][1][bW-1:0] + accbin_in[8][0][1][bW-1:0] + accbin_in[9][0][1][bW-1:0] + accbin_in[10][0][1][bW-1:0] + accbin_in[11][0][1][bW-1:0] + accbin_in[12][0][1][bW-1:0] + accbin_in[13][0][1][bW-1:0] + accbin_in[14][0][1][bW-1:0] + accbin_in[15][0][1][bW-1:0] + accbin_in[16][0][1][bW-1:0] + accbin_in[17][0][1][bW-1:0];
assign sum_out[0][2][bW-1:0] = accbin_in[0][0][2][bW-1:0] + accbin_in[1][0][2][bW-1:0] + accbin_in[2][0][2][bW-1:0] + accbin_in[3][0][2][bW-1:0] + accbin_in[4][0][2][bW-1:0] + accbin_in[5][0][2][bW-1:0] + accbin_in[6][0][2][bW-1:0] + accbin_in[7][0][2][bW-1:0] + accbin_in[8][0][2][bW-1:0] + accbin_in[9][0][2][bW-1:0] + accbin_in[10][0][2][bW-1:0] + accbin_in[11][0][2][bW-1:0] + accbin_in[12][0][2][bW-1:0] + accbin_in[13][0][2][bW-1:0] + accbin_in[14][0][2][bW-1:0] + accbin_in[15][0][2][bW-1:0] + accbin_in[16][0][2][bW-1:0] + accbin_in[17][0][2][bW-1:0];
assign sum_out[0][3][bW-1:0] = accbin_in[0][0][3][bW-1:0] + accbin_in[1][0][3][bW-1:0] + accbin_in[2][0][3][bW-1:0] + accbin_in[3][0][3][bW-1:0] + accbin_in[4][0][3][bW-1:0] + accbin_in[5][0][3][bW-1:0] + accbin_in[6][0][3][bW-1:0] + accbin_in[7][0][3][bW-1:0] + accbin_in[8][0][3][bW-1:0] + accbin_in[9][0][3][bW-1:0] + accbin_in[10][0][3][bW-1:0] + accbin_in[11][0][3][bW-1:0] + accbin_in[12][0][3][bW-1:0] + accbin_in[13][0][3][bW-1:0] + accbin_in[14][0][3][bW-1:0] + accbin_in[15][0][3][bW-1:0] + accbin_in[16][0][3][bW-1:0] + accbin_in[17][0][3][bW-1:0];
assign sum_out[0][4][bW-1:0] = accbin_in[0][0][4][bW-1:0] + accbin_in[1][0][4][bW-1:0] + accbin_in[2][0][4][bW-1:0] + accbin_in[3][0][4][bW-1:0] + accbin_in[4][0][4][bW-1:0] + accbin_in[5][0][4][bW-1:0] + accbin_in[6][0][4][bW-1:0] + accbin_in[7][0][4][bW-1:0] + accbin_in[8][0][4][bW-1:0] + accbin_in[9][0][4][bW-1:0] + accbin_in[10][0][4][bW-1:0] + accbin_in[11][0][4][bW-1:0] + accbin_in[12][0][4][bW-1:0] + accbin_in[13][0][4][bW-1:0] + accbin_in[14][0][4][bW-1:0] + accbin_in[15][0][4][bW-1:0] + accbin_in[16][0][4][bW-1:0] + accbin_in[17][0][4][bW-1:0];
assign sum_out[0][5][bW-1:0] = accbin_in[0][0][5][bW-1:0] + accbin_in[1][0][5][bW-1:0] + accbin_in[2][0][5][bW-1:0] + accbin_in[3][0][5][bW-1:0] + accbin_in[4][0][5][bW-1:0] + accbin_in[5][0][5][bW-1:0] + accbin_in[6][0][5][bW-1:0] + accbin_in[7][0][5][bW-1:0] + accbin_in[8][0][5][bW-1:0] + accbin_in[9][0][5][bW-1:0] + accbin_in[10][0][5][bW-1:0] + accbin_in[11][0][5][bW-1:0] + accbin_in[12][0][5][bW-1:0] + accbin_in[13][0][5][bW-1:0] + accbin_in[14][0][5][bW-1:0] + accbin_in[15][0][5][bW-1:0] + accbin_in[16][0][5][bW-1:0] + accbin_in[17][0][5][bW-1:0];
assign sum_out[0][6][bW-1:0] = accbin_in[0][0][6][bW-1:0] + accbin_in[1][0][6][bW-1:0] + accbin_in[2][0][6][bW-1:0] + accbin_in[3][0][6][bW-1:0] + accbin_in[4][0][6][bW-1:0] + accbin_in[5][0][6][bW-1:0] + accbin_in[6][0][6][bW-1:0] + accbin_in[7][0][6][bW-1:0] + accbin_in[8][0][6][bW-1:0] + accbin_in[9][0][6][bW-1:0] + accbin_in[10][0][6][bW-1:0] + accbin_in[11][0][6][bW-1:0] + accbin_in[12][0][6][bW-1:0] + accbin_in[13][0][6][bW-1:0] + accbin_in[14][0][6][bW-1:0] + accbin_in[15][0][6][bW-1:0] + accbin_in[16][0][6][bW-1:0] + accbin_in[17][0][6][bW-1:0];
assign sum_out[0][7][bW-1:0] = accbin_in[0][0][7][bW-1:0] + accbin_in[1][0][7][bW-1:0] + accbin_in[2][0][7][bW-1:0] + accbin_in[3][0][7][bW-1:0] + accbin_in[4][0][7][bW-1:0] + accbin_in[5][0][7][bW-1:0] + accbin_in[6][0][7][bW-1:0] + accbin_in[7][0][7][bW-1:0] + accbin_in[8][0][7][bW-1:0] + accbin_in[9][0][7][bW-1:0] + accbin_in[10][0][7][bW-1:0] + accbin_in[11][0][7][bW-1:0] + accbin_in[12][0][7][bW-1:0] + accbin_in[13][0][7][bW-1:0] + accbin_in[14][0][7][bW-1:0] + accbin_in[15][0][7][bW-1:0] + accbin_in[16][0][7][bW-1:0] + accbin_in[17][0][7][bW-1:0];
assign sum_out[0][8][bW-1:0] = accbin_in[0][0][8][bW-1:0] + accbin_in[1][0][8][bW-1:0] + accbin_in[2][0][8][bW-1:0] + accbin_in[3][0][8][bW-1:0] + accbin_in[4][0][8][bW-1:0] + accbin_in[5][0][8][bW-1:0] + accbin_in[6][0][8][bW-1:0] + accbin_in[7][0][8][bW-1:0] + accbin_in[8][0][8][bW-1:0] + accbin_in[9][0][8][bW-1:0] + accbin_in[10][0][8][bW-1:0] + accbin_in[11][0][8][bW-1:0] + accbin_in[12][0][8][bW-1:0] + accbin_in[13][0][8][bW-1:0] + accbin_in[14][0][8][bW-1:0] + accbin_in[15][0][8][bW-1:0] + accbin_in[16][0][8][bW-1:0] + accbin_in[17][0][8][bW-1:0];
assign sum_out[0][9][bW-1:0] = accbin_in[0][0][9][bW-1:0] + accbin_in[1][0][9][bW-1:0] + accbin_in[2][0][9][bW-1:0] + accbin_in[3][0][9][bW-1:0] + accbin_in[4][0][9][bW-1:0] + accbin_in[5][0][9][bW-1:0] + accbin_in[6][0][9][bW-1:0] + accbin_in[7][0][9][bW-1:0] + accbin_in[8][0][9][bW-1:0] + accbin_in[9][0][9][bW-1:0] + accbin_in[10][0][9][bW-1:0] + accbin_in[11][0][9][bW-1:0] + accbin_in[12][0][9][bW-1:0] + accbin_in[13][0][9][bW-1:0] + accbin_in[14][0][9][bW-1:0] + accbin_in[15][0][9][bW-1:0] + accbin_in[16][0][9][bW-1:0] + accbin_in[17][0][9][bW-1:0];
assign sum_out[0][10][bW-1:0] = accbin_in[0][0][10][bW-1:0] + accbin_in[1][0][10][bW-1:0] + accbin_in[2][0][10][bW-1:0] + accbin_in[3][0][10][bW-1:0] + accbin_in[4][0][10][bW-1:0] + accbin_in[5][0][10][bW-1:0] + accbin_in[6][0][10][bW-1:0] + accbin_in[7][0][10][bW-1:0] + accbin_in[8][0][10][bW-1:0] + accbin_in[9][0][10][bW-1:0] + accbin_in[10][0][10][bW-1:0] + accbin_in[11][0][10][bW-1:0] + accbin_in[12][0][10][bW-1:0] + accbin_in[13][0][10][bW-1:0] + accbin_in[14][0][10][bW-1:0] + accbin_in[15][0][10][bW-1:0] + accbin_in[16][0][10][bW-1:0] + accbin_in[17][0][10][bW-1:0];
assign sum_out[0][11][bW-1:0] = accbin_in[0][0][11][bW-1:0] + accbin_in[1][0][11][bW-1:0] + accbin_in[2][0][11][bW-1:0] + accbin_in[3][0][11][bW-1:0] + accbin_in[4][0][11][bW-1:0] + accbin_in[5][0][11][bW-1:0] + accbin_in[6][0][11][bW-1:0] + accbin_in[7][0][11][bW-1:0] + accbin_in[8][0][11][bW-1:0] + accbin_in[9][0][11][bW-1:0] + accbin_in[10][0][11][bW-1:0] + accbin_in[11][0][11][bW-1:0] + accbin_in[12][0][11][bW-1:0] + accbin_in[13][0][11][bW-1:0] + accbin_in[14][0][11][bW-1:0] + accbin_in[15][0][11][bW-1:0] + accbin_in[16][0][11][bW-1:0] + accbin_in[17][0][11][bW-1:0];
assign sum_out[1][0][bW-1:0] = accbin_in[0][1][0][bW-1:0] + accbin_in[1][1][0][bW-1:0] + accbin_in[2][1][0][bW-1:0] + accbin_in[3][1][0][bW-1:0] + accbin_in[4][1][0][bW-1:0] + accbin_in[5][1][0][bW-1:0] + accbin_in[6][1][0][bW-1:0] + accbin_in[7][1][0][bW-1:0] + accbin_in[8][1][0][bW-1:0] + accbin_in[9][1][0][bW-1:0] + accbin_in[10][1][0][bW-1:0] + accbin_in[11][1][0][bW-1:0] + accbin_in[12][1][0][bW-1:0] + accbin_in[13][1][0][bW-1:0] + accbin_in[14][1][0][bW-1:0] + accbin_in[15][1][0][bW-1:0] + accbin_in[16][1][0][bW-1:0] + accbin_in[17][1][0][bW-1:0];
assign sum_out[1][1][bW-1:0] = accbin_in[0][1][1][bW-1:0] + accbin_in[1][1][1][bW-1:0] + accbin_in[2][1][1][bW-1:0] + accbin_in[3][1][1][bW-1:0] + accbin_in[4][1][1][bW-1:0] + accbin_in[5][1][1][bW-1:0] + accbin_in[6][1][1][bW-1:0] + accbin_in[7][1][1][bW-1:0] + accbin_in[8][1][1][bW-1:0] + accbin_in[9][1][1][bW-1:0] + accbin_in[10][1][1][bW-1:0] + accbin_in[11][1][1][bW-1:0] + accbin_in[12][1][1][bW-1:0] + accbin_in[13][1][1][bW-1:0] + accbin_in[14][1][1][bW-1:0] + accbin_in[15][1][1][bW-1:0] + accbin_in[16][1][1][bW-1:0] + accbin_in[17][1][1][bW-1:0];
assign sum_out[1][2][bW-1:0] = accbin_in[0][1][2][bW-1:0] + accbin_in[1][1][2][bW-1:0] + accbin_in[2][1][2][bW-1:0] + accbin_in[3][1][2][bW-1:0] + accbin_in[4][1][2][bW-1:0] + accbin_in[5][1][2][bW-1:0] + accbin_in[6][1][2][bW-1:0] + accbin_in[7][1][2][bW-1:0] + accbin_in[8][1][2][bW-1:0] + accbin_in[9][1][2][bW-1:0] + accbin_in[10][1][2][bW-1:0] + accbin_in[11][1][2][bW-1:0] + accbin_in[12][1][2][bW-1:0] + accbin_in[13][1][2][bW-1:0] + accbin_in[14][1][2][bW-1:0] + accbin_in[15][1][2][bW-1:0] + accbin_in[16][1][2][bW-1:0] + accbin_in[17][1][2][bW-1:0];
assign sum_out[1][3][bW-1:0] = accbin_in[0][1][3][bW-1:0] + accbin_in[1][1][3][bW-1:0] + accbin_in[2][1][3][bW-1:0] + accbin_in[3][1][3][bW-1:0] + accbin_in[4][1][3][bW-1:0] + accbin_in[5][1][3][bW-1:0] + accbin_in[6][1][3][bW-1:0] + accbin_in[7][1][3][bW-1:0] + accbin_in[8][1][3][bW-1:0] + accbin_in[9][1][3][bW-1:0] + accbin_in[10][1][3][bW-1:0] + accbin_in[11][1][3][bW-1:0] + accbin_in[12][1][3][bW-1:0] + accbin_in[13][1][3][bW-1:0] + accbin_in[14][1][3][bW-1:0] + accbin_in[15][1][3][bW-1:0] + accbin_in[16][1][3][bW-1:0] + accbin_in[17][1][3][bW-1:0];
assign sum_out[1][4][bW-1:0] = accbin_in[0][1][4][bW-1:0] + accbin_in[1][1][4][bW-1:0] + accbin_in[2][1][4][bW-1:0] + accbin_in[3][1][4][bW-1:0] + accbin_in[4][1][4][bW-1:0] + accbin_in[5][1][4][bW-1:0] + accbin_in[6][1][4][bW-1:0] + accbin_in[7][1][4][bW-1:0] + accbin_in[8][1][4][bW-1:0] + accbin_in[9][1][4][bW-1:0] + accbin_in[10][1][4][bW-1:0] + accbin_in[11][1][4][bW-1:0] + accbin_in[12][1][4][bW-1:0] + accbin_in[13][1][4][bW-1:0] + accbin_in[14][1][4][bW-1:0] + accbin_in[15][1][4][bW-1:0] + accbin_in[16][1][4][bW-1:0] + accbin_in[17][1][4][bW-1:0];
assign sum_out[1][5][bW-1:0] = accbin_in[0][1][5][bW-1:0] + accbin_in[1][1][5][bW-1:0] + accbin_in[2][1][5][bW-1:0] + accbin_in[3][1][5][bW-1:0] + accbin_in[4][1][5][bW-1:0] + accbin_in[5][1][5][bW-1:0] + accbin_in[6][1][5][bW-1:0] + accbin_in[7][1][5][bW-1:0] + accbin_in[8][1][5][bW-1:0] + accbin_in[9][1][5][bW-1:0] + accbin_in[10][1][5][bW-1:0] + accbin_in[11][1][5][bW-1:0] + accbin_in[12][1][5][bW-1:0] + accbin_in[13][1][5][bW-1:0] + accbin_in[14][1][5][bW-1:0] + accbin_in[15][1][5][bW-1:0] + accbin_in[16][1][5][bW-1:0] + accbin_in[17][1][5][bW-1:0];
assign sum_out[1][6][bW-1:0] = accbin_in[0][1][6][bW-1:0] + accbin_in[1][1][6][bW-1:0] + accbin_in[2][1][6][bW-1:0] + accbin_in[3][1][6][bW-1:0] + accbin_in[4][1][6][bW-1:0] + accbin_in[5][1][6][bW-1:0] + accbin_in[6][1][6][bW-1:0] + accbin_in[7][1][6][bW-1:0] + accbin_in[8][1][6][bW-1:0] + accbin_in[9][1][6][bW-1:0] + accbin_in[10][1][6][bW-1:0] + accbin_in[11][1][6][bW-1:0] + accbin_in[12][1][6][bW-1:0] + accbin_in[13][1][6][bW-1:0] + accbin_in[14][1][6][bW-1:0] + accbin_in[15][1][6][bW-1:0] + accbin_in[16][1][6][bW-1:0] + accbin_in[17][1][6][bW-1:0];
assign sum_out[1][7][bW-1:0] = accbin_in[0][1][7][bW-1:0] + accbin_in[1][1][7][bW-1:0] + accbin_in[2][1][7][bW-1:0] + accbin_in[3][1][7][bW-1:0] + accbin_in[4][1][7][bW-1:0] + accbin_in[5][1][7][bW-1:0] + accbin_in[6][1][7][bW-1:0] + accbin_in[7][1][7][bW-1:0] + accbin_in[8][1][7][bW-1:0] + accbin_in[9][1][7][bW-1:0] + accbin_in[10][1][7][bW-1:0] + accbin_in[11][1][7][bW-1:0] + accbin_in[12][1][7][bW-1:0] + accbin_in[13][1][7][bW-1:0] + accbin_in[14][1][7][bW-1:0] + accbin_in[15][1][7][bW-1:0] + accbin_in[16][1][7][bW-1:0] + accbin_in[17][1][7][bW-1:0];
assign sum_out[1][8][bW-1:0] = accbin_in[0][1][8][bW-1:0] + accbin_in[1][1][8][bW-1:0] + accbin_in[2][1][8][bW-1:0] + accbin_in[3][1][8][bW-1:0] + accbin_in[4][1][8][bW-1:0] + accbin_in[5][1][8][bW-1:0] + accbin_in[6][1][8][bW-1:0] + accbin_in[7][1][8][bW-1:0] + accbin_in[8][1][8][bW-1:0] + accbin_in[9][1][8][bW-1:0] + accbin_in[10][1][8][bW-1:0] + accbin_in[11][1][8][bW-1:0] + accbin_in[12][1][8][bW-1:0] + accbin_in[13][1][8][bW-1:0] + accbin_in[14][1][8][bW-1:0] + accbin_in[15][1][8][bW-1:0] + accbin_in[16][1][8][bW-1:0] + accbin_in[17][1][8][bW-1:0];
assign sum_out[1][9][bW-1:0] = accbin_in[0][1][9][bW-1:0] + accbin_in[1][1][9][bW-1:0] + accbin_in[2][1][9][bW-1:0] + accbin_in[3][1][9][bW-1:0] + accbin_in[4][1][9][bW-1:0] + accbin_in[5][1][9][bW-1:0] + accbin_in[6][1][9][bW-1:0] + accbin_in[7][1][9][bW-1:0] + accbin_in[8][1][9][bW-1:0] + accbin_in[9][1][9][bW-1:0] + accbin_in[10][1][9][bW-1:0] + accbin_in[11][1][9][bW-1:0] + accbin_in[12][1][9][bW-1:0] + accbin_in[13][1][9][bW-1:0] + accbin_in[14][1][9][bW-1:0] + accbin_in[15][1][9][bW-1:0] + accbin_in[16][1][9][bW-1:0] + accbin_in[17][1][9][bW-1:0];
assign sum_out[1][10][bW-1:0] = accbin_in[0][1][10][bW-1:0] + accbin_in[1][1][10][bW-1:0] + accbin_in[2][1][10][bW-1:0] + accbin_in[3][1][10][bW-1:0] + accbin_in[4][1][10][bW-1:0] + accbin_in[5][1][10][bW-1:0] + accbin_in[6][1][10][bW-1:0] + accbin_in[7][1][10][bW-1:0] + accbin_in[8][1][10][bW-1:0] + accbin_in[9][1][10][bW-1:0] + accbin_in[10][1][10][bW-1:0] + accbin_in[11][1][10][bW-1:0] + accbin_in[12][1][10][bW-1:0] + accbin_in[13][1][10][bW-1:0] + accbin_in[14][1][10][bW-1:0] + accbin_in[15][1][10][bW-1:0] + accbin_in[16][1][10][bW-1:0] + accbin_in[17][1][10][bW-1:0];
assign sum_out[1][11][bW-1:0] = accbin_in[0][1][11][bW-1:0] + accbin_in[1][1][11][bW-1:0] + accbin_in[2][1][11][bW-1:0] + accbin_in[3][1][11][bW-1:0] + accbin_in[4][1][11][bW-1:0] + accbin_in[5][1][11][bW-1:0] + accbin_in[6][1][11][bW-1:0] + accbin_in[7][1][11][bW-1:0] + accbin_in[8][1][11][bW-1:0] + accbin_in[9][1][11][bW-1:0] + accbin_in[10][1][11][bW-1:0] + accbin_in[11][1][11][bW-1:0] + accbin_in[12][1][11][bW-1:0] + accbin_in[13][1][11][bW-1:0] + accbin_in[14][1][11][bW-1:0] + accbin_in[15][1][11][bW-1:0] + accbin_in[16][1][11][bW-1:0] + accbin_in[17][1][11][bW-1:0];
assign sum_out[2][0][bW-1:0] = accbin_in[0][2][0][bW-1:0] + accbin_in[1][2][0][bW-1:0] + accbin_in[2][2][0][bW-1:0] + accbin_in[3][2][0][bW-1:0] + accbin_in[4][2][0][bW-1:0] + accbin_in[5][2][0][bW-1:0] + accbin_in[6][2][0][bW-1:0] + accbin_in[7][2][0][bW-1:0] + accbin_in[8][2][0][bW-1:0] + accbin_in[9][2][0][bW-1:0] + accbin_in[10][2][0][bW-1:0] + accbin_in[11][2][0][bW-1:0] + accbin_in[12][2][0][bW-1:0] + accbin_in[13][2][0][bW-1:0] + accbin_in[14][2][0][bW-1:0] + accbin_in[15][2][0][bW-1:0] + accbin_in[16][2][0][bW-1:0] + accbin_in[17][2][0][bW-1:0];
assign sum_out[2][1][bW-1:0] = accbin_in[0][2][1][bW-1:0] + accbin_in[1][2][1][bW-1:0] + accbin_in[2][2][1][bW-1:0] + accbin_in[3][2][1][bW-1:0] + accbin_in[4][2][1][bW-1:0] + accbin_in[5][2][1][bW-1:0] + accbin_in[6][2][1][bW-1:0] + accbin_in[7][2][1][bW-1:0] + accbin_in[8][2][1][bW-1:0] + accbin_in[9][2][1][bW-1:0] + accbin_in[10][2][1][bW-1:0] + accbin_in[11][2][1][bW-1:0] + accbin_in[12][2][1][bW-1:0] + accbin_in[13][2][1][bW-1:0] + accbin_in[14][2][1][bW-1:0] + accbin_in[15][2][1][bW-1:0] + accbin_in[16][2][1][bW-1:0] + accbin_in[17][2][1][bW-1:0];
assign sum_out[2][2][bW-1:0] = accbin_in[0][2][2][bW-1:0] + accbin_in[1][2][2][bW-1:0] + accbin_in[2][2][2][bW-1:0] + accbin_in[3][2][2][bW-1:0] + accbin_in[4][2][2][bW-1:0] + accbin_in[5][2][2][bW-1:0] + accbin_in[6][2][2][bW-1:0] + accbin_in[7][2][2][bW-1:0] + accbin_in[8][2][2][bW-1:0] + accbin_in[9][2][2][bW-1:0] + accbin_in[10][2][2][bW-1:0] + accbin_in[11][2][2][bW-1:0] + accbin_in[12][2][2][bW-1:0] + accbin_in[13][2][2][bW-1:0] + accbin_in[14][2][2][bW-1:0] + accbin_in[15][2][2][bW-1:0] + accbin_in[16][2][2][bW-1:0] + accbin_in[17][2][2][bW-1:0];
assign sum_out[2][3][bW-1:0] = accbin_in[0][2][3][bW-1:0] + accbin_in[1][2][3][bW-1:0] + accbin_in[2][2][3][bW-1:0] + accbin_in[3][2][3][bW-1:0] + accbin_in[4][2][3][bW-1:0] + accbin_in[5][2][3][bW-1:0] + accbin_in[6][2][3][bW-1:0] + accbin_in[7][2][3][bW-1:0] + accbin_in[8][2][3][bW-1:0] + accbin_in[9][2][3][bW-1:0] + accbin_in[10][2][3][bW-1:0] + accbin_in[11][2][3][bW-1:0] + accbin_in[12][2][3][bW-1:0] + accbin_in[13][2][3][bW-1:0] + accbin_in[14][2][3][bW-1:0] + accbin_in[15][2][3][bW-1:0] + accbin_in[16][2][3][bW-1:0] + accbin_in[17][2][3][bW-1:0];
assign sum_out[2][4][bW-1:0] = accbin_in[0][2][4][bW-1:0] + accbin_in[1][2][4][bW-1:0] + accbin_in[2][2][4][bW-1:0] + accbin_in[3][2][4][bW-1:0] + accbin_in[4][2][4][bW-1:0] + accbin_in[5][2][4][bW-1:0] + accbin_in[6][2][4][bW-1:0] + accbin_in[7][2][4][bW-1:0] + accbin_in[8][2][4][bW-1:0] + accbin_in[9][2][4][bW-1:0] + accbin_in[10][2][4][bW-1:0] + accbin_in[11][2][4][bW-1:0] + accbin_in[12][2][4][bW-1:0] + accbin_in[13][2][4][bW-1:0] + accbin_in[14][2][4][bW-1:0] + accbin_in[15][2][4][bW-1:0] + accbin_in[16][2][4][bW-1:0] + accbin_in[17][2][4][bW-1:0];
assign sum_out[2][5][bW-1:0] = accbin_in[0][2][5][bW-1:0] + accbin_in[1][2][5][bW-1:0] + accbin_in[2][2][5][bW-1:0] + accbin_in[3][2][5][bW-1:0] + accbin_in[4][2][5][bW-1:0] + accbin_in[5][2][5][bW-1:0] + accbin_in[6][2][5][bW-1:0] + accbin_in[7][2][5][bW-1:0] + accbin_in[8][2][5][bW-1:0] + accbin_in[9][2][5][bW-1:0] + accbin_in[10][2][5][bW-1:0] + accbin_in[11][2][5][bW-1:0] + accbin_in[12][2][5][bW-1:0] + accbin_in[13][2][5][bW-1:0] + accbin_in[14][2][5][bW-1:0] + accbin_in[15][2][5][bW-1:0] + accbin_in[16][2][5][bW-1:0] + accbin_in[17][2][5][bW-1:0];
assign sum_out[2][6][bW-1:0] = accbin_in[0][2][6][bW-1:0] + accbin_in[1][2][6][bW-1:0] + accbin_in[2][2][6][bW-1:0] + accbin_in[3][2][6][bW-1:0] + accbin_in[4][2][6][bW-1:0] + accbin_in[5][2][6][bW-1:0] + accbin_in[6][2][6][bW-1:0] + accbin_in[7][2][6][bW-1:0] + accbin_in[8][2][6][bW-1:0] + accbin_in[9][2][6][bW-1:0] + accbin_in[10][2][6][bW-1:0] + accbin_in[11][2][6][bW-1:0] + accbin_in[12][2][6][bW-1:0] + accbin_in[13][2][6][bW-1:0] + accbin_in[14][2][6][bW-1:0] + accbin_in[15][2][6][bW-1:0] + accbin_in[16][2][6][bW-1:0] + accbin_in[17][2][6][bW-1:0];
assign sum_out[2][7][bW-1:0] = accbin_in[0][2][7][bW-1:0] + accbin_in[1][2][7][bW-1:0] + accbin_in[2][2][7][bW-1:0] + accbin_in[3][2][7][bW-1:0] + accbin_in[4][2][7][bW-1:0] + accbin_in[5][2][7][bW-1:0] + accbin_in[6][2][7][bW-1:0] + accbin_in[7][2][7][bW-1:0] + accbin_in[8][2][7][bW-1:0] + accbin_in[9][2][7][bW-1:0] + accbin_in[10][2][7][bW-1:0] + accbin_in[11][2][7][bW-1:0] + accbin_in[12][2][7][bW-1:0] + accbin_in[13][2][7][bW-1:0] + accbin_in[14][2][7][bW-1:0] + accbin_in[15][2][7][bW-1:0] + accbin_in[16][2][7][bW-1:0] + accbin_in[17][2][7][bW-1:0];
assign sum_out[2][8][bW-1:0] = accbin_in[0][2][8][bW-1:0] + accbin_in[1][2][8][bW-1:0] + accbin_in[2][2][8][bW-1:0] + accbin_in[3][2][8][bW-1:0] + accbin_in[4][2][8][bW-1:0] + accbin_in[5][2][8][bW-1:0] + accbin_in[6][2][8][bW-1:0] + accbin_in[7][2][8][bW-1:0] + accbin_in[8][2][8][bW-1:0] + accbin_in[9][2][8][bW-1:0] + accbin_in[10][2][8][bW-1:0] + accbin_in[11][2][8][bW-1:0] + accbin_in[12][2][8][bW-1:0] + accbin_in[13][2][8][bW-1:0] + accbin_in[14][2][8][bW-1:0] + accbin_in[15][2][8][bW-1:0] + accbin_in[16][2][8][bW-1:0] + accbin_in[17][2][8][bW-1:0];
assign sum_out[2][9][bW-1:0] = accbin_in[0][2][9][bW-1:0] + accbin_in[1][2][9][bW-1:0] + accbin_in[2][2][9][bW-1:0] + accbin_in[3][2][9][bW-1:0] + accbin_in[4][2][9][bW-1:0] + accbin_in[5][2][9][bW-1:0] + accbin_in[6][2][9][bW-1:0] + accbin_in[7][2][9][bW-1:0] + accbin_in[8][2][9][bW-1:0] + accbin_in[9][2][9][bW-1:0] + accbin_in[10][2][9][bW-1:0] + accbin_in[11][2][9][bW-1:0] + accbin_in[12][2][9][bW-1:0] + accbin_in[13][2][9][bW-1:0] + accbin_in[14][2][9][bW-1:0] + accbin_in[15][2][9][bW-1:0] + accbin_in[16][2][9][bW-1:0] + accbin_in[17][2][9][bW-1:0];
assign sum_out[2][10][bW-1:0] = accbin_in[0][2][10][bW-1:0] + accbin_in[1][2][10][bW-1:0] + accbin_in[2][2][10][bW-1:0] + accbin_in[3][2][10][bW-1:0] + accbin_in[4][2][10][bW-1:0] + accbin_in[5][2][10][bW-1:0] + accbin_in[6][2][10][bW-1:0] + accbin_in[7][2][10][bW-1:0] + accbin_in[8][2][10][bW-1:0] + accbin_in[9][2][10][bW-1:0] + accbin_in[10][2][10][bW-1:0] + accbin_in[11][2][10][bW-1:0] + accbin_in[12][2][10][bW-1:0] + accbin_in[13][2][10][bW-1:0] + accbin_in[14][2][10][bW-1:0] + accbin_in[15][2][10][bW-1:0] + accbin_in[16][2][10][bW-1:0] + accbin_in[17][2][10][bW-1:0];
assign sum_out[2][11][bW-1:0] = accbin_in[0][2][11][bW-1:0] + accbin_in[1][2][11][bW-1:0] + accbin_in[2][2][11][bW-1:0] + accbin_in[3][2][11][bW-1:0] + accbin_in[4][2][11][bW-1:0] + accbin_in[5][2][11][bW-1:0] + accbin_in[6][2][11][bW-1:0] + accbin_in[7][2][11][bW-1:0] + accbin_in[8][2][11][bW-1:0] + accbin_in[9][2][11][bW-1:0] + accbin_in[10][2][11][bW-1:0] + accbin_in[11][2][11][bW-1:0] + accbin_in[12][2][11][bW-1:0] + accbin_in[13][2][11][bW-1:0] + accbin_in[14][2][11][bW-1:0] + accbin_in[15][2][11][bW-1:0] + accbin_in[16][2][11][bW-1:0] + accbin_in[17][2][11][bW-1:0];
assign sum_out[3][0][bW-1:0] = accbin_in[0][3][0][bW-1:0] + accbin_in[1][3][0][bW-1:0] + accbin_in[2][3][0][bW-1:0] + accbin_in[3][3][0][bW-1:0] + accbin_in[4][3][0][bW-1:0] + accbin_in[5][3][0][bW-1:0] + accbin_in[6][3][0][bW-1:0] + accbin_in[7][3][0][bW-1:0] + accbin_in[8][3][0][bW-1:0] + accbin_in[9][3][0][bW-1:0] + accbin_in[10][3][0][bW-1:0] + accbin_in[11][3][0][bW-1:0] + accbin_in[12][3][0][bW-1:0] + accbin_in[13][3][0][bW-1:0] + accbin_in[14][3][0][bW-1:0] + accbin_in[15][3][0][bW-1:0] + accbin_in[16][3][0][bW-1:0] + accbin_in[17][3][0][bW-1:0];
assign sum_out[3][1][bW-1:0] = accbin_in[0][3][1][bW-1:0] + accbin_in[1][3][1][bW-1:0] + accbin_in[2][3][1][bW-1:0] + accbin_in[3][3][1][bW-1:0] + accbin_in[4][3][1][bW-1:0] + accbin_in[5][3][1][bW-1:0] + accbin_in[6][3][1][bW-1:0] + accbin_in[7][3][1][bW-1:0] + accbin_in[8][3][1][bW-1:0] + accbin_in[9][3][1][bW-1:0] + accbin_in[10][3][1][bW-1:0] + accbin_in[11][3][1][bW-1:0] + accbin_in[12][3][1][bW-1:0] + accbin_in[13][3][1][bW-1:0] + accbin_in[14][3][1][bW-1:0] + accbin_in[15][3][1][bW-1:0] + accbin_in[16][3][1][bW-1:0] + accbin_in[17][3][1][bW-1:0];
assign sum_out[3][2][bW-1:0] = accbin_in[0][3][2][bW-1:0] + accbin_in[1][3][2][bW-1:0] + accbin_in[2][3][2][bW-1:0] + accbin_in[3][3][2][bW-1:0] + accbin_in[4][3][2][bW-1:0] + accbin_in[5][3][2][bW-1:0] + accbin_in[6][3][2][bW-1:0] + accbin_in[7][3][2][bW-1:0] + accbin_in[8][3][2][bW-1:0] + accbin_in[9][3][2][bW-1:0] + accbin_in[10][3][2][bW-1:0] + accbin_in[11][3][2][bW-1:0] + accbin_in[12][3][2][bW-1:0] + accbin_in[13][3][2][bW-1:0] + accbin_in[14][3][2][bW-1:0] + accbin_in[15][3][2][bW-1:0] + accbin_in[16][3][2][bW-1:0] + accbin_in[17][3][2][bW-1:0];
assign sum_out[3][3][bW-1:0] = accbin_in[0][3][3][bW-1:0] + accbin_in[1][3][3][bW-1:0] + accbin_in[2][3][3][bW-1:0] + accbin_in[3][3][3][bW-1:0] + accbin_in[4][3][3][bW-1:0] + accbin_in[5][3][3][bW-1:0] + accbin_in[6][3][3][bW-1:0] + accbin_in[7][3][3][bW-1:0] + accbin_in[8][3][3][bW-1:0] + accbin_in[9][3][3][bW-1:0] + accbin_in[10][3][3][bW-1:0] + accbin_in[11][3][3][bW-1:0] + accbin_in[12][3][3][bW-1:0] + accbin_in[13][3][3][bW-1:0] + accbin_in[14][3][3][bW-1:0] + accbin_in[15][3][3][bW-1:0] + accbin_in[16][3][3][bW-1:0] + accbin_in[17][3][3][bW-1:0];
assign sum_out[3][4][bW-1:0] = accbin_in[0][3][4][bW-1:0] + accbin_in[1][3][4][bW-1:0] + accbin_in[2][3][4][bW-1:0] + accbin_in[3][3][4][bW-1:0] + accbin_in[4][3][4][bW-1:0] + accbin_in[5][3][4][bW-1:0] + accbin_in[6][3][4][bW-1:0] + accbin_in[7][3][4][bW-1:0] + accbin_in[8][3][4][bW-1:0] + accbin_in[9][3][4][bW-1:0] + accbin_in[10][3][4][bW-1:0] + accbin_in[11][3][4][bW-1:0] + accbin_in[12][3][4][bW-1:0] + accbin_in[13][3][4][bW-1:0] + accbin_in[14][3][4][bW-1:0] + accbin_in[15][3][4][bW-1:0] + accbin_in[16][3][4][bW-1:0] + accbin_in[17][3][4][bW-1:0];
assign sum_out[3][5][bW-1:0] = accbin_in[0][3][5][bW-1:0] + accbin_in[1][3][5][bW-1:0] + accbin_in[2][3][5][bW-1:0] + accbin_in[3][3][5][bW-1:0] + accbin_in[4][3][5][bW-1:0] + accbin_in[5][3][5][bW-1:0] + accbin_in[6][3][5][bW-1:0] + accbin_in[7][3][5][bW-1:0] + accbin_in[8][3][5][bW-1:0] + accbin_in[9][3][5][bW-1:0] + accbin_in[10][3][5][bW-1:0] + accbin_in[11][3][5][bW-1:0] + accbin_in[12][3][5][bW-1:0] + accbin_in[13][3][5][bW-1:0] + accbin_in[14][3][5][bW-1:0] + accbin_in[15][3][5][bW-1:0] + accbin_in[16][3][5][bW-1:0] + accbin_in[17][3][5][bW-1:0];
assign sum_out[3][6][bW-1:0] = accbin_in[0][3][6][bW-1:0] + accbin_in[1][3][6][bW-1:0] + accbin_in[2][3][6][bW-1:0] + accbin_in[3][3][6][bW-1:0] + accbin_in[4][3][6][bW-1:0] + accbin_in[5][3][6][bW-1:0] + accbin_in[6][3][6][bW-1:0] + accbin_in[7][3][6][bW-1:0] + accbin_in[8][3][6][bW-1:0] + accbin_in[9][3][6][bW-1:0] + accbin_in[10][3][6][bW-1:0] + accbin_in[11][3][6][bW-1:0] + accbin_in[12][3][6][bW-1:0] + accbin_in[13][3][6][bW-1:0] + accbin_in[14][3][6][bW-1:0] + accbin_in[15][3][6][bW-1:0] + accbin_in[16][3][6][bW-1:0] + accbin_in[17][3][6][bW-1:0];
assign sum_out[3][7][bW-1:0] = accbin_in[0][3][7][bW-1:0] + accbin_in[1][3][7][bW-1:0] + accbin_in[2][3][7][bW-1:0] + accbin_in[3][3][7][bW-1:0] + accbin_in[4][3][7][bW-1:0] + accbin_in[5][3][7][bW-1:0] + accbin_in[6][3][7][bW-1:0] + accbin_in[7][3][7][bW-1:0] + accbin_in[8][3][7][bW-1:0] + accbin_in[9][3][7][bW-1:0] + accbin_in[10][3][7][bW-1:0] + accbin_in[11][3][7][bW-1:0] + accbin_in[12][3][7][bW-1:0] + accbin_in[13][3][7][bW-1:0] + accbin_in[14][3][7][bW-1:0] + accbin_in[15][3][7][bW-1:0] + accbin_in[16][3][7][bW-1:0] + accbin_in[17][3][7][bW-1:0];
assign sum_out[3][8][bW-1:0] = accbin_in[0][3][8][bW-1:0] + accbin_in[1][3][8][bW-1:0] + accbin_in[2][3][8][bW-1:0] + accbin_in[3][3][8][bW-1:0] + accbin_in[4][3][8][bW-1:0] + accbin_in[5][3][8][bW-1:0] + accbin_in[6][3][8][bW-1:0] + accbin_in[7][3][8][bW-1:0] + accbin_in[8][3][8][bW-1:0] + accbin_in[9][3][8][bW-1:0] + accbin_in[10][3][8][bW-1:0] + accbin_in[11][3][8][bW-1:0] + accbin_in[12][3][8][bW-1:0] + accbin_in[13][3][8][bW-1:0] + accbin_in[14][3][8][bW-1:0] + accbin_in[15][3][8][bW-1:0] + accbin_in[16][3][8][bW-1:0] + accbin_in[17][3][8][bW-1:0];
assign sum_out[3][9][bW-1:0] = accbin_in[0][3][9][bW-1:0] + accbin_in[1][3][9][bW-1:0] + accbin_in[2][3][9][bW-1:0] + accbin_in[3][3][9][bW-1:0] + accbin_in[4][3][9][bW-1:0] + accbin_in[5][3][9][bW-1:0] + accbin_in[6][3][9][bW-1:0] + accbin_in[7][3][9][bW-1:0] + accbin_in[8][3][9][bW-1:0] + accbin_in[9][3][9][bW-1:0] + accbin_in[10][3][9][bW-1:0] + accbin_in[11][3][9][bW-1:0] + accbin_in[12][3][9][bW-1:0] + accbin_in[13][3][9][bW-1:0] + accbin_in[14][3][9][bW-1:0] + accbin_in[15][3][9][bW-1:0] + accbin_in[16][3][9][bW-1:0] + accbin_in[17][3][9][bW-1:0];
assign sum_out[3][10][bW-1:0] = accbin_in[0][3][10][bW-1:0] + accbin_in[1][3][10][bW-1:0] + accbin_in[2][3][10][bW-1:0] + accbin_in[3][3][10][bW-1:0] + accbin_in[4][3][10][bW-1:0] + accbin_in[5][3][10][bW-1:0] + accbin_in[6][3][10][bW-1:0] + accbin_in[7][3][10][bW-1:0] + accbin_in[8][3][10][bW-1:0] + accbin_in[9][3][10][bW-1:0] + accbin_in[10][3][10][bW-1:0] + accbin_in[11][3][10][bW-1:0] + accbin_in[12][3][10][bW-1:0] + accbin_in[13][3][10][bW-1:0] + accbin_in[14][3][10][bW-1:0] + accbin_in[15][3][10][bW-1:0] + accbin_in[16][3][10][bW-1:0] + accbin_in[17][3][10][bW-1:0];
assign sum_out[3][11][bW-1:0] = accbin_in[0][3][11][bW-1:0] + accbin_in[1][3][11][bW-1:0] + accbin_in[2][3][11][bW-1:0] + accbin_in[3][3][11][bW-1:0] + accbin_in[4][3][11][bW-1:0] + accbin_in[5][3][11][bW-1:0] + accbin_in[6][3][11][bW-1:0] + accbin_in[7][3][11][bW-1:0] + accbin_in[8][3][11][bW-1:0] + accbin_in[9][3][11][bW-1:0] + accbin_in[10][3][11][bW-1:0] + accbin_in[11][3][11][bW-1:0] + accbin_in[12][3][11][bW-1:0] + accbin_in[13][3][11][bW-1:0] + accbin_in[14][3][11][bW-1:0] + accbin_in[15][3][11][bW-1:0] + accbin_in[16][3][11][bW-1:0] + accbin_in[17][3][11][bW-1:0];
assign sum_out[4][0][bW-1:0] = accbin_in[0][4][0][bW-1:0] + accbin_in[1][4][0][bW-1:0] + accbin_in[2][4][0][bW-1:0] + accbin_in[3][4][0][bW-1:0] + accbin_in[4][4][0][bW-1:0] + accbin_in[5][4][0][bW-1:0] + accbin_in[6][4][0][bW-1:0] + accbin_in[7][4][0][bW-1:0] + accbin_in[8][4][0][bW-1:0] + accbin_in[9][4][0][bW-1:0] + accbin_in[10][4][0][bW-1:0] + accbin_in[11][4][0][bW-1:0] + accbin_in[12][4][0][bW-1:0] + accbin_in[13][4][0][bW-1:0] + accbin_in[14][4][0][bW-1:0] + accbin_in[15][4][0][bW-1:0] + accbin_in[16][4][0][bW-1:0] + accbin_in[17][4][0][bW-1:0];
assign sum_out[4][1][bW-1:0] = accbin_in[0][4][1][bW-1:0] + accbin_in[1][4][1][bW-1:0] + accbin_in[2][4][1][bW-1:0] + accbin_in[3][4][1][bW-1:0] + accbin_in[4][4][1][bW-1:0] + accbin_in[5][4][1][bW-1:0] + accbin_in[6][4][1][bW-1:0] + accbin_in[7][4][1][bW-1:0] + accbin_in[8][4][1][bW-1:0] + accbin_in[9][4][1][bW-1:0] + accbin_in[10][4][1][bW-1:0] + accbin_in[11][4][1][bW-1:0] + accbin_in[12][4][1][bW-1:0] + accbin_in[13][4][1][bW-1:0] + accbin_in[14][4][1][bW-1:0] + accbin_in[15][4][1][bW-1:0] + accbin_in[16][4][1][bW-1:0] + accbin_in[17][4][1][bW-1:0];
assign sum_out[4][2][bW-1:0] = accbin_in[0][4][2][bW-1:0] + accbin_in[1][4][2][bW-1:0] + accbin_in[2][4][2][bW-1:0] + accbin_in[3][4][2][bW-1:0] + accbin_in[4][4][2][bW-1:0] + accbin_in[5][4][2][bW-1:0] + accbin_in[6][4][2][bW-1:0] + accbin_in[7][4][2][bW-1:0] + accbin_in[8][4][2][bW-1:0] + accbin_in[9][4][2][bW-1:0] + accbin_in[10][4][2][bW-1:0] + accbin_in[11][4][2][bW-1:0] + accbin_in[12][4][2][bW-1:0] + accbin_in[13][4][2][bW-1:0] + accbin_in[14][4][2][bW-1:0] + accbin_in[15][4][2][bW-1:0] + accbin_in[16][4][2][bW-1:0] + accbin_in[17][4][2][bW-1:0];
assign sum_out[4][3][bW-1:0] = accbin_in[0][4][3][bW-1:0] + accbin_in[1][4][3][bW-1:0] + accbin_in[2][4][3][bW-1:0] + accbin_in[3][4][3][bW-1:0] + accbin_in[4][4][3][bW-1:0] + accbin_in[5][4][3][bW-1:0] + accbin_in[6][4][3][bW-1:0] + accbin_in[7][4][3][bW-1:0] + accbin_in[8][4][3][bW-1:0] + accbin_in[9][4][3][bW-1:0] + accbin_in[10][4][3][bW-1:0] + accbin_in[11][4][3][bW-1:0] + accbin_in[12][4][3][bW-1:0] + accbin_in[13][4][3][bW-1:0] + accbin_in[14][4][3][bW-1:0] + accbin_in[15][4][3][bW-1:0] + accbin_in[16][4][3][bW-1:0] + accbin_in[17][4][3][bW-1:0];
assign sum_out[4][4][bW-1:0] = accbin_in[0][4][4][bW-1:0] + accbin_in[1][4][4][bW-1:0] + accbin_in[2][4][4][bW-1:0] + accbin_in[3][4][4][bW-1:0] + accbin_in[4][4][4][bW-1:0] + accbin_in[5][4][4][bW-1:0] + accbin_in[6][4][4][bW-1:0] + accbin_in[7][4][4][bW-1:0] + accbin_in[8][4][4][bW-1:0] + accbin_in[9][4][4][bW-1:0] + accbin_in[10][4][4][bW-1:0] + accbin_in[11][4][4][bW-1:0] + accbin_in[12][4][4][bW-1:0] + accbin_in[13][4][4][bW-1:0] + accbin_in[14][4][4][bW-1:0] + accbin_in[15][4][4][bW-1:0] + accbin_in[16][4][4][bW-1:0] + accbin_in[17][4][4][bW-1:0];
assign sum_out[4][5][bW-1:0] = accbin_in[0][4][5][bW-1:0] + accbin_in[1][4][5][bW-1:0] + accbin_in[2][4][5][bW-1:0] + accbin_in[3][4][5][bW-1:0] + accbin_in[4][4][5][bW-1:0] + accbin_in[5][4][5][bW-1:0] + accbin_in[6][4][5][bW-1:0] + accbin_in[7][4][5][bW-1:0] + accbin_in[8][4][5][bW-1:0] + accbin_in[9][4][5][bW-1:0] + accbin_in[10][4][5][bW-1:0] + accbin_in[11][4][5][bW-1:0] + accbin_in[12][4][5][bW-1:0] + accbin_in[13][4][5][bW-1:0] + accbin_in[14][4][5][bW-1:0] + accbin_in[15][4][5][bW-1:0] + accbin_in[16][4][5][bW-1:0] + accbin_in[17][4][5][bW-1:0];
assign sum_out[4][6][bW-1:0] = accbin_in[0][4][6][bW-1:0] + accbin_in[1][4][6][bW-1:0] + accbin_in[2][4][6][bW-1:0] + accbin_in[3][4][6][bW-1:0] + accbin_in[4][4][6][bW-1:0] + accbin_in[5][4][6][bW-1:0] + accbin_in[6][4][6][bW-1:0] + accbin_in[7][4][6][bW-1:0] + accbin_in[8][4][6][bW-1:0] + accbin_in[9][4][6][bW-1:0] + accbin_in[10][4][6][bW-1:0] + accbin_in[11][4][6][bW-1:0] + accbin_in[12][4][6][bW-1:0] + accbin_in[13][4][6][bW-1:0] + accbin_in[14][4][6][bW-1:0] + accbin_in[15][4][6][bW-1:0] + accbin_in[16][4][6][bW-1:0] + accbin_in[17][4][6][bW-1:0];
assign sum_out[4][7][bW-1:0] = accbin_in[0][4][7][bW-1:0] + accbin_in[1][4][7][bW-1:0] + accbin_in[2][4][7][bW-1:0] + accbin_in[3][4][7][bW-1:0] + accbin_in[4][4][7][bW-1:0] + accbin_in[5][4][7][bW-1:0] + accbin_in[6][4][7][bW-1:0] + accbin_in[7][4][7][bW-1:0] + accbin_in[8][4][7][bW-1:0] + accbin_in[9][4][7][bW-1:0] + accbin_in[10][4][7][bW-1:0] + accbin_in[11][4][7][bW-1:0] + accbin_in[12][4][7][bW-1:0] + accbin_in[13][4][7][bW-1:0] + accbin_in[14][4][7][bW-1:0] + accbin_in[15][4][7][bW-1:0] + accbin_in[16][4][7][bW-1:0] + accbin_in[17][4][7][bW-1:0];
assign sum_out[4][8][bW-1:0] = accbin_in[0][4][8][bW-1:0] + accbin_in[1][4][8][bW-1:0] + accbin_in[2][4][8][bW-1:0] + accbin_in[3][4][8][bW-1:0] + accbin_in[4][4][8][bW-1:0] + accbin_in[5][4][8][bW-1:0] + accbin_in[6][4][8][bW-1:0] + accbin_in[7][4][8][bW-1:0] + accbin_in[8][4][8][bW-1:0] + accbin_in[9][4][8][bW-1:0] + accbin_in[10][4][8][bW-1:0] + accbin_in[11][4][8][bW-1:0] + accbin_in[12][4][8][bW-1:0] + accbin_in[13][4][8][bW-1:0] + accbin_in[14][4][8][bW-1:0] + accbin_in[15][4][8][bW-1:0] + accbin_in[16][4][8][bW-1:0] + accbin_in[17][4][8][bW-1:0];
assign sum_out[4][9][bW-1:0] = accbin_in[0][4][9][bW-1:0] + accbin_in[1][4][9][bW-1:0] + accbin_in[2][4][9][bW-1:0] + accbin_in[3][4][9][bW-1:0] + accbin_in[4][4][9][bW-1:0] + accbin_in[5][4][9][bW-1:0] + accbin_in[6][4][9][bW-1:0] + accbin_in[7][4][9][bW-1:0] + accbin_in[8][4][9][bW-1:0] + accbin_in[9][4][9][bW-1:0] + accbin_in[10][4][9][bW-1:0] + accbin_in[11][4][9][bW-1:0] + accbin_in[12][4][9][bW-1:0] + accbin_in[13][4][9][bW-1:0] + accbin_in[14][4][9][bW-1:0] + accbin_in[15][4][9][bW-1:0] + accbin_in[16][4][9][bW-1:0] + accbin_in[17][4][9][bW-1:0];
assign sum_out[4][10][bW-1:0] = accbin_in[0][4][10][bW-1:0] + accbin_in[1][4][10][bW-1:0] + accbin_in[2][4][10][bW-1:0] + accbin_in[3][4][10][bW-1:0] + accbin_in[4][4][10][bW-1:0] + accbin_in[5][4][10][bW-1:0] + accbin_in[6][4][10][bW-1:0] + accbin_in[7][4][10][bW-1:0] + accbin_in[8][4][10][bW-1:0] + accbin_in[9][4][10][bW-1:0] + accbin_in[10][4][10][bW-1:0] + accbin_in[11][4][10][bW-1:0] + accbin_in[12][4][10][bW-1:0] + accbin_in[13][4][10][bW-1:0] + accbin_in[14][4][10][bW-1:0] + accbin_in[15][4][10][bW-1:0] + accbin_in[16][4][10][bW-1:0] + accbin_in[17][4][10][bW-1:0];
assign sum_out[4][11][bW-1:0] = accbin_in[0][4][11][bW-1:0] + accbin_in[1][4][11][bW-1:0] + accbin_in[2][4][11][bW-1:0] + accbin_in[3][4][11][bW-1:0] + accbin_in[4][4][11][bW-1:0] + accbin_in[5][4][11][bW-1:0] + accbin_in[6][4][11][bW-1:0] + accbin_in[7][4][11][bW-1:0] + accbin_in[8][4][11][bW-1:0] + accbin_in[9][4][11][bW-1:0] + accbin_in[10][4][11][bW-1:0] + accbin_in[11][4][11][bW-1:0] + accbin_in[12][4][11][bW-1:0] + accbin_in[13][4][11][bW-1:0] + accbin_in[14][4][11][bW-1:0] + accbin_in[15][4][11][bW-1:0] + accbin_in[16][4][11][bW-1:0] + accbin_in[17][4][11][bW-1:0];
assign sum_out[5][0][bW-1:0] = accbin_in[0][5][0][bW-1:0] + accbin_in[1][5][0][bW-1:0] + accbin_in[2][5][0][bW-1:0] + accbin_in[3][5][0][bW-1:0] + accbin_in[4][5][0][bW-1:0] + accbin_in[5][5][0][bW-1:0] + accbin_in[6][5][0][bW-1:0] + accbin_in[7][5][0][bW-1:0] + accbin_in[8][5][0][bW-1:0] + accbin_in[9][5][0][bW-1:0] + accbin_in[10][5][0][bW-1:0] + accbin_in[11][5][0][bW-1:0] + accbin_in[12][5][0][bW-1:0] + accbin_in[13][5][0][bW-1:0] + accbin_in[14][5][0][bW-1:0] + accbin_in[15][5][0][bW-1:0] + accbin_in[16][5][0][bW-1:0] + accbin_in[17][5][0][bW-1:0];
assign sum_out[5][1][bW-1:0] = accbin_in[0][5][1][bW-1:0] + accbin_in[1][5][1][bW-1:0] + accbin_in[2][5][1][bW-1:0] + accbin_in[3][5][1][bW-1:0] + accbin_in[4][5][1][bW-1:0] + accbin_in[5][5][1][bW-1:0] + accbin_in[6][5][1][bW-1:0] + accbin_in[7][5][1][bW-1:0] + accbin_in[8][5][1][bW-1:0] + accbin_in[9][5][1][bW-1:0] + accbin_in[10][5][1][bW-1:0] + accbin_in[11][5][1][bW-1:0] + accbin_in[12][5][1][bW-1:0] + accbin_in[13][5][1][bW-1:0] + accbin_in[14][5][1][bW-1:0] + accbin_in[15][5][1][bW-1:0] + accbin_in[16][5][1][bW-1:0] + accbin_in[17][5][1][bW-1:0];
assign sum_out[5][2][bW-1:0] = accbin_in[0][5][2][bW-1:0] + accbin_in[1][5][2][bW-1:0] + accbin_in[2][5][2][bW-1:0] + accbin_in[3][5][2][bW-1:0] + accbin_in[4][5][2][bW-1:0] + accbin_in[5][5][2][bW-1:0] + accbin_in[6][5][2][bW-1:0] + accbin_in[7][5][2][bW-1:0] + accbin_in[8][5][2][bW-1:0] + accbin_in[9][5][2][bW-1:0] + accbin_in[10][5][2][bW-1:0] + accbin_in[11][5][2][bW-1:0] + accbin_in[12][5][2][bW-1:0] + accbin_in[13][5][2][bW-1:0] + accbin_in[14][5][2][bW-1:0] + accbin_in[15][5][2][bW-1:0] + accbin_in[16][5][2][bW-1:0] + accbin_in[17][5][2][bW-1:0];
assign sum_out[5][3][bW-1:0] = accbin_in[0][5][3][bW-1:0] + accbin_in[1][5][3][bW-1:0] + accbin_in[2][5][3][bW-1:0] + accbin_in[3][5][3][bW-1:0] + accbin_in[4][5][3][bW-1:0] + accbin_in[5][5][3][bW-1:0] + accbin_in[6][5][3][bW-1:0] + accbin_in[7][5][3][bW-1:0] + accbin_in[8][5][3][bW-1:0] + accbin_in[9][5][3][bW-1:0] + accbin_in[10][5][3][bW-1:0] + accbin_in[11][5][3][bW-1:0] + accbin_in[12][5][3][bW-1:0] + accbin_in[13][5][3][bW-1:0] + accbin_in[14][5][3][bW-1:0] + accbin_in[15][5][3][bW-1:0] + accbin_in[16][5][3][bW-1:0] + accbin_in[17][5][3][bW-1:0];
assign sum_out[5][4][bW-1:0] = accbin_in[0][5][4][bW-1:0] + accbin_in[1][5][4][bW-1:0] + accbin_in[2][5][4][bW-1:0] + accbin_in[3][5][4][bW-1:0] + accbin_in[4][5][4][bW-1:0] + accbin_in[5][5][4][bW-1:0] + accbin_in[6][5][4][bW-1:0] + accbin_in[7][5][4][bW-1:0] + accbin_in[8][5][4][bW-1:0] + accbin_in[9][5][4][bW-1:0] + accbin_in[10][5][4][bW-1:0] + accbin_in[11][5][4][bW-1:0] + accbin_in[12][5][4][bW-1:0] + accbin_in[13][5][4][bW-1:0] + accbin_in[14][5][4][bW-1:0] + accbin_in[15][5][4][bW-1:0] + accbin_in[16][5][4][bW-1:0] + accbin_in[17][5][4][bW-1:0];
assign sum_out[5][5][bW-1:0] = accbin_in[0][5][5][bW-1:0] + accbin_in[1][5][5][bW-1:0] + accbin_in[2][5][5][bW-1:0] + accbin_in[3][5][5][bW-1:0] + accbin_in[4][5][5][bW-1:0] + accbin_in[5][5][5][bW-1:0] + accbin_in[6][5][5][bW-1:0] + accbin_in[7][5][5][bW-1:0] + accbin_in[8][5][5][bW-1:0] + accbin_in[9][5][5][bW-1:0] + accbin_in[10][5][5][bW-1:0] + accbin_in[11][5][5][bW-1:0] + accbin_in[12][5][5][bW-1:0] + accbin_in[13][5][5][bW-1:0] + accbin_in[14][5][5][bW-1:0] + accbin_in[15][5][5][bW-1:0] + accbin_in[16][5][5][bW-1:0] + accbin_in[17][5][5][bW-1:0];
assign sum_out[5][6][bW-1:0] = accbin_in[0][5][6][bW-1:0] + accbin_in[1][5][6][bW-1:0] + accbin_in[2][5][6][bW-1:0] + accbin_in[3][5][6][bW-1:0] + accbin_in[4][5][6][bW-1:0] + accbin_in[5][5][6][bW-1:0] + accbin_in[6][5][6][bW-1:0] + accbin_in[7][5][6][bW-1:0] + accbin_in[8][5][6][bW-1:0] + accbin_in[9][5][6][bW-1:0] + accbin_in[10][5][6][bW-1:0] + accbin_in[11][5][6][bW-1:0] + accbin_in[12][5][6][bW-1:0] + accbin_in[13][5][6][bW-1:0] + accbin_in[14][5][6][bW-1:0] + accbin_in[15][5][6][bW-1:0] + accbin_in[16][5][6][bW-1:0] + accbin_in[17][5][6][bW-1:0];
assign sum_out[5][7][bW-1:0] = accbin_in[0][5][7][bW-1:0] + accbin_in[1][5][7][bW-1:0] + accbin_in[2][5][7][bW-1:0] + accbin_in[3][5][7][bW-1:0] + accbin_in[4][5][7][bW-1:0] + accbin_in[5][5][7][bW-1:0] + accbin_in[6][5][7][bW-1:0] + accbin_in[7][5][7][bW-1:0] + accbin_in[8][5][7][bW-1:0] + accbin_in[9][5][7][bW-1:0] + accbin_in[10][5][7][bW-1:0] + accbin_in[11][5][7][bW-1:0] + accbin_in[12][5][7][bW-1:0] + accbin_in[13][5][7][bW-1:0] + accbin_in[14][5][7][bW-1:0] + accbin_in[15][5][7][bW-1:0] + accbin_in[16][5][7][bW-1:0] + accbin_in[17][5][7][bW-1:0];
assign sum_out[5][8][bW-1:0] = accbin_in[0][5][8][bW-1:0] + accbin_in[1][5][8][bW-1:0] + accbin_in[2][5][8][bW-1:0] + accbin_in[3][5][8][bW-1:0] + accbin_in[4][5][8][bW-1:0] + accbin_in[5][5][8][bW-1:0] + accbin_in[6][5][8][bW-1:0] + accbin_in[7][5][8][bW-1:0] + accbin_in[8][5][8][bW-1:0] + accbin_in[9][5][8][bW-1:0] + accbin_in[10][5][8][bW-1:0] + accbin_in[11][5][8][bW-1:0] + accbin_in[12][5][8][bW-1:0] + accbin_in[13][5][8][bW-1:0] + accbin_in[14][5][8][bW-1:0] + accbin_in[15][5][8][bW-1:0] + accbin_in[16][5][8][bW-1:0] + accbin_in[17][5][8][bW-1:0];
assign sum_out[5][9][bW-1:0] = accbin_in[0][5][9][bW-1:0] + accbin_in[1][5][9][bW-1:0] + accbin_in[2][5][9][bW-1:0] + accbin_in[3][5][9][bW-1:0] + accbin_in[4][5][9][bW-1:0] + accbin_in[5][5][9][bW-1:0] + accbin_in[6][5][9][bW-1:0] + accbin_in[7][5][9][bW-1:0] + accbin_in[8][5][9][bW-1:0] + accbin_in[9][5][9][bW-1:0] + accbin_in[10][5][9][bW-1:0] + accbin_in[11][5][9][bW-1:0] + accbin_in[12][5][9][bW-1:0] + accbin_in[13][5][9][bW-1:0] + accbin_in[14][5][9][bW-1:0] + accbin_in[15][5][9][bW-1:0] + accbin_in[16][5][9][bW-1:0] + accbin_in[17][5][9][bW-1:0];
assign sum_out[5][10][bW-1:0] = accbin_in[0][5][10][bW-1:0] + accbin_in[1][5][10][bW-1:0] + accbin_in[2][5][10][bW-1:0] + accbin_in[3][5][10][bW-1:0] + accbin_in[4][5][10][bW-1:0] + accbin_in[5][5][10][bW-1:0] + accbin_in[6][5][10][bW-1:0] + accbin_in[7][5][10][bW-1:0] + accbin_in[8][5][10][bW-1:0] + accbin_in[9][5][10][bW-1:0] + accbin_in[10][5][10][bW-1:0] + accbin_in[11][5][10][bW-1:0] + accbin_in[12][5][10][bW-1:0] + accbin_in[13][5][10][bW-1:0] + accbin_in[14][5][10][bW-1:0] + accbin_in[15][5][10][bW-1:0] + accbin_in[16][5][10][bW-1:0] + accbin_in[17][5][10][bW-1:0];
assign sum_out[5][11][bW-1:0] = accbin_in[0][5][11][bW-1:0] + accbin_in[1][5][11][bW-1:0] + accbin_in[2][5][11][bW-1:0] + accbin_in[3][5][11][bW-1:0] + accbin_in[4][5][11][bW-1:0] + accbin_in[5][5][11][bW-1:0] + accbin_in[6][5][11][bW-1:0] + accbin_in[7][5][11][bW-1:0] + accbin_in[8][5][11][bW-1:0] + accbin_in[9][5][11][bW-1:0] + accbin_in[10][5][11][bW-1:0] + accbin_in[11][5][11][bW-1:0] + accbin_in[12][5][11][bW-1:0] + accbin_in[13][5][11][bW-1:0] + accbin_in[14][5][11][bW-1:0] + accbin_in[15][5][11][bW-1:0] + accbin_in[16][5][11][bW-1:0] + accbin_in[17][5][11][bW-1:0];
assign sum_out[6][0][bW-1:0] = accbin_in[0][6][0][bW-1:0] + accbin_in[1][6][0][bW-1:0] + accbin_in[2][6][0][bW-1:0] + accbin_in[3][6][0][bW-1:0] + accbin_in[4][6][0][bW-1:0] + accbin_in[5][6][0][bW-1:0] + accbin_in[6][6][0][bW-1:0] + accbin_in[7][6][0][bW-1:0] + accbin_in[8][6][0][bW-1:0] + accbin_in[9][6][0][bW-1:0] + accbin_in[10][6][0][bW-1:0] + accbin_in[11][6][0][bW-1:0] + accbin_in[12][6][0][bW-1:0] + accbin_in[13][6][0][bW-1:0] + accbin_in[14][6][0][bW-1:0] + accbin_in[15][6][0][bW-1:0] + accbin_in[16][6][0][bW-1:0] + accbin_in[17][6][0][bW-1:0];
assign sum_out[6][1][bW-1:0] = accbin_in[0][6][1][bW-1:0] + accbin_in[1][6][1][bW-1:0] + accbin_in[2][6][1][bW-1:0] + accbin_in[3][6][1][bW-1:0] + accbin_in[4][6][1][bW-1:0] + accbin_in[5][6][1][bW-1:0] + accbin_in[6][6][1][bW-1:0] + accbin_in[7][6][1][bW-1:0] + accbin_in[8][6][1][bW-1:0] + accbin_in[9][6][1][bW-1:0] + accbin_in[10][6][1][bW-1:0] + accbin_in[11][6][1][bW-1:0] + accbin_in[12][6][1][bW-1:0] + accbin_in[13][6][1][bW-1:0] + accbin_in[14][6][1][bW-1:0] + accbin_in[15][6][1][bW-1:0] + accbin_in[16][6][1][bW-1:0] + accbin_in[17][6][1][bW-1:0];
assign sum_out[6][2][bW-1:0] = accbin_in[0][6][2][bW-1:0] + accbin_in[1][6][2][bW-1:0] + accbin_in[2][6][2][bW-1:0] + accbin_in[3][6][2][bW-1:0] + accbin_in[4][6][2][bW-1:0] + accbin_in[5][6][2][bW-1:0] + accbin_in[6][6][2][bW-1:0] + accbin_in[7][6][2][bW-1:0] + accbin_in[8][6][2][bW-1:0] + accbin_in[9][6][2][bW-1:0] + accbin_in[10][6][2][bW-1:0] + accbin_in[11][6][2][bW-1:0] + accbin_in[12][6][2][bW-1:0] + accbin_in[13][6][2][bW-1:0] + accbin_in[14][6][2][bW-1:0] + accbin_in[15][6][2][bW-1:0] + accbin_in[16][6][2][bW-1:0] + accbin_in[17][6][2][bW-1:0];
assign sum_out[6][3][bW-1:0] = accbin_in[0][6][3][bW-1:0] + accbin_in[1][6][3][bW-1:0] + accbin_in[2][6][3][bW-1:0] + accbin_in[3][6][3][bW-1:0] + accbin_in[4][6][3][bW-1:0] + accbin_in[5][6][3][bW-1:0] + accbin_in[6][6][3][bW-1:0] + accbin_in[7][6][3][bW-1:0] + accbin_in[8][6][3][bW-1:0] + accbin_in[9][6][3][bW-1:0] + accbin_in[10][6][3][bW-1:0] + accbin_in[11][6][3][bW-1:0] + accbin_in[12][6][3][bW-1:0] + accbin_in[13][6][3][bW-1:0] + accbin_in[14][6][3][bW-1:0] + accbin_in[15][6][3][bW-1:0] + accbin_in[16][6][3][bW-1:0] + accbin_in[17][6][3][bW-1:0];
assign sum_out[6][4][bW-1:0] = accbin_in[0][6][4][bW-1:0] + accbin_in[1][6][4][bW-1:0] + accbin_in[2][6][4][bW-1:0] + accbin_in[3][6][4][bW-1:0] + accbin_in[4][6][4][bW-1:0] + accbin_in[5][6][4][bW-1:0] + accbin_in[6][6][4][bW-1:0] + accbin_in[7][6][4][bW-1:0] + accbin_in[8][6][4][bW-1:0] + accbin_in[9][6][4][bW-1:0] + accbin_in[10][6][4][bW-1:0] + accbin_in[11][6][4][bW-1:0] + accbin_in[12][6][4][bW-1:0] + accbin_in[13][6][4][bW-1:0] + accbin_in[14][6][4][bW-1:0] + accbin_in[15][6][4][bW-1:0] + accbin_in[16][6][4][bW-1:0] + accbin_in[17][6][4][bW-1:0];
assign sum_out[6][5][bW-1:0] = accbin_in[0][6][5][bW-1:0] + accbin_in[1][6][5][bW-1:0] + accbin_in[2][6][5][bW-1:0] + accbin_in[3][6][5][bW-1:0] + accbin_in[4][6][5][bW-1:0] + accbin_in[5][6][5][bW-1:0] + accbin_in[6][6][5][bW-1:0] + accbin_in[7][6][5][bW-1:0] + accbin_in[8][6][5][bW-1:0] + accbin_in[9][6][5][bW-1:0] + accbin_in[10][6][5][bW-1:0] + accbin_in[11][6][5][bW-1:0] + accbin_in[12][6][5][bW-1:0] + accbin_in[13][6][5][bW-1:0] + accbin_in[14][6][5][bW-1:0] + accbin_in[15][6][5][bW-1:0] + accbin_in[16][6][5][bW-1:0] + accbin_in[17][6][5][bW-1:0];
assign sum_out[6][6][bW-1:0] = accbin_in[0][6][6][bW-1:0] + accbin_in[1][6][6][bW-1:0] + accbin_in[2][6][6][bW-1:0] + accbin_in[3][6][6][bW-1:0] + accbin_in[4][6][6][bW-1:0] + accbin_in[5][6][6][bW-1:0] + accbin_in[6][6][6][bW-1:0] + accbin_in[7][6][6][bW-1:0] + accbin_in[8][6][6][bW-1:0] + accbin_in[9][6][6][bW-1:0] + accbin_in[10][6][6][bW-1:0] + accbin_in[11][6][6][bW-1:0] + accbin_in[12][6][6][bW-1:0] + accbin_in[13][6][6][bW-1:0] + accbin_in[14][6][6][bW-1:0] + accbin_in[15][6][6][bW-1:0] + accbin_in[16][6][6][bW-1:0] + accbin_in[17][6][6][bW-1:0];
assign sum_out[6][7][bW-1:0] = accbin_in[0][6][7][bW-1:0] + accbin_in[1][6][7][bW-1:0] + accbin_in[2][6][7][bW-1:0] + accbin_in[3][6][7][bW-1:0] + accbin_in[4][6][7][bW-1:0] + accbin_in[5][6][7][bW-1:0] + accbin_in[6][6][7][bW-1:0] + accbin_in[7][6][7][bW-1:0] + accbin_in[8][6][7][bW-1:0] + accbin_in[9][6][7][bW-1:0] + accbin_in[10][6][7][bW-1:0] + accbin_in[11][6][7][bW-1:0] + accbin_in[12][6][7][bW-1:0] + accbin_in[13][6][7][bW-1:0] + accbin_in[14][6][7][bW-1:0] + accbin_in[15][6][7][bW-1:0] + accbin_in[16][6][7][bW-1:0] + accbin_in[17][6][7][bW-1:0];
assign sum_out[6][8][bW-1:0] = accbin_in[0][6][8][bW-1:0] + accbin_in[1][6][8][bW-1:0] + accbin_in[2][6][8][bW-1:0] + accbin_in[3][6][8][bW-1:0] + accbin_in[4][6][8][bW-1:0] + accbin_in[5][6][8][bW-1:0] + accbin_in[6][6][8][bW-1:0] + accbin_in[7][6][8][bW-1:0] + accbin_in[8][6][8][bW-1:0] + accbin_in[9][6][8][bW-1:0] + accbin_in[10][6][8][bW-1:0] + accbin_in[11][6][8][bW-1:0] + accbin_in[12][6][8][bW-1:0] + accbin_in[13][6][8][bW-1:0] + accbin_in[14][6][8][bW-1:0] + accbin_in[15][6][8][bW-1:0] + accbin_in[16][6][8][bW-1:0] + accbin_in[17][6][8][bW-1:0];
assign sum_out[6][9][bW-1:0] = accbin_in[0][6][9][bW-1:0] + accbin_in[1][6][9][bW-1:0] + accbin_in[2][6][9][bW-1:0] + accbin_in[3][6][9][bW-1:0] + accbin_in[4][6][9][bW-1:0] + accbin_in[5][6][9][bW-1:0] + accbin_in[6][6][9][bW-1:0] + accbin_in[7][6][9][bW-1:0] + accbin_in[8][6][9][bW-1:0] + accbin_in[9][6][9][bW-1:0] + accbin_in[10][6][9][bW-1:0] + accbin_in[11][6][9][bW-1:0] + accbin_in[12][6][9][bW-1:0] + accbin_in[13][6][9][bW-1:0] + accbin_in[14][6][9][bW-1:0] + accbin_in[15][6][9][bW-1:0] + accbin_in[16][6][9][bW-1:0] + accbin_in[17][6][9][bW-1:0];
assign sum_out[6][10][bW-1:0] = accbin_in[0][6][10][bW-1:0] + accbin_in[1][6][10][bW-1:0] + accbin_in[2][6][10][bW-1:0] + accbin_in[3][6][10][bW-1:0] + accbin_in[4][6][10][bW-1:0] + accbin_in[5][6][10][bW-1:0] + accbin_in[6][6][10][bW-1:0] + accbin_in[7][6][10][bW-1:0] + accbin_in[8][6][10][bW-1:0] + accbin_in[9][6][10][bW-1:0] + accbin_in[10][6][10][bW-1:0] + accbin_in[11][6][10][bW-1:0] + accbin_in[12][6][10][bW-1:0] + accbin_in[13][6][10][bW-1:0] + accbin_in[14][6][10][bW-1:0] + accbin_in[15][6][10][bW-1:0] + accbin_in[16][6][10][bW-1:0] + accbin_in[17][6][10][bW-1:0];
assign sum_out[6][11][bW-1:0] = accbin_in[0][6][11][bW-1:0] + accbin_in[1][6][11][bW-1:0] + accbin_in[2][6][11][bW-1:0] + accbin_in[3][6][11][bW-1:0] + accbin_in[4][6][11][bW-1:0] + accbin_in[5][6][11][bW-1:0] + accbin_in[6][6][11][bW-1:0] + accbin_in[7][6][11][bW-1:0] + accbin_in[8][6][11][bW-1:0] + accbin_in[9][6][11][bW-1:0] + accbin_in[10][6][11][bW-1:0] + accbin_in[11][6][11][bW-1:0] + accbin_in[12][6][11][bW-1:0] + accbin_in[13][6][11][bW-1:0] + accbin_in[14][6][11][bW-1:0] + accbin_in[15][6][11][bW-1:0] + accbin_in[16][6][11][bW-1:0] + accbin_in[17][6][11][bW-1:0];
assign sum_out[7][0][bW-1:0] = accbin_in[0][7][0][bW-1:0] + accbin_in[1][7][0][bW-1:0] + accbin_in[2][7][0][bW-1:0] + accbin_in[3][7][0][bW-1:0] + accbin_in[4][7][0][bW-1:0] + accbin_in[5][7][0][bW-1:0] + accbin_in[6][7][0][bW-1:0] + accbin_in[7][7][0][bW-1:0] + accbin_in[8][7][0][bW-1:0] + accbin_in[9][7][0][bW-1:0] + accbin_in[10][7][0][bW-1:0] + accbin_in[11][7][0][bW-1:0] + accbin_in[12][7][0][bW-1:0] + accbin_in[13][7][0][bW-1:0] + accbin_in[14][7][0][bW-1:0] + accbin_in[15][7][0][bW-1:0] + accbin_in[16][7][0][bW-1:0] + accbin_in[17][7][0][bW-1:0];
assign sum_out[7][1][bW-1:0] = accbin_in[0][7][1][bW-1:0] + accbin_in[1][7][1][bW-1:0] + accbin_in[2][7][1][bW-1:0] + accbin_in[3][7][1][bW-1:0] + accbin_in[4][7][1][bW-1:0] + accbin_in[5][7][1][bW-1:0] + accbin_in[6][7][1][bW-1:0] + accbin_in[7][7][1][bW-1:0] + accbin_in[8][7][1][bW-1:0] + accbin_in[9][7][1][bW-1:0] + accbin_in[10][7][1][bW-1:0] + accbin_in[11][7][1][bW-1:0] + accbin_in[12][7][1][bW-1:0] + accbin_in[13][7][1][bW-1:0] + accbin_in[14][7][1][bW-1:0] + accbin_in[15][7][1][bW-1:0] + accbin_in[16][7][1][bW-1:0] + accbin_in[17][7][1][bW-1:0];
assign sum_out[7][2][bW-1:0] = accbin_in[0][7][2][bW-1:0] + accbin_in[1][7][2][bW-1:0] + accbin_in[2][7][2][bW-1:0] + accbin_in[3][7][2][bW-1:0] + accbin_in[4][7][2][bW-1:0] + accbin_in[5][7][2][bW-1:0] + accbin_in[6][7][2][bW-1:0] + accbin_in[7][7][2][bW-1:0] + accbin_in[8][7][2][bW-1:0] + accbin_in[9][7][2][bW-1:0] + accbin_in[10][7][2][bW-1:0] + accbin_in[11][7][2][bW-1:0] + accbin_in[12][7][2][bW-1:0] + accbin_in[13][7][2][bW-1:0] + accbin_in[14][7][2][bW-1:0] + accbin_in[15][7][2][bW-1:0] + accbin_in[16][7][2][bW-1:0] + accbin_in[17][7][2][bW-1:0];
assign sum_out[7][3][bW-1:0] = accbin_in[0][7][3][bW-1:0] + accbin_in[1][7][3][bW-1:0] + accbin_in[2][7][3][bW-1:0] + accbin_in[3][7][3][bW-1:0] + accbin_in[4][7][3][bW-1:0] + accbin_in[5][7][3][bW-1:0] + accbin_in[6][7][3][bW-1:0] + accbin_in[7][7][3][bW-1:0] + accbin_in[8][7][3][bW-1:0] + accbin_in[9][7][3][bW-1:0] + accbin_in[10][7][3][bW-1:0] + accbin_in[11][7][3][bW-1:0] + accbin_in[12][7][3][bW-1:0] + accbin_in[13][7][3][bW-1:0] + accbin_in[14][7][3][bW-1:0] + accbin_in[15][7][3][bW-1:0] + accbin_in[16][7][3][bW-1:0] + accbin_in[17][7][3][bW-1:0];
assign sum_out[7][4][bW-1:0] = accbin_in[0][7][4][bW-1:0] + accbin_in[1][7][4][bW-1:0] + accbin_in[2][7][4][bW-1:0] + accbin_in[3][7][4][bW-1:0] + accbin_in[4][7][4][bW-1:0] + accbin_in[5][7][4][bW-1:0] + accbin_in[6][7][4][bW-1:0] + accbin_in[7][7][4][bW-1:0] + accbin_in[8][7][4][bW-1:0] + accbin_in[9][7][4][bW-1:0] + accbin_in[10][7][4][bW-1:0] + accbin_in[11][7][4][bW-1:0] + accbin_in[12][7][4][bW-1:0] + accbin_in[13][7][4][bW-1:0] + accbin_in[14][7][4][bW-1:0] + accbin_in[15][7][4][bW-1:0] + accbin_in[16][7][4][bW-1:0] + accbin_in[17][7][4][bW-1:0];
assign sum_out[7][5][bW-1:0] = accbin_in[0][7][5][bW-1:0] + accbin_in[1][7][5][bW-1:0] + accbin_in[2][7][5][bW-1:0] + accbin_in[3][7][5][bW-1:0] + accbin_in[4][7][5][bW-1:0] + accbin_in[5][7][5][bW-1:0] + accbin_in[6][7][5][bW-1:0] + accbin_in[7][7][5][bW-1:0] + accbin_in[8][7][5][bW-1:0] + accbin_in[9][7][5][bW-1:0] + accbin_in[10][7][5][bW-1:0] + accbin_in[11][7][5][bW-1:0] + accbin_in[12][7][5][bW-1:0] + accbin_in[13][7][5][bW-1:0] + accbin_in[14][7][5][bW-1:0] + accbin_in[15][7][5][bW-1:0] + accbin_in[16][7][5][bW-1:0] + accbin_in[17][7][5][bW-1:0];
assign sum_out[7][6][bW-1:0] = accbin_in[0][7][6][bW-1:0] + accbin_in[1][7][6][bW-1:0] + accbin_in[2][7][6][bW-1:0] + accbin_in[3][7][6][bW-1:0] + accbin_in[4][7][6][bW-1:0] + accbin_in[5][7][6][bW-1:0] + accbin_in[6][7][6][bW-1:0] + accbin_in[7][7][6][bW-1:0] + accbin_in[8][7][6][bW-1:0] + accbin_in[9][7][6][bW-1:0] + accbin_in[10][7][6][bW-1:0] + accbin_in[11][7][6][bW-1:0] + accbin_in[12][7][6][bW-1:0] + accbin_in[13][7][6][bW-1:0] + accbin_in[14][7][6][bW-1:0] + accbin_in[15][7][6][bW-1:0] + accbin_in[16][7][6][bW-1:0] + accbin_in[17][7][6][bW-1:0];
assign sum_out[7][7][bW-1:0] = accbin_in[0][7][7][bW-1:0] + accbin_in[1][7][7][bW-1:0] + accbin_in[2][7][7][bW-1:0] + accbin_in[3][7][7][bW-1:0] + accbin_in[4][7][7][bW-1:0] + accbin_in[5][7][7][bW-1:0] + accbin_in[6][7][7][bW-1:0] + accbin_in[7][7][7][bW-1:0] + accbin_in[8][7][7][bW-1:0] + accbin_in[9][7][7][bW-1:0] + accbin_in[10][7][7][bW-1:0] + accbin_in[11][7][7][bW-1:0] + accbin_in[12][7][7][bW-1:0] + accbin_in[13][7][7][bW-1:0] + accbin_in[14][7][7][bW-1:0] + accbin_in[15][7][7][bW-1:0] + accbin_in[16][7][7][bW-1:0] + accbin_in[17][7][7][bW-1:0];
assign sum_out[7][8][bW-1:0] = accbin_in[0][7][8][bW-1:0] + accbin_in[1][7][8][bW-1:0] + accbin_in[2][7][8][bW-1:0] + accbin_in[3][7][8][bW-1:0] + accbin_in[4][7][8][bW-1:0] + accbin_in[5][7][8][bW-1:0] + accbin_in[6][7][8][bW-1:0] + accbin_in[7][7][8][bW-1:0] + accbin_in[8][7][8][bW-1:0] + accbin_in[9][7][8][bW-1:0] + accbin_in[10][7][8][bW-1:0] + accbin_in[11][7][8][bW-1:0] + accbin_in[12][7][8][bW-1:0] + accbin_in[13][7][8][bW-1:0] + accbin_in[14][7][8][bW-1:0] + accbin_in[15][7][8][bW-1:0] + accbin_in[16][7][8][bW-1:0] + accbin_in[17][7][8][bW-1:0];
assign sum_out[7][9][bW-1:0] = accbin_in[0][7][9][bW-1:0] + accbin_in[1][7][9][bW-1:0] + accbin_in[2][7][9][bW-1:0] + accbin_in[3][7][9][bW-1:0] + accbin_in[4][7][9][bW-1:0] + accbin_in[5][7][9][bW-1:0] + accbin_in[6][7][9][bW-1:0] + accbin_in[7][7][9][bW-1:0] + accbin_in[8][7][9][bW-1:0] + accbin_in[9][7][9][bW-1:0] + accbin_in[10][7][9][bW-1:0] + accbin_in[11][7][9][bW-1:0] + accbin_in[12][7][9][bW-1:0] + accbin_in[13][7][9][bW-1:0] + accbin_in[14][7][9][bW-1:0] + accbin_in[15][7][9][bW-1:0] + accbin_in[16][7][9][bW-1:0] + accbin_in[17][7][9][bW-1:0];
assign sum_out[7][10][bW-1:0] = accbin_in[0][7][10][bW-1:0] + accbin_in[1][7][10][bW-1:0] + accbin_in[2][7][10][bW-1:0] + accbin_in[3][7][10][bW-1:0] + accbin_in[4][7][10][bW-1:0] + accbin_in[5][7][10][bW-1:0] + accbin_in[6][7][10][bW-1:0] + accbin_in[7][7][10][bW-1:0] + accbin_in[8][7][10][bW-1:0] + accbin_in[9][7][10][bW-1:0] + accbin_in[10][7][10][bW-1:0] + accbin_in[11][7][10][bW-1:0] + accbin_in[12][7][10][bW-1:0] + accbin_in[13][7][10][bW-1:0] + accbin_in[14][7][10][bW-1:0] + accbin_in[15][7][10][bW-1:0] + accbin_in[16][7][10][bW-1:0] + accbin_in[17][7][10][bW-1:0];
assign sum_out[7][11][bW-1:0] = accbin_in[0][7][11][bW-1:0] + accbin_in[1][7][11][bW-1:0] + accbin_in[2][7][11][bW-1:0] + accbin_in[3][7][11][bW-1:0] + accbin_in[4][7][11][bW-1:0] + accbin_in[5][7][11][bW-1:0] + accbin_in[6][7][11][bW-1:0] + accbin_in[7][7][11][bW-1:0] + accbin_in[8][7][11][bW-1:0] + accbin_in[9][7][11][bW-1:0] + accbin_in[10][7][11][bW-1:0] + accbin_in[11][7][11][bW-1:0] + accbin_in[12][7][11][bW-1:0] + accbin_in[13][7][11][bW-1:0] + accbin_in[14][7][11][bW-1:0] + accbin_in[15][7][11][bW-1:0] + accbin_in[16][7][11][bW-1:0] + accbin_in[17][7][11][bW-1:0];
assign sum_out[8][0][bW-1:0] = accbin_in[0][8][0][bW-1:0] + accbin_in[1][8][0][bW-1:0] + accbin_in[2][8][0][bW-1:0] + accbin_in[3][8][0][bW-1:0] + accbin_in[4][8][0][bW-1:0] + accbin_in[5][8][0][bW-1:0] + accbin_in[6][8][0][bW-1:0] + accbin_in[7][8][0][bW-1:0] + accbin_in[8][8][0][bW-1:0] + accbin_in[9][8][0][bW-1:0] + accbin_in[10][8][0][bW-1:0] + accbin_in[11][8][0][bW-1:0] + accbin_in[12][8][0][bW-1:0] + accbin_in[13][8][0][bW-1:0] + accbin_in[14][8][0][bW-1:0] + accbin_in[15][8][0][bW-1:0] + accbin_in[16][8][0][bW-1:0] + accbin_in[17][8][0][bW-1:0];
assign sum_out[8][1][bW-1:0] = accbin_in[0][8][1][bW-1:0] + accbin_in[1][8][1][bW-1:0] + accbin_in[2][8][1][bW-1:0] + accbin_in[3][8][1][bW-1:0] + accbin_in[4][8][1][bW-1:0] + accbin_in[5][8][1][bW-1:0] + accbin_in[6][8][1][bW-1:0] + accbin_in[7][8][1][bW-1:0] + accbin_in[8][8][1][bW-1:0] + accbin_in[9][8][1][bW-1:0] + accbin_in[10][8][1][bW-1:0] + accbin_in[11][8][1][bW-1:0] + accbin_in[12][8][1][bW-1:0] + accbin_in[13][8][1][bW-1:0] + accbin_in[14][8][1][bW-1:0] + accbin_in[15][8][1][bW-1:0] + accbin_in[16][8][1][bW-1:0] + accbin_in[17][8][1][bW-1:0];
assign sum_out[8][2][bW-1:0] = accbin_in[0][8][2][bW-1:0] + accbin_in[1][8][2][bW-1:0] + accbin_in[2][8][2][bW-1:0] + accbin_in[3][8][2][bW-1:0] + accbin_in[4][8][2][bW-1:0] + accbin_in[5][8][2][bW-1:0] + accbin_in[6][8][2][bW-1:0] + accbin_in[7][8][2][bW-1:0] + accbin_in[8][8][2][bW-1:0] + accbin_in[9][8][2][bW-1:0] + accbin_in[10][8][2][bW-1:0] + accbin_in[11][8][2][bW-1:0] + accbin_in[12][8][2][bW-1:0] + accbin_in[13][8][2][bW-1:0] + accbin_in[14][8][2][bW-1:0] + accbin_in[15][8][2][bW-1:0] + accbin_in[16][8][2][bW-1:0] + accbin_in[17][8][2][bW-1:0];
assign sum_out[8][3][bW-1:0] = accbin_in[0][8][3][bW-1:0] + accbin_in[1][8][3][bW-1:0] + accbin_in[2][8][3][bW-1:0] + accbin_in[3][8][3][bW-1:0] + accbin_in[4][8][3][bW-1:0] + accbin_in[5][8][3][bW-1:0] + accbin_in[6][8][3][bW-1:0] + accbin_in[7][8][3][bW-1:0] + accbin_in[8][8][3][bW-1:0] + accbin_in[9][8][3][bW-1:0] + accbin_in[10][8][3][bW-1:0] + accbin_in[11][8][3][bW-1:0] + accbin_in[12][8][3][bW-1:0] + accbin_in[13][8][3][bW-1:0] + accbin_in[14][8][3][bW-1:0] + accbin_in[15][8][3][bW-1:0] + accbin_in[16][8][3][bW-1:0] + accbin_in[17][8][3][bW-1:0];
assign sum_out[8][4][bW-1:0] = accbin_in[0][8][4][bW-1:0] + accbin_in[1][8][4][bW-1:0] + accbin_in[2][8][4][bW-1:0] + accbin_in[3][8][4][bW-1:0] + accbin_in[4][8][4][bW-1:0] + accbin_in[5][8][4][bW-1:0] + accbin_in[6][8][4][bW-1:0] + accbin_in[7][8][4][bW-1:0] + accbin_in[8][8][4][bW-1:0] + accbin_in[9][8][4][bW-1:0] + accbin_in[10][8][4][bW-1:0] + accbin_in[11][8][4][bW-1:0] + accbin_in[12][8][4][bW-1:0] + accbin_in[13][8][4][bW-1:0] + accbin_in[14][8][4][bW-1:0] + accbin_in[15][8][4][bW-1:0] + accbin_in[16][8][4][bW-1:0] + accbin_in[17][8][4][bW-1:0];
assign sum_out[8][5][bW-1:0] = accbin_in[0][8][5][bW-1:0] + accbin_in[1][8][5][bW-1:0] + accbin_in[2][8][5][bW-1:0] + accbin_in[3][8][5][bW-1:0] + accbin_in[4][8][5][bW-1:0] + accbin_in[5][8][5][bW-1:0] + accbin_in[6][8][5][bW-1:0] + accbin_in[7][8][5][bW-1:0] + accbin_in[8][8][5][bW-1:0] + accbin_in[9][8][5][bW-1:0] + accbin_in[10][8][5][bW-1:0] + accbin_in[11][8][5][bW-1:0] + accbin_in[12][8][5][bW-1:0] + accbin_in[13][8][5][bW-1:0] + accbin_in[14][8][5][bW-1:0] + accbin_in[15][8][5][bW-1:0] + accbin_in[16][8][5][bW-1:0] + accbin_in[17][8][5][bW-1:0];
assign sum_out[8][6][bW-1:0] = accbin_in[0][8][6][bW-1:0] + accbin_in[1][8][6][bW-1:0] + accbin_in[2][8][6][bW-1:0] + accbin_in[3][8][6][bW-1:0] + accbin_in[4][8][6][bW-1:0] + accbin_in[5][8][6][bW-1:0] + accbin_in[6][8][6][bW-1:0] + accbin_in[7][8][6][bW-1:0] + accbin_in[8][8][6][bW-1:0] + accbin_in[9][8][6][bW-1:0] + accbin_in[10][8][6][bW-1:0] + accbin_in[11][8][6][bW-1:0] + accbin_in[12][8][6][bW-1:0] + accbin_in[13][8][6][bW-1:0] + accbin_in[14][8][6][bW-1:0] + accbin_in[15][8][6][bW-1:0] + accbin_in[16][8][6][bW-1:0] + accbin_in[17][8][6][bW-1:0];
assign sum_out[8][7][bW-1:0] = accbin_in[0][8][7][bW-1:0] + accbin_in[1][8][7][bW-1:0] + accbin_in[2][8][7][bW-1:0] + accbin_in[3][8][7][bW-1:0] + accbin_in[4][8][7][bW-1:0] + accbin_in[5][8][7][bW-1:0] + accbin_in[6][8][7][bW-1:0] + accbin_in[7][8][7][bW-1:0] + accbin_in[8][8][7][bW-1:0] + accbin_in[9][8][7][bW-1:0] + accbin_in[10][8][7][bW-1:0] + accbin_in[11][8][7][bW-1:0] + accbin_in[12][8][7][bW-1:0] + accbin_in[13][8][7][bW-1:0] + accbin_in[14][8][7][bW-1:0] + accbin_in[15][8][7][bW-1:0] + accbin_in[16][8][7][bW-1:0] + accbin_in[17][8][7][bW-1:0];
assign sum_out[8][8][bW-1:0] = accbin_in[0][8][8][bW-1:0] + accbin_in[1][8][8][bW-1:0] + accbin_in[2][8][8][bW-1:0] + accbin_in[3][8][8][bW-1:0] + accbin_in[4][8][8][bW-1:0] + accbin_in[5][8][8][bW-1:0] + accbin_in[6][8][8][bW-1:0] + accbin_in[7][8][8][bW-1:0] + accbin_in[8][8][8][bW-1:0] + accbin_in[9][8][8][bW-1:0] + accbin_in[10][8][8][bW-1:0] + accbin_in[11][8][8][bW-1:0] + accbin_in[12][8][8][bW-1:0] + accbin_in[13][8][8][bW-1:0] + accbin_in[14][8][8][bW-1:0] + accbin_in[15][8][8][bW-1:0] + accbin_in[16][8][8][bW-1:0] + accbin_in[17][8][8][bW-1:0];
assign sum_out[8][9][bW-1:0] = accbin_in[0][8][9][bW-1:0] + accbin_in[1][8][9][bW-1:0] + accbin_in[2][8][9][bW-1:0] + accbin_in[3][8][9][bW-1:0] + accbin_in[4][8][9][bW-1:0] + accbin_in[5][8][9][bW-1:0] + accbin_in[6][8][9][bW-1:0] + accbin_in[7][8][9][bW-1:0] + accbin_in[8][8][9][bW-1:0] + accbin_in[9][8][9][bW-1:0] + accbin_in[10][8][9][bW-1:0] + accbin_in[11][8][9][bW-1:0] + accbin_in[12][8][9][bW-1:0] + accbin_in[13][8][9][bW-1:0] + accbin_in[14][8][9][bW-1:0] + accbin_in[15][8][9][bW-1:0] + accbin_in[16][8][9][bW-1:0] + accbin_in[17][8][9][bW-1:0];
assign sum_out[8][10][bW-1:0] = accbin_in[0][8][10][bW-1:0] + accbin_in[1][8][10][bW-1:0] + accbin_in[2][8][10][bW-1:0] + accbin_in[3][8][10][bW-1:0] + accbin_in[4][8][10][bW-1:0] + accbin_in[5][8][10][bW-1:0] + accbin_in[6][8][10][bW-1:0] + accbin_in[7][8][10][bW-1:0] + accbin_in[8][8][10][bW-1:0] + accbin_in[9][8][10][bW-1:0] + accbin_in[10][8][10][bW-1:0] + accbin_in[11][8][10][bW-1:0] + accbin_in[12][8][10][bW-1:0] + accbin_in[13][8][10][bW-1:0] + accbin_in[14][8][10][bW-1:0] + accbin_in[15][8][10][bW-1:0] + accbin_in[16][8][10][bW-1:0] + accbin_in[17][8][10][bW-1:0];
assign sum_out[8][11][bW-1:0] = accbin_in[0][8][11][bW-1:0] + accbin_in[1][8][11][bW-1:0] + accbin_in[2][8][11][bW-1:0] + accbin_in[3][8][11][bW-1:0] + accbin_in[4][8][11][bW-1:0] + accbin_in[5][8][11][bW-1:0] + accbin_in[6][8][11][bW-1:0] + accbin_in[7][8][11][bW-1:0] + accbin_in[8][8][11][bW-1:0] + accbin_in[9][8][11][bW-1:0] + accbin_in[10][8][11][bW-1:0] + accbin_in[11][8][11][bW-1:0] + accbin_in[12][8][11][bW-1:0] + accbin_in[13][8][11][bW-1:0] + accbin_in[14][8][11][bW-1:0] + accbin_in[15][8][11][bW-1:0] + accbin_in[16][8][11][bW-1:0] + accbin_in[17][8][11][bW-1:0];
assign sum_out[9][0][bW-1:0] = accbin_in[0][9][0][bW-1:0] + accbin_in[1][9][0][bW-1:0] + accbin_in[2][9][0][bW-1:0] + accbin_in[3][9][0][bW-1:0] + accbin_in[4][9][0][bW-1:0] + accbin_in[5][9][0][bW-1:0] + accbin_in[6][9][0][bW-1:0] + accbin_in[7][9][0][bW-1:0] + accbin_in[8][9][0][bW-1:0] + accbin_in[9][9][0][bW-1:0] + accbin_in[10][9][0][bW-1:0] + accbin_in[11][9][0][bW-1:0] + accbin_in[12][9][0][bW-1:0] + accbin_in[13][9][0][bW-1:0] + accbin_in[14][9][0][bW-1:0] + accbin_in[15][9][0][bW-1:0] + accbin_in[16][9][0][bW-1:0] + accbin_in[17][9][0][bW-1:0];
assign sum_out[9][1][bW-1:0] = accbin_in[0][9][1][bW-1:0] + accbin_in[1][9][1][bW-1:0] + accbin_in[2][9][1][bW-1:0] + accbin_in[3][9][1][bW-1:0] + accbin_in[4][9][1][bW-1:0] + accbin_in[5][9][1][bW-1:0] + accbin_in[6][9][1][bW-1:0] + accbin_in[7][9][1][bW-1:0] + accbin_in[8][9][1][bW-1:0] + accbin_in[9][9][1][bW-1:0] + accbin_in[10][9][1][bW-1:0] + accbin_in[11][9][1][bW-1:0] + accbin_in[12][9][1][bW-1:0] + accbin_in[13][9][1][bW-1:0] + accbin_in[14][9][1][bW-1:0] + accbin_in[15][9][1][bW-1:0] + accbin_in[16][9][1][bW-1:0] + accbin_in[17][9][1][bW-1:0];
assign sum_out[9][2][bW-1:0] = accbin_in[0][9][2][bW-1:0] + accbin_in[1][9][2][bW-1:0] + accbin_in[2][9][2][bW-1:0] + accbin_in[3][9][2][bW-1:0] + accbin_in[4][9][2][bW-1:0] + accbin_in[5][9][2][bW-1:0] + accbin_in[6][9][2][bW-1:0] + accbin_in[7][9][2][bW-1:0] + accbin_in[8][9][2][bW-1:0] + accbin_in[9][9][2][bW-1:0] + accbin_in[10][9][2][bW-1:0] + accbin_in[11][9][2][bW-1:0] + accbin_in[12][9][2][bW-1:0] + accbin_in[13][9][2][bW-1:0] + accbin_in[14][9][2][bW-1:0] + accbin_in[15][9][2][bW-1:0] + accbin_in[16][9][2][bW-1:0] + accbin_in[17][9][2][bW-1:0];
assign sum_out[9][3][bW-1:0] = accbin_in[0][9][3][bW-1:0] + accbin_in[1][9][3][bW-1:0] + accbin_in[2][9][3][bW-1:0] + accbin_in[3][9][3][bW-1:0] + accbin_in[4][9][3][bW-1:0] + accbin_in[5][9][3][bW-1:0] + accbin_in[6][9][3][bW-1:0] + accbin_in[7][9][3][bW-1:0] + accbin_in[8][9][3][bW-1:0] + accbin_in[9][9][3][bW-1:0] + accbin_in[10][9][3][bW-1:0] + accbin_in[11][9][3][bW-1:0] + accbin_in[12][9][3][bW-1:0] + accbin_in[13][9][3][bW-1:0] + accbin_in[14][9][3][bW-1:0] + accbin_in[15][9][3][bW-1:0] + accbin_in[16][9][3][bW-1:0] + accbin_in[17][9][3][bW-1:0];
assign sum_out[9][4][bW-1:0] = accbin_in[0][9][4][bW-1:0] + accbin_in[1][9][4][bW-1:0] + accbin_in[2][9][4][bW-1:0] + accbin_in[3][9][4][bW-1:0] + accbin_in[4][9][4][bW-1:0] + accbin_in[5][9][4][bW-1:0] + accbin_in[6][9][4][bW-1:0] + accbin_in[7][9][4][bW-1:0] + accbin_in[8][9][4][bW-1:0] + accbin_in[9][9][4][bW-1:0] + accbin_in[10][9][4][bW-1:0] + accbin_in[11][9][4][bW-1:0] + accbin_in[12][9][4][bW-1:0] + accbin_in[13][9][4][bW-1:0] + accbin_in[14][9][4][bW-1:0] + accbin_in[15][9][4][bW-1:0] + accbin_in[16][9][4][bW-1:0] + accbin_in[17][9][4][bW-1:0];
assign sum_out[9][5][bW-1:0] = accbin_in[0][9][5][bW-1:0] + accbin_in[1][9][5][bW-1:0] + accbin_in[2][9][5][bW-1:0] + accbin_in[3][9][5][bW-1:0] + accbin_in[4][9][5][bW-1:0] + accbin_in[5][9][5][bW-1:0] + accbin_in[6][9][5][bW-1:0] + accbin_in[7][9][5][bW-1:0] + accbin_in[8][9][5][bW-1:0] + accbin_in[9][9][5][bW-1:0] + accbin_in[10][9][5][bW-1:0] + accbin_in[11][9][5][bW-1:0] + accbin_in[12][9][5][bW-1:0] + accbin_in[13][9][5][bW-1:0] + accbin_in[14][9][5][bW-1:0] + accbin_in[15][9][5][bW-1:0] + accbin_in[16][9][5][bW-1:0] + accbin_in[17][9][5][bW-1:0];
assign sum_out[9][6][bW-1:0] = accbin_in[0][9][6][bW-1:0] + accbin_in[1][9][6][bW-1:0] + accbin_in[2][9][6][bW-1:0] + accbin_in[3][9][6][bW-1:0] + accbin_in[4][9][6][bW-1:0] + accbin_in[5][9][6][bW-1:0] + accbin_in[6][9][6][bW-1:0] + accbin_in[7][9][6][bW-1:0] + accbin_in[8][9][6][bW-1:0] + accbin_in[9][9][6][bW-1:0] + accbin_in[10][9][6][bW-1:0] + accbin_in[11][9][6][bW-1:0] + accbin_in[12][9][6][bW-1:0] + accbin_in[13][9][6][bW-1:0] + accbin_in[14][9][6][bW-1:0] + accbin_in[15][9][6][bW-1:0] + accbin_in[16][9][6][bW-1:0] + accbin_in[17][9][6][bW-1:0];
assign sum_out[9][7][bW-1:0] = accbin_in[0][9][7][bW-1:0] + accbin_in[1][9][7][bW-1:0] + accbin_in[2][9][7][bW-1:0] + accbin_in[3][9][7][bW-1:0] + accbin_in[4][9][7][bW-1:0] + accbin_in[5][9][7][bW-1:0] + accbin_in[6][9][7][bW-1:0] + accbin_in[7][9][7][bW-1:0] + accbin_in[8][9][7][bW-1:0] + accbin_in[9][9][7][bW-1:0] + accbin_in[10][9][7][bW-1:0] + accbin_in[11][9][7][bW-1:0] + accbin_in[12][9][7][bW-1:0] + accbin_in[13][9][7][bW-1:0] + accbin_in[14][9][7][bW-1:0] + accbin_in[15][9][7][bW-1:0] + accbin_in[16][9][7][bW-1:0] + accbin_in[17][9][7][bW-1:0];
assign sum_out[9][8][bW-1:0] = accbin_in[0][9][8][bW-1:0] + accbin_in[1][9][8][bW-1:0] + accbin_in[2][9][8][bW-1:0] + accbin_in[3][9][8][bW-1:0] + accbin_in[4][9][8][bW-1:0] + accbin_in[5][9][8][bW-1:0] + accbin_in[6][9][8][bW-1:0] + accbin_in[7][9][8][bW-1:0] + accbin_in[8][9][8][bW-1:0] + accbin_in[9][9][8][bW-1:0] + accbin_in[10][9][8][bW-1:0] + accbin_in[11][9][8][bW-1:0] + accbin_in[12][9][8][bW-1:0] + accbin_in[13][9][8][bW-1:0] + accbin_in[14][9][8][bW-1:0] + accbin_in[15][9][8][bW-1:0] + accbin_in[16][9][8][bW-1:0] + accbin_in[17][9][8][bW-1:0];
assign sum_out[9][9][bW-1:0] = accbin_in[0][9][9][bW-1:0] + accbin_in[1][9][9][bW-1:0] + accbin_in[2][9][9][bW-1:0] + accbin_in[3][9][9][bW-1:0] + accbin_in[4][9][9][bW-1:0] + accbin_in[5][9][9][bW-1:0] + accbin_in[6][9][9][bW-1:0] + accbin_in[7][9][9][bW-1:0] + accbin_in[8][9][9][bW-1:0] + accbin_in[9][9][9][bW-1:0] + accbin_in[10][9][9][bW-1:0] + accbin_in[11][9][9][bW-1:0] + accbin_in[12][9][9][bW-1:0] + accbin_in[13][9][9][bW-1:0] + accbin_in[14][9][9][bW-1:0] + accbin_in[15][9][9][bW-1:0] + accbin_in[16][9][9][bW-1:0] + accbin_in[17][9][9][bW-1:0];
assign sum_out[9][10][bW-1:0] = accbin_in[0][9][10][bW-1:0] + accbin_in[1][9][10][bW-1:0] + accbin_in[2][9][10][bW-1:0] + accbin_in[3][9][10][bW-1:0] + accbin_in[4][9][10][bW-1:0] + accbin_in[5][9][10][bW-1:0] + accbin_in[6][9][10][bW-1:0] + accbin_in[7][9][10][bW-1:0] + accbin_in[8][9][10][bW-1:0] + accbin_in[9][9][10][bW-1:0] + accbin_in[10][9][10][bW-1:0] + accbin_in[11][9][10][bW-1:0] + accbin_in[12][9][10][bW-1:0] + accbin_in[13][9][10][bW-1:0] + accbin_in[14][9][10][bW-1:0] + accbin_in[15][9][10][bW-1:0] + accbin_in[16][9][10][bW-1:0] + accbin_in[17][9][10][bW-1:0];
assign sum_out[9][11][bW-1:0] = accbin_in[0][9][11][bW-1:0] + accbin_in[1][9][11][bW-1:0] + accbin_in[2][9][11][bW-1:0] + accbin_in[3][9][11][bW-1:0] + accbin_in[4][9][11][bW-1:0] + accbin_in[5][9][11][bW-1:0] + accbin_in[6][9][11][bW-1:0] + accbin_in[7][9][11][bW-1:0] + accbin_in[8][9][11][bW-1:0] + accbin_in[9][9][11][bW-1:0] + accbin_in[10][9][11][bW-1:0] + accbin_in[11][9][11][bW-1:0] + accbin_in[12][9][11][bW-1:0] + accbin_in[13][9][11][bW-1:0] + accbin_in[14][9][11][bW-1:0] + accbin_in[15][9][11][bW-1:0] + accbin_in[16][9][11][bW-1:0] + accbin_in[17][9][11][bW-1:0];
assign sum_out[10][0][bW-1:0] = accbin_in[0][10][0][bW-1:0] + accbin_in[1][10][0][bW-1:0] + accbin_in[2][10][0][bW-1:0] + accbin_in[3][10][0][bW-1:0] + accbin_in[4][10][0][bW-1:0] + accbin_in[5][10][0][bW-1:0] + accbin_in[6][10][0][bW-1:0] + accbin_in[7][10][0][bW-1:0] + accbin_in[8][10][0][bW-1:0] + accbin_in[9][10][0][bW-1:0] + accbin_in[10][10][0][bW-1:0] + accbin_in[11][10][0][bW-1:0] + accbin_in[12][10][0][bW-1:0] + accbin_in[13][10][0][bW-1:0] + accbin_in[14][10][0][bW-1:0] + accbin_in[15][10][0][bW-1:0] + accbin_in[16][10][0][bW-1:0] + accbin_in[17][10][0][bW-1:0];
assign sum_out[10][1][bW-1:0] = accbin_in[0][10][1][bW-1:0] + accbin_in[1][10][1][bW-1:0] + accbin_in[2][10][1][bW-1:0] + accbin_in[3][10][1][bW-1:0] + accbin_in[4][10][1][bW-1:0] + accbin_in[5][10][1][bW-1:0] + accbin_in[6][10][1][bW-1:0] + accbin_in[7][10][1][bW-1:0] + accbin_in[8][10][1][bW-1:0] + accbin_in[9][10][1][bW-1:0] + accbin_in[10][10][1][bW-1:0] + accbin_in[11][10][1][bW-1:0] + accbin_in[12][10][1][bW-1:0] + accbin_in[13][10][1][bW-1:0] + accbin_in[14][10][1][bW-1:0] + accbin_in[15][10][1][bW-1:0] + accbin_in[16][10][1][bW-1:0] + accbin_in[17][10][1][bW-1:0];
assign sum_out[10][2][bW-1:0] = accbin_in[0][10][2][bW-1:0] + accbin_in[1][10][2][bW-1:0] + accbin_in[2][10][2][bW-1:0] + accbin_in[3][10][2][bW-1:0] + accbin_in[4][10][2][bW-1:0] + accbin_in[5][10][2][bW-1:0] + accbin_in[6][10][2][bW-1:0] + accbin_in[7][10][2][bW-1:0] + accbin_in[8][10][2][bW-1:0] + accbin_in[9][10][2][bW-1:0] + accbin_in[10][10][2][bW-1:0] + accbin_in[11][10][2][bW-1:0] + accbin_in[12][10][2][bW-1:0] + accbin_in[13][10][2][bW-1:0] + accbin_in[14][10][2][bW-1:0] + accbin_in[15][10][2][bW-1:0] + accbin_in[16][10][2][bW-1:0] + accbin_in[17][10][2][bW-1:0];
assign sum_out[10][3][bW-1:0] = accbin_in[0][10][3][bW-1:0] + accbin_in[1][10][3][bW-1:0] + accbin_in[2][10][3][bW-1:0] + accbin_in[3][10][3][bW-1:0] + accbin_in[4][10][3][bW-1:0] + accbin_in[5][10][3][bW-1:0] + accbin_in[6][10][3][bW-1:0] + accbin_in[7][10][3][bW-1:0] + accbin_in[8][10][3][bW-1:0] + accbin_in[9][10][3][bW-1:0] + accbin_in[10][10][3][bW-1:0] + accbin_in[11][10][3][bW-1:0] + accbin_in[12][10][3][bW-1:0] + accbin_in[13][10][3][bW-1:0] + accbin_in[14][10][3][bW-1:0] + accbin_in[15][10][3][bW-1:0] + accbin_in[16][10][3][bW-1:0] + accbin_in[17][10][3][bW-1:0];
assign sum_out[10][4][bW-1:0] = accbin_in[0][10][4][bW-1:0] + accbin_in[1][10][4][bW-1:0] + accbin_in[2][10][4][bW-1:0] + accbin_in[3][10][4][bW-1:0] + accbin_in[4][10][4][bW-1:0] + accbin_in[5][10][4][bW-1:0] + accbin_in[6][10][4][bW-1:0] + accbin_in[7][10][4][bW-1:0] + accbin_in[8][10][4][bW-1:0] + accbin_in[9][10][4][bW-1:0] + accbin_in[10][10][4][bW-1:0] + accbin_in[11][10][4][bW-1:0] + accbin_in[12][10][4][bW-1:0] + accbin_in[13][10][4][bW-1:0] + accbin_in[14][10][4][bW-1:0] + accbin_in[15][10][4][bW-1:0] + accbin_in[16][10][4][bW-1:0] + accbin_in[17][10][4][bW-1:0];
assign sum_out[10][5][bW-1:0] = accbin_in[0][10][5][bW-1:0] + accbin_in[1][10][5][bW-1:0] + accbin_in[2][10][5][bW-1:0] + accbin_in[3][10][5][bW-1:0] + accbin_in[4][10][5][bW-1:0] + accbin_in[5][10][5][bW-1:0] + accbin_in[6][10][5][bW-1:0] + accbin_in[7][10][5][bW-1:0] + accbin_in[8][10][5][bW-1:0] + accbin_in[9][10][5][bW-1:0] + accbin_in[10][10][5][bW-1:0] + accbin_in[11][10][5][bW-1:0] + accbin_in[12][10][5][bW-1:0] + accbin_in[13][10][5][bW-1:0] + accbin_in[14][10][5][bW-1:0] + accbin_in[15][10][5][bW-1:0] + accbin_in[16][10][5][bW-1:0] + accbin_in[17][10][5][bW-1:0];
assign sum_out[10][6][bW-1:0] = accbin_in[0][10][6][bW-1:0] + accbin_in[1][10][6][bW-1:0] + accbin_in[2][10][6][bW-1:0] + accbin_in[3][10][6][bW-1:0] + accbin_in[4][10][6][bW-1:0] + accbin_in[5][10][6][bW-1:0] + accbin_in[6][10][6][bW-1:0] + accbin_in[7][10][6][bW-1:0] + accbin_in[8][10][6][bW-1:0] + accbin_in[9][10][6][bW-1:0] + accbin_in[10][10][6][bW-1:0] + accbin_in[11][10][6][bW-1:0] + accbin_in[12][10][6][bW-1:0] + accbin_in[13][10][6][bW-1:0] + accbin_in[14][10][6][bW-1:0] + accbin_in[15][10][6][bW-1:0] + accbin_in[16][10][6][bW-1:0] + accbin_in[17][10][6][bW-1:0];
assign sum_out[10][7][bW-1:0] = accbin_in[0][10][7][bW-1:0] + accbin_in[1][10][7][bW-1:0] + accbin_in[2][10][7][bW-1:0] + accbin_in[3][10][7][bW-1:0] + accbin_in[4][10][7][bW-1:0] + accbin_in[5][10][7][bW-1:0] + accbin_in[6][10][7][bW-1:0] + accbin_in[7][10][7][bW-1:0] + accbin_in[8][10][7][bW-1:0] + accbin_in[9][10][7][bW-1:0] + accbin_in[10][10][7][bW-1:0] + accbin_in[11][10][7][bW-1:0] + accbin_in[12][10][7][bW-1:0] + accbin_in[13][10][7][bW-1:0] + accbin_in[14][10][7][bW-1:0] + accbin_in[15][10][7][bW-1:0] + accbin_in[16][10][7][bW-1:0] + accbin_in[17][10][7][bW-1:0];
assign sum_out[10][8][bW-1:0] = accbin_in[0][10][8][bW-1:0] + accbin_in[1][10][8][bW-1:0] + accbin_in[2][10][8][bW-1:0] + accbin_in[3][10][8][bW-1:0] + accbin_in[4][10][8][bW-1:0] + accbin_in[5][10][8][bW-1:0] + accbin_in[6][10][8][bW-1:0] + accbin_in[7][10][8][bW-1:0] + accbin_in[8][10][8][bW-1:0] + accbin_in[9][10][8][bW-1:0] + accbin_in[10][10][8][bW-1:0] + accbin_in[11][10][8][bW-1:0] + accbin_in[12][10][8][bW-1:0] + accbin_in[13][10][8][bW-1:0] + accbin_in[14][10][8][bW-1:0] + accbin_in[15][10][8][bW-1:0] + accbin_in[16][10][8][bW-1:0] + accbin_in[17][10][8][bW-1:0];
assign sum_out[10][9][bW-1:0] = accbin_in[0][10][9][bW-1:0] + accbin_in[1][10][9][bW-1:0] + accbin_in[2][10][9][bW-1:0] + accbin_in[3][10][9][bW-1:0] + accbin_in[4][10][9][bW-1:0] + accbin_in[5][10][9][bW-1:0] + accbin_in[6][10][9][bW-1:0] + accbin_in[7][10][9][bW-1:0] + accbin_in[8][10][9][bW-1:0] + accbin_in[9][10][9][bW-1:0] + accbin_in[10][10][9][bW-1:0] + accbin_in[11][10][9][bW-1:0] + accbin_in[12][10][9][bW-1:0] + accbin_in[13][10][9][bW-1:0] + accbin_in[14][10][9][bW-1:0] + accbin_in[15][10][9][bW-1:0] + accbin_in[16][10][9][bW-1:0] + accbin_in[17][10][9][bW-1:0];
assign sum_out[10][10][bW-1:0] = accbin_in[0][10][10][bW-1:0] + accbin_in[1][10][10][bW-1:0] + accbin_in[2][10][10][bW-1:0] + accbin_in[3][10][10][bW-1:0] + accbin_in[4][10][10][bW-1:0] + accbin_in[5][10][10][bW-1:0] + accbin_in[6][10][10][bW-1:0] + accbin_in[7][10][10][bW-1:0] + accbin_in[8][10][10][bW-1:0] + accbin_in[9][10][10][bW-1:0] + accbin_in[10][10][10][bW-1:0] + accbin_in[11][10][10][bW-1:0] + accbin_in[12][10][10][bW-1:0] + accbin_in[13][10][10][bW-1:0] + accbin_in[14][10][10][bW-1:0] + accbin_in[15][10][10][bW-1:0] + accbin_in[16][10][10][bW-1:0] + accbin_in[17][10][10][bW-1:0];
assign sum_out[10][11][bW-1:0] = accbin_in[0][10][11][bW-1:0] + accbin_in[1][10][11][bW-1:0] + accbin_in[2][10][11][bW-1:0] + accbin_in[3][10][11][bW-1:0] + accbin_in[4][10][11][bW-1:0] + accbin_in[5][10][11][bW-1:0] + accbin_in[6][10][11][bW-1:0] + accbin_in[7][10][11][bW-1:0] + accbin_in[8][10][11][bW-1:0] + accbin_in[9][10][11][bW-1:0] + accbin_in[10][10][11][bW-1:0] + accbin_in[11][10][11][bW-1:0] + accbin_in[12][10][11][bW-1:0] + accbin_in[13][10][11][bW-1:0] + accbin_in[14][10][11][bW-1:0] + accbin_in[15][10][11][bW-1:0] + accbin_in[16][10][11][bW-1:0] + accbin_in[17][10][11][bW-1:0];
assign sum_out[11][0][bW-1:0] = accbin_in[0][11][0][bW-1:0] + accbin_in[1][11][0][bW-1:0] + accbin_in[2][11][0][bW-1:0] + accbin_in[3][11][0][bW-1:0] + accbin_in[4][11][0][bW-1:0] + accbin_in[5][11][0][bW-1:0] + accbin_in[6][11][0][bW-1:0] + accbin_in[7][11][0][bW-1:0] + accbin_in[8][11][0][bW-1:0] + accbin_in[9][11][0][bW-1:0] + accbin_in[10][11][0][bW-1:0] + accbin_in[11][11][0][bW-1:0] + accbin_in[12][11][0][bW-1:0] + accbin_in[13][11][0][bW-1:0] + accbin_in[14][11][0][bW-1:0] + accbin_in[15][11][0][bW-1:0] + accbin_in[16][11][0][bW-1:0] + accbin_in[17][11][0][bW-1:0];
assign sum_out[11][1][bW-1:0] = accbin_in[0][11][1][bW-1:0] + accbin_in[1][11][1][bW-1:0] + accbin_in[2][11][1][bW-1:0] + accbin_in[3][11][1][bW-1:0] + accbin_in[4][11][1][bW-1:0] + accbin_in[5][11][1][bW-1:0] + accbin_in[6][11][1][bW-1:0] + accbin_in[7][11][1][bW-1:0] + accbin_in[8][11][1][bW-1:0] + accbin_in[9][11][1][bW-1:0] + accbin_in[10][11][1][bW-1:0] + accbin_in[11][11][1][bW-1:0] + accbin_in[12][11][1][bW-1:0] + accbin_in[13][11][1][bW-1:0] + accbin_in[14][11][1][bW-1:0] + accbin_in[15][11][1][bW-1:0] + accbin_in[16][11][1][bW-1:0] + accbin_in[17][11][1][bW-1:0];
assign sum_out[11][2][bW-1:0] = accbin_in[0][11][2][bW-1:0] + accbin_in[1][11][2][bW-1:0] + accbin_in[2][11][2][bW-1:0] + accbin_in[3][11][2][bW-1:0] + accbin_in[4][11][2][bW-1:0] + accbin_in[5][11][2][bW-1:0] + accbin_in[6][11][2][bW-1:0] + accbin_in[7][11][2][bW-1:0] + accbin_in[8][11][2][bW-1:0] + accbin_in[9][11][2][bW-1:0] + accbin_in[10][11][2][bW-1:0] + accbin_in[11][11][2][bW-1:0] + accbin_in[12][11][2][bW-1:0] + accbin_in[13][11][2][bW-1:0] + accbin_in[14][11][2][bW-1:0] + accbin_in[15][11][2][bW-1:0] + accbin_in[16][11][2][bW-1:0] + accbin_in[17][11][2][bW-1:0];
assign sum_out[11][3][bW-1:0] = accbin_in[0][11][3][bW-1:0] + accbin_in[1][11][3][bW-1:0] + accbin_in[2][11][3][bW-1:0] + accbin_in[3][11][3][bW-1:0] + accbin_in[4][11][3][bW-1:0] + accbin_in[5][11][3][bW-1:0] + accbin_in[6][11][3][bW-1:0] + accbin_in[7][11][3][bW-1:0] + accbin_in[8][11][3][bW-1:0] + accbin_in[9][11][3][bW-1:0] + accbin_in[10][11][3][bW-1:0] + accbin_in[11][11][3][bW-1:0] + accbin_in[12][11][3][bW-1:0] + accbin_in[13][11][3][bW-1:0] + accbin_in[14][11][3][bW-1:0] + accbin_in[15][11][3][bW-1:0] + accbin_in[16][11][3][bW-1:0] + accbin_in[17][11][3][bW-1:0];
assign sum_out[11][4][bW-1:0] = accbin_in[0][11][4][bW-1:0] + accbin_in[1][11][4][bW-1:0] + accbin_in[2][11][4][bW-1:0] + accbin_in[3][11][4][bW-1:0] + accbin_in[4][11][4][bW-1:0] + accbin_in[5][11][4][bW-1:0] + accbin_in[6][11][4][bW-1:0] + accbin_in[7][11][4][bW-1:0] + accbin_in[8][11][4][bW-1:0] + accbin_in[9][11][4][bW-1:0] + accbin_in[10][11][4][bW-1:0] + accbin_in[11][11][4][bW-1:0] + accbin_in[12][11][4][bW-1:0] + accbin_in[13][11][4][bW-1:0] + accbin_in[14][11][4][bW-1:0] + accbin_in[15][11][4][bW-1:0] + accbin_in[16][11][4][bW-1:0] + accbin_in[17][11][4][bW-1:0];
assign sum_out[11][5][bW-1:0] = accbin_in[0][11][5][bW-1:0] + accbin_in[1][11][5][bW-1:0] + accbin_in[2][11][5][bW-1:0] + accbin_in[3][11][5][bW-1:0] + accbin_in[4][11][5][bW-1:0] + accbin_in[5][11][5][bW-1:0] + accbin_in[6][11][5][bW-1:0] + accbin_in[7][11][5][bW-1:0] + accbin_in[8][11][5][bW-1:0] + accbin_in[9][11][5][bW-1:0] + accbin_in[10][11][5][bW-1:0] + accbin_in[11][11][5][bW-1:0] + accbin_in[12][11][5][bW-1:0] + accbin_in[13][11][5][bW-1:0] + accbin_in[14][11][5][bW-1:0] + accbin_in[15][11][5][bW-1:0] + accbin_in[16][11][5][bW-1:0] + accbin_in[17][11][5][bW-1:0];
assign sum_out[11][6][bW-1:0] = accbin_in[0][11][6][bW-1:0] + accbin_in[1][11][6][bW-1:0] + accbin_in[2][11][6][bW-1:0] + accbin_in[3][11][6][bW-1:0] + accbin_in[4][11][6][bW-1:0] + accbin_in[5][11][6][bW-1:0] + accbin_in[6][11][6][bW-1:0] + accbin_in[7][11][6][bW-1:0] + accbin_in[8][11][6][bW-1:0] + accbin_in[9][11][6][bW-1:0] + accbin_in[10][11][6][bW-1:0] + accbin_in[11][11][6][bW-1:0] + accbin_in[12][11][6][bW-1:0] + accbin_in[13][11][6][bW-1:0] + accbin_in[14][11][6][bW-1:0] + accbin_in[15][11][6][bW-1:0] + accbin_in[16][11][6][bW-1:0] + accbin_in[17][11][6][bW-1:0];
assign sum_out[11][7][bW-1:0] = accbin_in[0][11][7][bW-1:0] + accbin_in[1][11][7][bW-1:0] + accbin_in[2][11][7][bW-1:0] + accbin_in[3][11][7][bW-1:0] + accbin_in[4][11][7][bW-1:0] + accbin_in[5][11][7][bW-1:0] + accbin_in[6][11][7][bW-1:0] + accbin_in[7][11][7][bW-1:0] + accbin_in[8][11][7][bW-1:0] + accbin_in[9][11][7][bW-1:0] + accbin_in[10][11][7][bW-1:0] + accbin_in[11][11][7][bW-1:0] + accbin_in[12][11][7][bW-1:0] + accbin_in[13][11][7][bW-1:0] + accbin_in[14][11][7][bW-1:0] + accbin_in[15][11][7][bW-1:0] + accbin_in[16][11][7][bW-1:0] + accbin_in[17][11][7][bW-1:0];
assign sum_out[11][8][bW-1:0] = accbin_in[0][11][8][bW-1:0] + accbin_in[1][11][8][bW-1:0] + accbin_in[2][11][8][bW-1:0] + accbin_in[3][11][8][bW-1:0] + accbin_in[4][11][8][bW-1:0] + accbin_in[5][11][8][bW-1:0] + accbin_in[6][11][8][bW-1:0] + accbin_in[7][11][8][bW-1:0] + accbin_in[8][11][8][bW-1:0] + accbin_in[9][11][8][bW-1:0] + accbin_in[10][11][8][bW-1:0] + accbin_in[11][11][8][bW-1:0] + accbin_in[12][11][8][bW-1:0] + accbin_in[13][11][8][bW-1:0] + accbin_in[14][11][8][bW-1:0] + accbin_in[15][11][8][bW-1:0] + accbin_in[16][11][8][bW-1:0] + accbin_in[17][11][8][bW-1:0];
assign sum_out[11][9][bW-1:0] = accbin_in[0][11][9][bW-1:0] + accbin_in[1][11][9][bW-1:0] + accbin_in[2][11][9][bW-1:0] + accbin_in[3][11][9][bW-1:0] + accbin_in[4][11][9][bW-1:0] + accbin_in[5][11][9][bW-1:0] + accbin_in[6][11][9][bW-1:0] + accbin_in[7][11][9][bW-1:0] + accbin_in[8][11][9][bW-1:0] + accbin_in[9][11][9][bW-1:0] + accbin_in[10][11][9][bW-1:0] + accbin_in[11][11][9][bW-1:0] + accbin_in[12][11][9][bW-1:0] + accbin_in[13][11][9][bW-1:0] + accbin_in[14][11][9][bW-1:0] + accbin_in[15][11][9][bW-1:0] + accbin_in[16][11][9][bW-1:0] + accbin_in[17][11][9][bW-1:0];
assign sum_out[11][10][bW-1:0] = accbin_in[0][11][10][bW-1:0] + accbin_in[1][11][10][bW-1:0] + accbin_in[2][11][10][bW-1:0] + accbin_in[3][11][10][bW-1:0] + accbin_in[4][11][10][bW-1:0] + accbin_in[5][11][10][bW-1:0] + accbin_in[6][11][10][bW-1:0] + accbin_in[7][11][10][bW-1:0] + accbin_in[8][11][10][bW-1:0] + accbin_in[9][11][10][bW-1:0] + accbin_in[10][11][10][bW-1:0] + accbin_in[11][11][10][bW-1:0] + accbin_in[12][11][10][bW-1:0] + accbin_in[13][11][10][bW-1:0] + accbin_in[14][11][10][bW-1:0] + accbin_in[15][11][10][bW-1:0] + accbin_in[16][11][10][bW-1:0] + accbin_in[17][11][10][bW-1:0];
assign sum_out[11][11][bW-1:0] = accbin_in[0][11][11][bW-1:0] + accbin_in[1][11][11][bW-1:0] + accbin_in[2][11][11][bW-1:0] + accbin_in[3][11][11][bW-1:0] + accbin_in[4][11][11][bW-1:0] + accbin_in[5][11][11][bW-1:0] + accbin_in[6][11][11][bW-1:0] + accbin_in[7][11][11][bW-1:0] + accbin_in[8][11][11][bW-1:0] + accbin_in[9][11][11][bW-1:0] + accbin_in[10][11][11][bW-1:0] + accbin_in[11][11][11][bW-1:0] + accbin_in[12][11][11][bW-1:0] + accbin_in[13][11][11][bW-1:0] + accbin_in[14][11][11][bW-1:0] + accbin_in[15][11][11][bW-1:0] + accbin_in[16][11][11][bW-1:0] + accbin_in[17][11][11][bW-1:0];

assign accbin_out[0][0] = (sum_out[0][0][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[0][1] = (sum_out[0][1][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[0][2] = (sum_out[0][2][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[0][3] = (sum_out[0][3][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[0][4] = (sum_out[0][4][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[0][5] = (sum_out[0][5][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[0][6] = (sum_out[0][6][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[0][7] = (sum_out[0][7][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[0][8] = (sum_out[0][8][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[0][9] = (sum_out[0][9][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[0][10] = (sum_out[0][10][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[0][11] = (sum_out[0][11][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[1][0] = (sum_out[1][0][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[1][1] = (sum_out[1][1][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[1][2] = (sum_out[1][2][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[1][3] = (sum_out[1][3][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[1][4] = (sum_out[1][4][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[1][5] = (sum_out[1][5][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[1][6] = (sum_out[1][6][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[1][7] = (sum_out[1][7][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[1][8] = (sum_out[1][8][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[1][9] = (sum_out[1][9][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[1][10] = (sum_out[1][10][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[1][11] = (sum_out[1][11][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[2][0] = (sum_out[2][0][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[2][1] = (sum_out[2][1][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[2][2] = (sum_out[2][2][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[2][3] = (sum_out[2][3][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[2][4] = (sum_out[2][4][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[2][5] = (sum_out[2][5][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[2][6] = (sum_out[2][6][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[2][7] = (sum_out[2][7][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[2][8] = (sum_out[2][8][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[2][9] = (sum_out[2][9][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[2][10] = (sum_out[2][10][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[2][11] = (sum_out[2][11][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[3][0] = (sum_out[3][0][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[3][1] = (sum_out[3][1][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[3][2] = (sum_out[3][2][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[3][3] = (sum_out[3][3][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[3][4] = (sum_out[3][4][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[3][5] = (sum_out[3][5][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[3][6] = (sum_out[3][6][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[3][7] = (sum_out[3][7][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[3][8] = (sum_out[3][8][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[3][9] = (sum_out[3][9][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[3][10] = (sum_out[3][10][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[3][11] = (sum_out[3][11][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[4][0] = (sum_out[4][0][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[4][1] = (sum_out[4][1][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[4][2] = (sum_out[4][2][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[4][3] = (sum_out[4][3][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[4][4] = (sum_out[4][4][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[4][5] = (sum_out[4][5][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[4][6] = (sum_out[4][6][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[4][7] = (sum_out[4][7][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[4][8] = (sum_out[4][8][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[4][9] = (sum_out[4][9][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[4][10] = (sum_out[4][10][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[4][11] = (sum_out[4][11][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[5][0] = (sum_out[5][0][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[5][1] = (sum_out[5][1][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[5][2] = (sum_out[5][2][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[5][3] = (sum_out[5][3][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[5][4] = (sum_out[5][4][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[5][5] = (sum_out[5][5][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[5][6] = (sum_out[5][6][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[5][7] = (sum_out[5][7][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[5][8] = (sum_out[5][8][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[5][9] = (sum_out[5][9][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[5][10] = (sum_out[5][10][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[5][11] = (sum_out[5][11][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[6][0] = (sum_out[6][0][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[6][1] = (sum_out[6][1][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[6][2] = (sum_out[6][2][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[6][3] = (sum_out[6][3][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[6][4] = (sum_out[6][4][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[6][5] = (sum_out[6][5][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[6][6] = (sum_out[6][6][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[6][7] = (sum_out[6][7][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[6][8] = (sum_out[6][8][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[6][9] = (sum_out[6][9][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[6][10] = (sum_out[6][10][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[6][11] = (sum_out[6][11][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[7][0] = (sum_out[7][0][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[7][1] = (sum_out[7][1][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[7][2] = (sum_out[7][2][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[7][3] = (sum_out[7][3][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[7][4] = (sum_out[7][4][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[7][5] = (sum_out[7][5][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[7][6] = (sum_out[7][6][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[7][7] = (sum_out[7][7][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[7][8] = (sum_out[7][8][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[7][9] = (sum_out[7][9][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[7][10] = (sum_out[7][10][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[7][11] = (sum_out[7][11][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[8][0] = (sum_out[8][0][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[8][1] = (sum_out[8][1][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[8][2] = (sum_out[8][2][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[8][3] = (sum_out[8][3][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[8][4] = (sum_out[8][4][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[8][5] = (sum_out[8][5][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[8][6] = (sum_out[8][6][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[8][7] = (sum_out[8][7][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[8][8] = (sum_out[8][8][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[8][9] = (sum_out[8][9][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[8][10] = (sum_out[8][10][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[8][11] = (sum_out[8][11][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[9][0] = (sum_out[9][0][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[9][1] = (sum_out[9][1][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[9][2] = (sum_out[9][2][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[9][3] = (sum_out[9][3][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[9][4] = (sum_out[9][4][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[9][5] = (sum_out[9][5][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[9][6] = (sum_out[9][6][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[9][7] = (sum_out[9][7][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[9][8] = (sum_out[9][8][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[9][9] = (sum_out[9][9][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[9][10] = (sum_out[9][10][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[9][11] = (sum_out[9][11][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[10][0] = (sum_out[10][0][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[10][1] = (sum_out[10][1][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[10][2] = (sum_out[10][2][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[10][3] = (sum_out[10][3][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[10][4] = (sum_out[10][4][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[10][5] = (sum_out[10][5][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[10][6] = (sum_out[10][6][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[10][7] = (sum_out[10][7][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[10][8] = (sum_out[10][8][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[10][9] = (sum_out[10][9][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[10][10] = (sum_out[10][10][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[10][11] = (sum_out[10][11][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[11][0] = (sum_out[11][0][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[11][1] = (sum_out[11][1][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[11][2] = (sum_out[11][2][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[11][3] = (sum_out[11][3][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[11][4] = (sum_out[11][4][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[11][5] = (sum_out[11][5][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[11][6] = (sum_out[11][6][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[11][7] = (sum_out[11][7][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[11][8] = (sum_out[11][8][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[11][9] = (sum_out[11][9][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[11][10] = (sum_out[11][10][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;
assign accbin_out[11][11] = (sum_out[11][11][bW-1:0] > kernel_offset[bW-1:0]) ? 1'b1 : 1'b0;

endmodule