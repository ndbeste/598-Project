module convchan2( 
    input  logic signed image     [0:11][0:11],
    input  logic        kernel    [0:4] [0:4],
    output logic        out_fmap  [0:7][0:7]
    );

logic signed [bW-1:0] xor_sum       [0:7][0:7];
logic signed [1   :0] signed_kernel [0:4][0:4];


// Make kernel signed 

always_ff @(posedge clk) begin
    if(~rst_n) begin
        for(i=0; i<5; i=i+1) begin
            for(j=0; j<5; j=j+1) begin
                signed_kernel[i][j] <= 2'b00;
            end
        end
    end else begin
        for(i=0; i<5; i=i+1) begin
            for(j=0; j<5; j=j+1) begin
                signed_kernel[i][j] <= (kernel[i][j] == 1'b1) ? 2'b01 : 2'b11;
            end
        end
    end
end

assign xor_sum[0][0] = kernel[0][0] ~^ image[0][0] + kernel[0][1] ~^ image[0][1] + kernel[0][2] ~^ image[0][2] + kernel[0][3] ~^ image[0][3] + kernel[0][4] ~^ image[0][4] + kernel[1][0] ~^ image[1][0] + kernel[1][1] ~^ image[1][1] + kernel[1][2] ~^ image[1][2] + kernel[1][3] ~^ image[1][3] + kernel[1][4] ~^ image[1][4] + kernel[2][0] ~^ image[2][0] + kernel[2][1] ~^ image[2][1] + kernel[2][2] ~^ image[2][2] + kernel[2][3] ~^ image[2][3] + kernel[2][4] ~^ image[2][4] + kernel[3][0] ~^ image[3][0] + kernel[3][1] ~^ image[3][1] + kernel[3][2] ~^ image[3][2] + kernel[3][3] ~^ image[3][3] + kernel[3][4] ~^ image[3][4] + kernel[4][0] ~^ image[4][0] + kernel[4][1] ~^ image[4][1] + kernel[4][2] ~^ image[4][2] + kernel[4][3] ~^ image[4][3] + kernel[4][4] ~^ image[4][4];
assign xor_sum[0][1] = kernel[0][0] ~^ image[0][1] + kernel[0][1] ~^ image[0][2] + kernel[0][2] ~^ image[0][3] + kernel[0][3] ~^ image[0][4] + kernel[0][4] ~^ image[0][5] + kernel[1][0] ~^ image[1][1] + kernel[1][1] ~^ image[1][2] + kernel[1][2] ~^ image[1][3] + kernel[1][3] ~^ image[1][4] + kernel[1][4] ~^ image[1][5] + kernel[2][0] ~^ image[2][1] + kernel[2][1] ~^ image[2][2] + kernel[2][2] ~^ image[2][3] + kernel[2][3] ~^ image[2][4] + kernel[2][4] ~^ image[2][5] + kernel[3][0] ~^ image[3][1] + kernel[3][1] ~^ image[3][2] + kernel[3][2] ~^ image[3][3] + kernel[3][3] ~^ image[3][4] + kernel[3][4] ~^ image[3][5] + kernel[4][0] ~^ image[4][1] + kernel[4][1] ~^ image[4][2] + kernel[4][2] ~^ image[4][3] + kernel[4][3] ~^ image[4][4] + kernel[4][4] ~^ image[4][5];
assign xor_sum[0][2] = kernel[0][0] ~^ image[0][2] + kernel[0][1] ~^ image[0][3] + kernel[0][2] ~^ image[0][4] + kernel[0][3] ~^ image[0][5] + kernel[0][4] ~^ image[0][6] + kernel[1][0] ~^ image[1][2] + kernel[1][1] ~^ image[1][3] + kernel[1][2] ~^ image[1][4] + kernel[1][3] ~^ image[1][5] + kernel[1][4] ~^ image[1][6] + kernel[2][0] ~^ image[2][2] + kernel[2][1] ~^ image[2][3] + kernel[2][2] ~^ image[2][4] + kernel[2][3] ~^ image[2][5] + kernel[2][4] ~^ image[2][6] + kernel[3][0] ~^ image[3][2] + kernel[3][1] ~^ image[3][3] + kernel[3][2] ~^ image[3][4] + kernel[3][3] ~^ image[3][5] + kernel[3][4] ~^ image[3][6] + kernel[4][0] ~^ image[4][2] + kernel[4][1] ~^ image[4][3] + kernel[4][2] ~^ image[4][4] + kernel[4][3] ~^ image[4][5] + kernel[4][4] ~^ image[4][6];
assign xor_sum[0][3] = kernel[0][0] ~^ image[0][3] + kernel[0][1] ~^ image[0][4] + kernel[0][2] ~^ image[0][5] + kernel[0][3] ~^ image[0][6] + kernel[0][4] ~^ image[0][7] + kernel[1][0] ~^ image[1][3] + kernel[1][1] ~^ image[1][4] + kernel[1][2] ~^ image[1][5] + kernel[1][3] ~^ image[1][6] + kernel[1][4] ~^ image[1][7] + kernel[2][0] ~^ image[2][3] + kernel[2][1] ~^ image[2][4] + kernel[2][2] ~^ image[2][5] + kernel[2][3] ~^ image[2][6] + kernel[2][4] ~^ image[2][7] + kernel[3][0] ~^ image[3][3] + kernel[3][1] ~^ image[3][4] + kernel[3][2] ~^ image[3][5] + kernel[3][3] ~^ image[3][6] + kernel[3][4] ~^ image[3][7] + kernel[4][0] ~^ image[4][3] + kernel[4][1] ~^ image[4][4] + kernel[4][2] ~^ image[4][5] + kernel[4][3] ~^ image[4][6] + kernel[4][4] ~^ image[4][7];
assign xor_sum[0][4] = kernel[0][0] ~^ image[0][4] + kernel[0][1] ~^ image[0][5] + kernel[0][2] ~^ image[0][6] + kernel[0][3] ~^ image[0][7] + kernel[0][4] ~^ image[0][8] + kernel[1][0] ~^ image[1][4] + kernel[1][1] ~^ image[1][5] + kernel[1][2] ~^ image[1][6] + kernel[1][3] ~^ image[1][7] + kernel[1][4] ~^ image[1][8] + kernel[2][0] ~^ image[2][4] + kernel[2][1] ~^ image[2][5] + kernel[2][2] ~^ image[2][6] + kernel[2][3] ~^ image[2][7] + kernel[2][4] ~^ image[2][8] + kernel[3][0] ~^ image[3][4] + kernel[3][1] ~^ image[3][5] + kernel[3][2] ~^ image[3][6] + kernel[3][3] ~^ image[3][7] + kernel[3][4] ~^ image[3][8] + kernel[4][0] ~^ image[4][4] + kernel[4][1] ~^ image[4][5] + kernel[4][2] ~^ image[4][6] + kernel[4][3] ~^ image[4][7] + kernel[4][4] ~^ image[4][8];
assign xor_sum[0][5] = kernel[0][0] ~^ image[0][5] + kernel[0][1] ~^ image[0][6] + kernel[0][2] ~^ image[0][7] + kernel[0][3] ~^ image[0][8] + kernel[0][4] ~^ image[0][9] + kernel[1][0] ~^ image[1][5] + kernel[1][1] ~^ image[1][6] + kernel[1][2] ~^ image[1][7] + kernel[1][3] ~^ image[1][8] + kernel[1][4] ~^ image[1][9] + kernel[2][0] ~^ image[2][5] + kernel[2][1] ~^ image[2][6] + kernel[2][2] ~^ image[2][7] + kernel[2][3] ~^ image[2][8] + kernel[2][4] ~^ image[2][9] + kernel[3][0] ~^ image[3][5] + kernel[3][1] ~^ image[3][6] + kernel[3][2] ~^ image[3][7] + kernel[3][3] ~^ image[3][8] + kernel[3][4] ~^ image[3][9] + kernel[4][0] ~^ image[4][5] + kernel[4][1] ~^ image[4][6] + kernel[4][2] ~^ image[4][7] + kernel[4][3] ~^ image[4][8] + kernel[4][4] ~^ image[4][9];
assign xor_sum[0][6] = kernel[0][0] ~^ image[0][6] + kernel[0][1] ~^ image[0][7] + kernel[0][2] ~^ image[0][8] + kernel[0][3] ~^ image[0][9] + kernel[0][4] ~^ image[0][10] + kernel[1][0] ~^ image[1][6] + kernel[1][1] ~^ image[1][7] + kernel[1][2] ~^ image[1][8] + kernel[1][3] ~^ image[1][9] + kernel[1][4] ~^ image[1][10] + kernel[2][0] ~^ image[2][6] + kernel[2][1] ~^ image[2][7] + kernel[2][2] ~^ image[2][8] + kernel[2][3] ~^ image[2][9] + kernel[2][4] ~^ image[2][10] + kernel[3][0] ~^ image[3][6] + kernel[3][1] ~^ image[3][7] + kernel[3][2] ~^ image[3][8] + kernel[3][3] ~^ image[3][9] + kernel[3][4] ~^ image[3][10] + kernel[4][0] ~^ image[4][6] + kernel[4][1] ~^ image[4][7] + kernel[4][2] ~^ image[4][8] + kernel[4][3] ~^ image[4][9] + kernel[4][4] ~^ image[4][10];
assign xor_sum[0][7] = kernel[0][0] ~^ image[0][7] + kernel[0][1] ~^ image[0][8] + kernel[0][2] ~^ image[0][9] + kernel[0][3] ~^ image[0][10] + kernel[0][4] ~^ image[0][11] + kernel[1][0] ~^ image[1][7] + kernel[1][1] ~^ image[1][8] + kernel[1][2] ~^ image[1][9] + kernel[1][3] ~^ image[1][10] + kernel[1][4] ~^ image[1][11] + kernel[2][0] ~^ image[2][7] + kernel[2][1] ~^ image[2][8] + kernel[2][2] ~^ image[2][9] + kernel[2][3] ~^ image[2][10] + kernel[2][4] ~^ image[2][11] + kernel[3][0] ~^ image[3][7] + kernel[3][1] ~^ image[3][8] + kernel[3][2] ~^ image[3][9] + kernel[3][3] ~^ image[3][10] + kernel[3][4] ~^ image[3][11] + kernel[4][0] ~^ image[4][7] + kernel[4][1] ~^ image[4][8] + kernel[4][2] ~^ image[4][9] + kernel[4][3] ~^ image[4][10] + kernel[4][4] ~^ image[4][11];
assign xor_sum[1][0] = kernel[0][0] ~^ image[1][0] + kernel[0][1] ~^ image[1][1] + kernel[0][2] ~^ image[1][2] + kernel[0][3] ~^ image[1][3] + kernel[0][4] ~^ image[1][4] + kernel[1][0] ~^ image[2][0] + kernel[1][1] ~^ image[2][1] + kernel[1][2] ~^ image[2][2] + kernel[1][3] ~^ image[2][3] + kernel[1][4] ~^ image[2][4] + kernel[2][0] ~^ image[3][0] + kernel[2][1] ~^ image[3][1] + kernel[2][2] ~^ image[3][2] + kernel[2][3] ~^ image[3][3] + kernel[2][4] ~^ image[3][4] + kernel[3][0] ~^ image[4][0] + kernel[3][1] ~^ image[4][1] + kernel[3][2] ~^ image[4][2] + kernel[3][3] ~^ image[4][3] + kernel[3][4] ~^ image[4][4] + kernel[4][0] ~^ image[5][0] + kernel[4][1] ~^ image[5][1] + kernel[4][2] ~^ image[5][2] + kernel[4][3] ~^ image[5][3] + kernel[4][4] ~^ image[5][4];
assign xor_sum[1][1] = kernel[0][0] ~^ image[1][1] + kernel[0][1] ~^ image[1][2] + kernel[0][2] ~^ image[1][3] + kernel[0][3] ~^ image[1][4] + kernel[0][4] ~^ image[1][5] + kernel[1][0] ~^ image[2][1] + kernel[1][1] ~^ image[2][2] + kernel[1][2] ~^ image[2][3] + kernel[1][3] ~^ image[2][4] + kernel[1][4] ~^ image[2][5] + kernel[2][0] ~^ image[3][1] + kernel[2][1] ~^ image[3][2] + kernel[2][2] ~^ image[3][3] + kernel[2][3] ~^ image[3][4] + kernel[2][4] ~^ image[3][5] + kernel[3][0] ~^ image[4][1] + kernel[3][1] ~^ image[4][2] + kernel[3][2] ~^ image[4][3] + kernel[3][3] ~^ image[4][4] + kernel[3][4] ~^ image[4][5] + kernel[4][0] ~^ image[5][1] + kernel[4][1] ~^ image[5][2] + kernel[4][2] ~^ image[5][3] + kernel[4][3] ~^ image[5][4] + kernel[4][4] ~^ image[5][5];
assign xor_sum[1][2] = kernel[0][0] ~^ image[1][2] + kernel[0][1] ~^ image[1][3] + kernel[0][2] ~^ image[1][4] + kernel[0][3] ~^ image[1][5] + kernel[0][4] ~^ image[1][6] + kernel[1][0] ~^ image[2][2] + kernel[1][1] ~^ image[2][3] + kernel[1][2] ~^ image[2][4] + kernel[1][3] ~^ image[2][5] + kernel[1][4] ~^ image[2][6] + kernel[2][0] ~^ image[3][2] + kernel[2][1] ~^ image[3][3] + kernel[2][2] ~^ image[3][4] + kernel[2][3] ~^ image[3][5] + kernel[2][4] ~^ image[3][6] + kernel[3][0] ~^ image[4][2] + kernel[3][1] ~^ image[4][3] + kernel[3][2] ~^ image[4][4] + kernel[3][3] ~^ image[4][5] + kernel[3][4] ~^ image[4][6] + kernel[4][0] ~^ image[5][2] + kernel[4][1] ~^ image[5][3] + kernel[4][2] ~^ image[5][4] + kernel[4][3] ~^ image[5][5] + kernel[4][4] ~^ image[5][6];
assign xor_sum[1][3] = kernel[0][0] ~^ image[1][3] + kernel[0][1] ~^ image[1][4] + kernel[0][2] ~^ image[1][5] + kernel[0][3] ~^ image[1][6] + kernel[0][4] ~^ image[1][7] + kernel[1][0] ~^ image[2][3] + kernel[1][1] ~^ image[2][4] + kernel[1][2] ~^ image[2][5] + kernel[1][3] ~^ image[2][6] + kernel[1][4] ~^ image[2][7] + kernel[2][0] ~^ image[3][3] + kernel[2][1] ~^ image[3][4] + kernel[2][2] ~^ image[3][5] + kernel[2][3] ~^ image[3][6] + kernel[2][4] ~^ image[3][7] + kernel[3][0] ~^ image[4][3] + kernel[3][1] ~^ image[4][4] + kernel[3][2] ~^ image[4][5] + kernel[3][3] ~^ image[4][6] + kernel[3][4] ~^ image[4][7] + kernel[4][0] ~^ image[5][3] + kernel[4][1] ~^ image[5][4] + kernel[4][2] ~^ image[5][5] + kernel[4][3] ~^ image[5][6] + kernel[4][4] ~^ image[5][7];
assign xor_sum[1][4] = kernel[0][0] ~^ image[1][4] + kernel[0][1] ~^ image[1][5] + kernel[0][2] ~^ image[1][6] + kernel[0][3] ~^ image[1][7] + kernel[0][4] ~^ image[1][8] + kernel[1][0] ~^ image[2][4] + kernel[1][1] ~^ image[2][5] + kernel[1][2] ~^ image[2][6] + kernel[1][3] ~^ image[2][7] + kernel[1][4] ~^ image[2][8] + kernel[2][0] ~^ image[3][4] + kernel[2][1] ~^ image[3][5] + kernel[2][2] ~^ image[3][6] + kernel[2][3] ~^ image[3][7] + kernel[2][4] ~^ image[3][8] + kernel[3][0] ~^ image[4][4] + kernel[3][1] ~^ image[4][5] + kernel[3][2] ~^ image[4][6] + kernel[3][3] ~^ image[4][7] + kernel[3][4] ~^ image[4][8] + kernel[4][0] ~^ image[5][4] + kernel[4][1] ~^ image[5][5] + kernel[4][2] ~^ image[5][6] + kernel[4][3] ~^ image[5][7] + kernel[4][4] ~^ image[5][8];
assign xor_sum[1][5] = kernel[0][0] ~^ image[1][5] + kernel[0][1] ~^ image[1][6] + kernel[0][2] ~^ image[1][7] + kernel[0][3] ~^ image[1][8] + kernel[0][4] ~^ image[1][9] + kernel[1][0] ~^ image[2][5] + kernel[1][1] ~^ image[2][6] + kernel[1][2] ~^ image[2][7] + kernel[1][3] ~^ image[2][8] + kernel[1][4] ~^ image[2][9] + kernel[2][0] ~^ image[3][5] + kernel[2][1] ~^ image[3][6] + kernel[2][2] ~^ image[3][7] + kernel[2][3] ~^ image[3][8] + kernel[2][4] ~^ image[3][9] + kernel[3][0] ~^ image[4][5] + kernel[3][1] ~^ image[4][6] + kernel[3][2] ~^ image[4][7] + kernel[3][3] ~^ image[4][8] + kernel[3][4] ~^ image[4][9] + kernel[4][0] ~^ image[5][5] + kernel[4][1] ~^ image[5][6] + kernel[4][2] ~^ image[5][7] + kernel[4][3] ~^ image[5][8] + kernel[4][4] ~^ image[5][9];
assign xor_sum[1][6] = kernel[0][0] ~^ image[1][6] + kernel[0][1] ~^ image[1][7] + kernel[0][2] ~^ image[1][8] + kernel[0][3] ~^ image[1][9] + kernel[0][4] ~^ image[1][10] + kernel[1][0] ~^ image[2][6] + kernel[1][1] ~^ image[2][7] + kernel[1][2] ~^ image[2][8] + kernel[1][3] ~^ image[2][9] + kernel[1][4] ~^ image[2][10] + kernel[2][0] ~^ image[3][6] + kernel[2][1] ~^ image[3][7] + kernel[2][2] ~^ image[3][8] + kernel[2][3] ~^ image[3][9] + kernel[2][4] ~^ image[3][10] + kernel[3][0] ~^ image[4][6] + kernel[3][1] ~^ image[4][7] + kernel[3][2] ~^ image[4][8] + kernel[3][3] ~^ image[4][9] + kernel[3][4] ~^ image[4][10] + kernel[4][0] ~^ image[5][6] + kernel[4][1] ~^ image[5][7] + kernel[4][2] ~^ image[5][8] + kernel[4][3] ~^ image[5][9] + kernel[4][4] ~^ image[5][10];
assign xor_sum[1][7] = kernel[0][0] ~^ image[1][7] + kernel[0][1] ~^ image[1][8] + kernel[0][2] ~^ image[1][9] + kernel[0][3] ~^ image[1][10] + kernel[0][4] ~^ image[1][11] + kernel[1][0] ~^ image[2][7] + kernel[1][1] ~^ image[2][8] + kernel[1][2] ~^ image[2][9] + kernel[1][3] ~^ image[2][10] + kernel[1][4] ~^ image[2][11] + kernel[2][0] ~^ image[3][7] + kernel[2][1] ~^ image[3][8] + kernel[2][2] ~^ image[3][9] + kernel[2][3] ~^ image[3][10] + kernel[2][4] ~^ image[3][11] + kernel[3][0] ~^ image[4][7] + kernel[3][1] ~^ image[4][8] + kernel[3][2] ~^ image[4][9] + kernel[3][3] ~^ image[4][10] + kernel[3][4] ~^ image[4][11] + kernel[4][0] ~^ image[5][7] + kernel[4][1] ~^ image[5][8] + kernel[4][2] ~^ image[5][9] + kernel[4][3] ~^ image[5][10] + kernel[4][4] ~^ image[5][11];
assign xor_sum[2][0] = kernel[0][0] ~^ image[2][0] + kernel[0][1] ~^ image[2][1] + kernel[0][2] ~^ image[2][2] + kernel[0][3] ~^ image[2][3] + kernel[0][4] ~^ image[2][4] + kernel[1][0] ~^ image[3][0] + kernel[1][1] ~^ image[3][1] + kernel[1][2] ~^ image[3][2] + kernel[1][3] ~^ image[3][3] + kernel[1][4] ~^ image[3][4] + kernel[2][0] ~^ image[4][0] + kernel[2][1] ~^ image[4][1] + kernel[2][2] ~^ image[4][2] + kernel[2][3] ~^ image[4][3] + kernel[2][4] ~^ image[4][4] + kernel[3][0] ~^ image[5][0] + kernel[3][1] ~^ image[5][1] + kernel[3][2] ~^ image[5][2] + kernel[3][3] ~^ image[5][3] + kernel[3][4] ~^ image[5][4] + kernel[4][0] ~^ image[6][0] + kernel[4][1] ~^ image[6][1] + kernel[4][2] ~^ image[6][2] + kernel[4][3] ~^ image[6][3] + kernel[4][4] ~^ image[6][4];
assign xor_sum[2][1] = kernel[0][0] ~^ image[2][1] + kernel[0][1] ~^ image[2][2] + kernel[0][2] ~^ image[2][3] + kernel[0][3] ~^ image[2][4] + kernel[0][4] ~^ image[2][5] + kernel[1][0] ~^ image[3][1] + kernel[1][1] ~^ image[3][2] + kernel[1][2] ~^ image[3][3] + kernel[1][3] ~^ image[3][4] + kernel[1][4] ~^ image[3][5] + kernel[2][0] ~^ image[4][1] + kernel[2][1] ~^ image[4][2] + kernel[2][2] ~^ image[4][3] + kernel[2][3] ~^ image[4][4] + kernel[2][4] ~^ image[4][5] + kernel[3][0] ~^ image[5][1] + kernel[3][1] ~^ image[5][2] + kernel[3][2] ~^ image[5][3] + kernel[3][3] ~^ image[5][4] + kernel[3][4] ~^ image[5][5] + kernel[4][0] ~^ image[6][1] + kernel[4][1] ~^ image[6][2] + kernel[4][2] ~^ image[6][3] + kernel[4][3] ~^ image[6][4] + kernel[4][4] ~^ image[6][5];
assign xor_sum[2][2] = kernel[0][0] ~^ image[2][2] + kernel[0][1] ~^ image[2][3] + kernel[0][2] ~^ image[2][4] + kernel[0][3] ~^ image[2][5] + kernel[0][4] ~^ image[2][6] + kernel[1][0] ~^ image[3][2] + kernel[1][1] ~^ image[3][3] + kernel[1][2] ~^ image[3][4] + kernel[1][3] ~^ image[3][5] + kernel[1][4] ~^ image[3][6] + kernel[2][0] ~^ image[4][2] + kernel[2][1] ~^ image[4][3] + kernel[2][2] ~^ image[4][4] + kernel[2][3] ~^ image[4][5] + kernel[2][4] ~^ image[4][6] + kernel[3][0] ~^ image[5][2] + kernel[3][1] ~^ image[5][3] + kernel[3][2] ~^ image[5][4] + kernel[3][3] ~^ image[5][5] + kernel[3][4] ~^ image[5][6] + kernel[4][0] ~^ image[6][2] + kernel[4][1] ~^ image[6][3] + kernel[4][2] ~^ image[6][4] + kernel[4][3] ~^ image[6][5] + kernel[4][4] ~^ image[6][6];
assign xor_sum[2][3] = kernel[0][0] ~^ image[2][3] + kernel[0][1] ~^ image[2][4] + kernel[0][2] ~^ image[2][5] + kernel[0][3] ~^ image[2][6] + kernel[0][4] ~^ image[2][7] + kernel[1][0] ~^ image[3][3] + kernel[1][1] ~^ image[3][4] + kernel[1][2] ~^ image[3][5] + kernel[1][3] ~^ image[3][6] + kernel[1][4] ~^ image[3][7] + kernel[2][0] ~^ image[4][3] + kernel[2][1] ~^ image[4][4] + kernel[2][2] ~^ image[4][5] + kernel[2][3] ~^ image[4][6] + kernel[2][4] ~^ image[4][7] + kernel[3][0] ~^ image[5][3] + kernel[3][1] ~^ image[5][4] + kernel[3][2] ~^ image[5][5] + kernel[3][3] ~^ image[5][6] + kernel[3][4] ~^ image[5][7] + kernel[4][0] ~^ image[6][3] + kernel[4][1] ~^ image[6][4] + kernel[4][2] ~^ image[6][5] + kernel[4][3] ~^ image[6][6] + kernel[4][4] ~^ image[6][7];
assign xor_sum[2][4] = kernel[0][0] ~^ image[2][4] + kernel[0][1] ~^ image[2][5] + kernel[0][2] ~^ image[2][6] + kernel[0][3] ~^ image[2][7] + kernel[0][4] ~^ image[2][8] + kernel[1][0] ~^ image[3][4] + kernel[1][1] ~^ image[3][5] + kernel[1][2] ~^ image[3][6] + kernel[1][3] ~^ image[3][7] + kernel[1][4] ~^ image[3][8] + kernel[2][0] ~^ image[4][4] + kernel[2][1] ~^ image[4][5] + kernel[2][2] ~^ image[4][6] + kernel[2][3] ~^ image[4][7] + kernel[2][4] ~^ image[4][8] + kernel[3][0] ~^ image[5][4] + kernel[3][1] ~^ image[5][5] + kernel[3][2] ~^ image[5][6] + kernel[3][3] ~^ image[5][7] + kernel[3][4] ~^ image[5][8] + kernel[4][0] ~^ image[6][4] + kernel[4][1] ~^ image[6][5] + kernel[4][2] ~^ image[6][6] + kernel[4][3] ~^ image[6][7] + kernel[4][4] ~^ image[6][8];
assign xor_sum[2][5] = kernel[0][0] ~^ image[2][5] + kernel[0][1] ~^ image[2][6] + kernel[0][2] ~^ image[2][7] + kernel[0][3] ~^ image[2][8] + kernel[0][4] ~^ image[2][9] + kernel[1][0] ~^ image[3][5] + kernel[1][1] ~^ image[3][6] + kernel[1][2] ~^ image[3][7] + kernel[1][3] ~^ image[3][8] + kernel[1][4] ~^ image[3][9] + kernel[2][0] ~^ image[4][5] + kernel[2][1] ~^ image[4][6] + kernel[2][2] ~^ image[4][7] + kernel[2][3] ~^ image[4][8] + kernel[2][4] ~^ image[4][9] + kernel[3][0] ~^ image[5][5] + kernel[3][1] ~^ image[5][6] + kernel[3][2] ~^ image[5][7] + kernel[3][3] ~^ image[5][8] + kernel[3][4] ~^ image[5][9] + kernel[4][0] ~^ image[6][5] + kernel[4][1] ~^ image[6][6] + kernel[4][2] ~^ image[6][7] + kernel[4][3] ~^ image[6][8] + kernel[4][4] ~^ image[6][9];
assign xor_sum[2][6] = kernel[0][0] ~^ image[2][6] + kernel[0][1] ~^ image[2][7] + kernel[0][2] ~^ image[2][8] + kernel[0][3] ~^ image[2][9] + kernel[0][4] ~^ image[2][10] + kernel[1][0] ~^ image[3][6] + kernel[1][1] ~^ image[3][7] + kernel[1][2] ~^ image[3][8] + kernel[1][3] ~^ image[3][9] + kernel[1][4] ~^ image[3][10] + kernel[2][0] ~^ image[4][6] + kernel[2][1] ~^ image[4][7] + kernel[2][2] ~^ image[4][8] + kernel[2][3] ~^ image[4][9] + kernel[2][4] ~^ image[4][10] + kernel[3][0] ~^ image[5][6] + kernel[3][1] ~^ image[5][7] + kernel[3][2] ~^ image[5][8] + kernel[3][3] ~^ image[5][9] + kernel[3][4] ~^ image[5][10] + kernel[4][0] ~^ image[6][6] + kernel[4][1] ~^ image[6][7] + kernel[4][2] ~^ image[6][8] + kernel[4][3] ~^ image[6][9] + kernel[4][4] ~^ image[6][10];
assign xor_sum[2][7] = kernel[0][0] ~^ image[2][7] + kernel[0][1] ~^ image[2][8] + kernel[0][2] ~^ image[2][9] + kernel[0][3] ~^ image[2][10] + kernel[0][4] ~^ image[2][11] + kernel[1][0] ~^ image[3][7] + kernel[1][1] ~^ image[3][8] + kernel[1][2] ~^ image[3][9] + kernel[1][3] ~^ image[3][10] + kernel[1][4] ~^ image[3][11] + kernel[2][0] ~^ image[4][7] + kernel[2][1] ~^ image[4][8] + kernel[2][2] ~^ image[4][9] + kernel[2][3] ~^ image[4][10] + kernel[2][4] ~^ image[4][11] + kernel[3][0] ~^ image[5][7] + kernel[3][1] ~^ image[5][8] + kernel[3][2] ~^ image[5][9] + kernel[3][3] ~^ image[5][10] + kernel[3][4] ~^ image[5][11] + kernel[4][0] ~^ image[6][7] + kernel[4][1] ~^ image[6][8] + kernel[4][2] ~^ image[6][9] + kernel[4][3] ~^ image[6][10] + kernel[4][4] ~^ image[6][11];
assign xor_sum[3][0] = kernel[0][0] ~^ image[3][0] + kernel[0][1] ~^ image[3][1] + kernel[0][2] ~^ image[3][2] + kernel[0][3] ~^ image[3][3] + kernel[0][4] ~^ image[3][4] + kernel[1][0] ~^ image[4][0] + kernel[1][1] ~^ image[4][1] + kernel[1][2] ~^ image[4][2] + kernel[1][3] ~^ image[4][3] + kernel[1][4] ~^ image[4][4] + kernel[2][0] ~^ image[5][0] + kernel[2][1] ~^ image[5][1] + kernel[2][2] ~^ image[5][2] + kernel[2][3] ~^ image[5][3] + kernel[2][4] ~^ image[5][4] + kernel[3][0] ~^ image[6][0] + kernel[3][1] ~^ image[6][1] + kernel[3][2] ~^ image[6][2] + kernel[3][3] ~^ image[6][3] + kernel[3][4] ~^ image[6][4] + kernel[4][0] ~^ image[7][0] + kernel[4][1] ~^ image[7][1] + kernel[4][2] ~^ image[7][2] + kernel[4][3] ~^ image[7][3] + kernel[4][4] ~^ image[7][4];
assign xor_sum[3][1] = kernel[0][0] ~^ image[3][1] + kernel[0][1] ~^ image[3][2] + kernel[0][2] ~^ image[3][3] + kernel[0][3] ~^ image[3][4] + kernel[0][4] ~^ image[3][5] + kernel[1][0] ~^ image[4][1] + kernel[1][1] ~^ image[4][2] + kernel[1][2] ~^ image[4][3] + kernel[1][3] ~^ image[4][4] + kernel[1][4] ~^ image[4][5] + kernel[2][0] ~^ image[5][1] + kernel[2][1] ~^ image[5][2] + kernel[2][2] ~^ image[5][3] + kernel[2][3] ~^ image[5][4] + kernel[2][4] ~^ image[5][5] + kernel[3][0] ~^ image[6][1] + kernel[3][1] ~^ image[6][2] + kernel[3][2] ~^ image[6][3] + kernel[3][3] ~^ image[6][4] + kernel[3][4] ~^ image[6][5] + kernel[4][0] ~^ image[7][1] + kernel[4][1] ~^ image[7][2] + kernel[4][2] ~^ image[7][3] + kernel[4][3] ~^ image[7][4] + kernel[4][4] ~^ image[7][5];
assign xor_sum[3][2] = kernel[0][0] ~^ image[3][2] + kernel[0][1] ~^ image[3][3] + kernel[0][2] ~^ image[3][4] + kernel[0][3] ~^ image[3][5] + kernel[0][4] ~^ image[3][6] + kernel[1][0] ~^ image[4][2] + kernel[1][1] ~^ image[4][3] + kernel[1][2] ~^ image[4][4] + kernel[1][3] ~^ image[4][5] + kernel[1][4] ~^ image[4][6] + kernel[2][0] ~^ image[5][2] + kernel[2][1] ~^ image[5][3] + kernel[2][2] ~^ image[5][4] + kernel[2][3] ~^ image[5][5] + kernel[2][4] ~^ image[5][6] + kernel[3][0] ~^ image[6][2] + kernel[3][1] ~^ image[6][3] + kernel[3][2] ~^ image[6][4] + kernel[3][3] ~^ image[6][5] + kernel[3][4] ~^ image[6][6] + kernel[4][0] ~^ image[7][2] + kernel[4][1] ~^ image[7][3] + kernel[4][2] ~^ image[7][4] + kernel[4][3] ~^ image[7][5] + kernel[4][4] ~^ image[7][6];
assign xor_sum[3][3] = kernel[0][0] ~^ image[3][3] + kernel[0][1] ~^ image[3][4] + kernel[0][2] ~^ image[3][5] + kernel[0][3] ~^ image[3][6] + kernel[0][4] ~^ image[3][7] + kernel[1][0] ~^ image[4][3] + kernel[1][1] ~^ image[4][4] + kernel[1][2] ~^ image[4][5] + kernel[1][3] ~^ image[4][6] + kernel[1][4] ~^ image[4][7] + kernel[2][0] ~^ image[5][3] + kernel[2][1] ~^ image[5][4] + kernel[2][2] ~^ image[5][5] + kernel[2][3] ~^ image[5][6] + kernel[2][4] ~^ image[5][7] + kernel[3][0] ~^ image[6][3] + kernel[3][1] ~^ image[6][4] + kernel[3][2] ~^ image[6][5] + kernel[3][3] ~^ image[6][6] + kernel[3][4] ~^ image[6][7] + kernel[4][0] ~^ image[7][3] + kernel[4][1] ~^ image[7][4] + kernel[4][2] ~^ image[7][5] + kernel[4][3] ~^ image[7][6] + kernel[4][4] ~^ image[7][7];
assign xor_sum[3][4] = kernel[0][0] ~^ image[3][4] + kernel[0][1] ~^ image[3][5] + kernel[0][2] ~^ image[3][6] + kernel[0][3] ~^ image[3][7] + kernel[0][4] ~^ image[3][8] + kernel[1][0] ~^ image[4][4] + kernel[1][1] ~^ image[4][5] + kernel[1][2] ~^ image[4][6] + kernel[1][3] ~^ image[4][7] + kernel[1][4] ~^ image[4][8] + kernel[2][0] ~^ image[5][4] + kernel[2][1] ~^ image[5][5] + kernel[2][2] ~^ image[5][6] + kernel[2][3] ~^ image[5][7] + kernel[2][4] ~^ image[5][8] + kernel[3][0] ~^ image[6][4] + kernel[3][1] ~^ image[6][5] + kernel[3][2] ~^ image[6][6] + kernel[3][3] ~^ image[6][7] + kernel[3][4] ~^ image[6][8] + kernel[4][0] ~^ image[7][4] + kernel[4][1] ~^ image[7][5] + kernel[4][2] ~^ image[7][6] + kernel[4][3] ~^ image[7][7] + kernel[4][4] ~^ image[7][8];
assign xor_sum[3][5] = kernel[0][0] ~^ image[3][5] + kernel[0][1] ~^ image[3][6] + kernel[0][2] ~^ image[3][7] + kernel[0][3] ~^ image[3][8] + kernel[0][4] ~^ image[3][9] + kernel[1][0] ~^ image[4][5] + kernel[1][1] ~^ image[4][6] + kernel[1][2] ~^ image[4][7] + kernel[1][3] ~^ image[4][8] + kernel[1][4] ~^ image[4][9] + kernel[2][0] ~^ image[5][5] + kernel[2][1] ~^ image[5][6] + kernel[2][2] ~^ image[5][7] + kernel[2][3] ~^ image[5][8] + kernel[2][4] ~^ image[5][9] + kernel[3][0] ~^ image[6][5] + kernel[3][1] ~^ image[6][6] + kernel[3][2] ~^ image[6][7] + kernel[3][3] ~^ image[6][8] + kernel[3][4] ~^ image[6][9] + kernel[4][0] ~^ image[7][5] + kernel[4][1] ~^ image[7][6] + kernel[4][2] ~^ image[7][7] + kernel[4][3] ~^ image[7][8] + kernel[4][4] ~^ image[7][9];
assign xor_sum[3][6] = kernel[0][0] ~^ image[3][6] + kernel[0][1] ~^ image[3][7] + kernel[0][2] ~^ image[3][8] + kernel[0][3] ~^ image[3][9] + kernel[0][4] ~^ image[3][10] + kernel[1][0] ~^ image[4][6] + kernel[1][1] ~^ image[4][7] + kernel[1][2] ~^ image[4][8] + kernel[1][3] ~^ image[4][9] + kernel[1][4] ~^ image[4][10] + kernel[2][0] ~^ image[5][6] + kernel[2][1] ~^ image[5][7] + kernel[2][2] ~^ image[5][8] + kernel[2][3] ~^ image[5][9] + kernel[2][4] ~^ image[5][10] + kernel[3][0] ~^ image[6][6] + kernel[3][1] ~^ image[6][7] + kernel[3][2] ~^ image[6][8] + kernel[3][3] ~^ image[6][9] + kernel[3][4] ~^ image[6][10] + kernel[4][0] ~^ image[7][6] + kernel[4][1] ~^ image[7][7] + kernel[4][2] ~^ image[7][8] + kernel[4][3] ~^ image[7][9] + kernel[4][4] ~^ image[7][10];
assign xor_sum[3][7] = kernel[0][0] ~^ image[3][7] + kernel[0][1] ~^ image[3][8] + kernel[0][2] ~^ image[3][9] + kernel[0][3] ~^ image[3][10] + kernel[0][4] ~^ image[3][11] + kernel[1][0] ~^ image[4][7] + kernel[1][1] ~^ image[4][8] + kernel[1][2] ~^ image[4][9] + kernel[1][3] ~^ image[4][10] + kernel[1][4] ~^ image[4][11] + kernel[2][0] ~^ image[5][7] + kernel[2][1] ~^ image[5][8] + kernel[2][2] ~^ image[5][9] + kernel[2][3] ~^ image[5][10] + kernel[2][4] ~^ image[5][11] + kernel[3][0] ~^ image[6][7] + kernel[3][1] ~^ image[6][8] + kernel[3][2] ~^ image[6][9] + kernel[3][3] ~^ image[6][10] + kernel[3][4] ~^ image[6][11] + kernel[4][0] ~^ image[7][7] + kernel[4][1] ~^ image[7][8] + kernel[4][2] ~^ image[7][9] + kernel[4][3] ~^ image[7][10] + kernel[4][4] ~^ image[7][11];
assign xor_sum[4][0] = kernel[0][0] ~^ image[4][0] + kernel[0][1] ~^ image[4][1] + kernel[0][2] ~^ image[4][2] + kernel[0][3] ~^ image[4][3] + kernel[0][4] ~^ image[4][4] + kernel[1][0] ~^ image[5][0] + kernel[1][1] ~^ image[5][1] + kernel[1][2] ~^ image[5][2] + kernel[1][3] ~^ image[5][3] + kernel[1][4] ~^ image[5][4] + kernel[2][0] ~^ image[6][0] + kernel[2][1] ~^ image[6][1] + kernel[2][2] ~^ image[6][2] + kernel[2][3] ~^ image[6][3] + kernel[2][4] ~^ image[6][4] + kernel[3][0] ~^ image[7][0] + kernel[3][1] ~^ image[7][1] + kernel[3][2] ~^ image[7][2] + kernel[3][3] ~^ image[7][3] + kernel[3][4] ~^ image[7][4] + kernel[4][0] ~^ image[8][0] + kernel[4][1] ~^ image[8][1] + kernel[4][2] ~^ image[8][2] + kernel[4][3] ~^ image[8][3] + kernel[4][4] ~^ image[8][4];
assign xor_sum[4][1] = kernel[0][0] ~^ image[4][1] + kernel[0][1] ~^ image[4][2] + kernel[0][2] ~^ image[4][3] + kernel[0][3] ~^ image[4][4] + kernel[0][4] ~^ image[4][5] + kernel[1][0] ~^ image[5][1] + kernel[1][1] ~^ image[5][2] + kernel[1][2] ~^ image[5][3] + kernel[1][3] ~^ image[5][4] + kernel[1][4] ~^ image[5][5] + kernel[2][0] ~^ image[6][1] + kernel[2][1] ~^ image[6][2] + kernel[2][2] ~^ image[6][3] + kernel[2][3] ~^ image[6][4] + kernel[2][4] ~^ image[6][5] + kernel[3][0] ~^ image[7][1] + kernel[3][1] ~^ image[7][2] + kernel[3][2] ~^ image[7][3] + kernel[3][3] ~^ image[7][4] + kernel[3][4] ~^ image[7][5] + kernel[4][0] ~^ image[8][1] + kernel[4][1] ~^ image[8][2] + kernel[4][2] ~^ image[8][3] + kernel[4][3] ~^ image[8][4] + kernel[4][4] ~^ image[8][5];
assign xor_sum[4][2] = kernel[0][0] ~^ image[4][2] + kernel[0][1] ~^ image[4][3] + kernel[0][2] ~^ image[4][4] + kernel[0][3] ~^ image[4][5] + kernel[0][4] ~^ image[4][6] + kernel[1][0] ~^ image[5][2] + kernel[1][1] ~^ image[5][3] + kernel[1][2] ~^ image[5][4] + kernel[1][3] ~^ image[5][5] + kernel[1][4] ~^ image[5][6] + kernel[2][0] ~^ image[6][2] + kernel[2][1] ~^ image[6][3] + kernel[2][2] ~^ image[6][4] + kernel[2][3] ~^ image[6][5] + kernel[2][4] ~^ image[6][6] + kernel[3][0] ~^ image[7][2] + kernel[3][1] ~^ image[7][3] + kernel[3][2] ~^ image[7][4] + kernel[3][3] ~^ image[7][5] + kernel[3][4] ~^ image[7][6] + kernel[4][0] ~^ image[8][2] + kernel[4][1] ~^ image[8][3] + kernel[4][2] ~^ image[8][4] + kernel[4][3] ~^ image[8][5] + kernel[4][4] ~^ image[8][6];
assign xor_sum[4][3] = kernel[0][0] ~^ image[4][3] + kernel[0][1] ~^ image[4][4] + kernel[0][2] ~^ image[4][5] + kernel[0][3] ~^ image[4][6] + kernel[0][4] ~^ image[4][7] + kernel[1][0] ~^ image[5][3] + kernel[1][1] ~^ image[5][4] + kernel[1][2] ~^ image[5][5] + kernel[1][3] ~^ image[5][6] + kernel[1][4] ~^ image[5][7] + kernel[2][0] ~^ image[6][3] + kernel[2][1] ~^ image[6][4] + kernel[2][2] ~^ image[6][5] + kernel[2][3] ~^ image[6][6] + kernel[2][4] ~^ image[6][7] + kernel[3][0] ~^ image[7][3] + kernel[3][1] ~^ image[7][4] + kernel[3][2] ~^ image[7][5] + kernel[3][3] ~^ image[7][6] + kernel[3][4] ~^ image[7][7] + kernel[4][0] ~^ image[8][3] + kernel[4][1] ~^ image[8][4] + kernel[4][2] ~^ image[8][5] + kernel[4][3] ~^ image[8][6] + kernel[4][4] ~^ image[8][7];
assign xor_sum[4][4] = kernel[0][0] ~^ image[4][4] + kernel[0][1] ~^ image[4][5] + kernel[0][2] ~^ image[4][6] + kernel[0][3] ~^ image[4][7] + kernel[0][4] ~^ image[4][8] + kernel[1][0] ~^ image[5][4] + kernel[1][1] ~^ image[5][5] + kernel[1][2] ~^ image[5][6] + kernel[1][3] ~^ image[5][7] + kernel[1][4] ~^ image[5][8] + kernel[2][0] ~^ image[6][4] + kernel[2][1] ~^ image[6][5] + kernel[2][2] ~^ image[6][6] + kernel[2][3] ~^ image[6][7] + kernel[2][4] ~^ image[6][8] + kernel[3][0] ~^ image[7][4] + kernel[3][1] ~^ image[7][5] + kernel[3][2] ~^ image[7][6] + kernel[3][3] ~^ image[7][7] + kernel[3][4] ~^ image[7][8] + kernel[4][0] ~^ image[8][4] + kernel[4][1] ~^ image[8][5] + kernel[4][2] ~^ image[8][6] + kernel[4][3] ~^ image[8][7] + kernel[4][4] ~^ image[8][8];
assign xor_sum[4][5] = kernel[0][0] ~^ image[4][5] + kernel[0][1] ~^ image[4][6] + kernel[0][2] ~^ image[4][7] + kernel[0][3] ~^ image[4][8] + kernel[0][4] ~^ image[4][9] + kernel[1][0] ~^ image[5][5] + kernel[1][1] ~^ image[5][6] + kernel[1][2] ~^ image[5][7] + kernel[1][3] ~^ image[5][8] + kernel[1][4] ~^ image[5][9] + kernel[2][0] ~^ image[6][5] + kernel[2][1] ~^ image[6][6] + kernel[2][2] ~^ image[6][7] + kernel[2][3] ~^ image[6][8] + kernel[2][4] ~^ image[6][9] + kernel[3][0] ~^ image[7][5] + kernel[3][1] ~^ image[7][6] + kernel[3][2] ~^ image[7][7] + kernel[3][3] ~^ image[7][8] + kernel[3][4] ~^ image[7][9] + kernel[4][0] ~^ image[8][5] + kernel[4][1] ~^ image[8][6] + kernel[4][2] ~^ image[8][7] + kernel[4][3] ~^ image[8][8] + kernel[4][4] ~^ image[8][9];
assign xor_sum[4][6] = kernel[0][0] ~^ image[4][6] + kernel[0][1] ~^ image[4][7] + kernel[0][2] ~^ image[4][8] + kernel[0][3] ~^ image[4][9] + kernel[0][4] ~^ image[4][10] + kernel[1][0] ~^ image[5][6] + kernel[1][1] ~^ image[5][7] + kernel[1][2] ~^ image[5][8] + kernel[1][3] ~^ image[5][9] + kernel[1][4] ~^ image[5][10] + kernel[2][0] ~^ image[6][6] + kernel[2][1] ~^ image[6][7] + kernel[2][2] ~^ image[6][8] + kernel[2][3] ~^ image[6][9] + kernel[2][4] ~^ image[6][10] + kernel[3][0] ~^ image[7][6] + kernel[3][1] ~^ image[7][7] + kernel[3][2] ~^ image[7][8] + kernel[3][3] ~^ image[7][9] + kernel[3][4] ~^ image[7][10] + kernel[4][0] ~^ image[8][6] + kernel[4][1] ~^ image[8][7] + kernel[4][2] ~^ image[8][8] + kernel[4][3] ~^ image[8][9] + kernel[4][4] ~^ image[8][10];
assign xor_sum[4][7] = kernel[0][0] ~^ image[4][7] + kernel[0][1] ~^ image[4][8] + kernel[0][2] ~^ image[4][9] + kernel[0][3] ~^ image[4][10] + kernel[0][4] ~^ image[4][11] + kernel[1][0] ~^ image[5][7] + kernel[1][1] ~^ image[5][8] + kernel[1][2] ~^ image[5][9] + kernel[1][3] ~^ image[5][10] + kernel[1][4] ~^ image[5][11] + kernel[2][0] ~^ image[6][7] + kernel[2][1] ~^ image[6][8] + kernel[2][2] ~^ image[6][9] + kernel[2][3] ~^ image[6][10] + kernel[2][4] ~^ image[6][11] + kernel[3][0] ~^ image[7][7] + kernel[3][1] ~^ image[7][8] + kernel[3][2] ~^ image[7][9] + kernel[3][3] ~^ image[7][10] + kernel[3][4] ~^ image[7][11] + kernel[4][0] ~^ image[8][7] + kernel[4][1] ~^ image[8][8] + kernel[4][2] ~^ image[8][9] + kernel[4][3] ~^ image[8][10] + kernel[4][4] ~^ image[8][11];
assign xor_sum[5][0] = kernel[0][0] ~^ image[5][0] + kernel[0][1] ~^ image[5][1] + kernel[0][2] ~^ image[5][2] + kernel[0][3] ~^ image[5][3] + kernel[0][4] ~^ image[5][4] + kernel[1][0] ~^ image[6][0] + kernel[1][1] ~^ image[6][1] + kernel[1][2] ~^ image[6][2] + kernel[1][3] ~^ image[6][3] + kernel[1][4] ~^ image[6][4] + kernel[2][0] ~^ image[7][0] + kernel[2][1] ~^ image[7][1] + kernel[2][2] ~^ image[7][2] + kernel[2][3] ~^ image[7][3] + kernel[2][4] ~^ image[7][4] + kernel[3][0] ~^ image[8][0] + kernel[3][1] ~^ image[8][1] + kernel[3][2] ~^ image[8][2] + kernel[3][3] ~^ image[8][3] + kernel[3][4] ~^ image[8][4] + kernel[4][0] ~^ image[9][0] + kernel[4][1] ~^ image[9][1] + kernel[4][2] ~^ image[9][2] + kernel[4][3] ~^ image[9][3] + kernel[4][4] ~^ image[9][4];
assign xor_sum[5][1] = kernel[0][0] ~^ image[5][1] + kernel[0][1] ~^ image[5][2] + kernel[0][2] ~^ image[5][3] + kernel[0][3] ~^ image[5][4] + kernel[0][4] ~^ image[5][5] + kernel[1][0] ~^ image[6][1] + kernel[1][1] ~^ image[6][2] + kernel[1][2] ~^ image[6][3] + kernel[1][3] ~^ image[6][4] + kernel[1][4] ~^ image[6][5] + kernel[2][0] ~^ image[7][1] + kernel[2][1] ~^ image[7][2] + kernel[2][2] ~^ image[7][3] + kernel[2][3] ~^ image[7][4] + kernel[2][4] ~^ image[7][5] + kernel[3][0] ~^ image[8][1] + kernel[3][1] ~^ image[8][2] + kernel[3][2] ~^ image[8][3] + kernel[3][3] ~^ image[8][4] + kernel[3][4] ~^ image[8][5] + kernel[4][0] ~^ image[9][1] + kernel[4][1] ~^ image[9][2] + kernel[4][2] ~^ image[9][3] + kernel[4][3] ~^ image[9][4] + kernel[4][4] ~^ image[9][5];
assign xor_sum[5][2] = kernel[0][0] ~^ image[5][2] + kernel[0][1] ~^ image[5][3] + kernel[0][2] ~^ image[5][4] + kernel[0][3] ~^ image[5][5] + kernel[0][4] ~^ image[5][6] + kernel[1][0] ~^ image[6][2] + kernel[1][1] ~^ image[6][3] + kernel[1][2] ~^ image[6][4] + kernel[1][3] ~^ image[6][5] + kernel[1][4] ~^ image[6][6] + kernel[2][0] ~^ image[7][2] + kernel[2][1] ~^ image[7][3] + kernel[2][2] ~^ image[7][4] + kernel[2][3] ~^ image[7][5] + kernel[2][4] ~^ image[7][6] + kernel[3][0] ~^ image[8][2] + kernel[3][1] ~^ image[8][3] + kernel[3][2] ~^ image[8][4] + kernel[3][3] ~^ image[8][5] + kernel[3][4] ~^ image[8][6] + kernel[4][0] ~^ image[9][2] + kernel[4][1] ~^ image[9][3] + kernel[4][2] ~^ image[9][4] + kernel[4][3] ~^ image[9][5] + kernel[4][4] ~^ image[9][6];
assign xor_sum[5][3] = kernel[0][0] ~^ image[5][3] + kernel[0][1] ~^ image[5][4] + kernel[0][2] ~^ image[5][5] + kernel[0][3] ~^ image[5][6] + kernel[0][4] ~^ image[5][7] + kernel[1][0] ~^ image[6][3] + kernel[1][1] ~^ image[6][4] + kernel[1][2] ~^ image[6][5] + kernel[1][3] ~^ image[6][6] + kernel[1][4] ~^ image[6][7] + kernel[2][0] ~^ image[7][3] + kernel[2][1] ~^ image[7][4] + kernel[2][2] ~^ image[7][5] + kernel[2][3] ~^ image[7][6] + kernel[2][4] ~^ image[7][7] + kernel[3][0] ~^ image[8][3] + kernel[3][1] ~^ image[8][4] + kernel[3][2] ~^ image[8][5] + kernel[3][3] ~^ image[8][6] + kernel[3][4] ~^ image[8][7] + kernel[4][0] ~^ image[9][3] + kernel[4][1] ~^ image[9][4] + kernel[4][2] ~^ image[9][5] + kernel[4][3] ~^ image[9][6] + kernel[4][4] ~^ image[9][7];
assign xor_sum[5][4] = kernel[0][0] ~^ image[5][4] + kernel[0][1] ~^ image[5][5] + kernel[0][2] ~^ image[5][6] + kernel[0][3] ~^ image[5][7] + kernel[0][4] ~^ image[5][8] + kernel[1][0] ~^ image[6][4] + kernel[1][1] ~^ image[6][5] + kernel[1][2] ~^ image[6][6] + kernel[1][3] ~^ image[6][7] + kernel[1][4] ~^ image[6][8] + kernel[2][0] ~^ image[7][4] + kernel[2][1] ~^ image[7][5] + kernel[2][2] ~^ image[7][6] + kernel[2][3] ~^ image[7][7] + kernel[2][4] ~^ image[7][8] + kernel[3][0] ~^ image[8][4] + kernel[3][1] ~^ image[8][5] + kernel[3][2] ~^ image[8][6] + kernel[3][3] ~^ image[8][7] + kernel[3][4] ~^ image[8][8] + kernel[4][0] ~^ image[9][4] + kernel[4][1] ~^ image[9][5] + kernel[4][2] ~^ image[9][6] + kernel[4][3] ~^ image[9][7] + kernel[4][4] ~^ image[9][8];
assign xor_sum[5][5] = kernel[0][0] ~^ image[5][5] + kernel[0][1] ~^ image[5][6] + kernel[0][2] ~^ image[5][7] + kernel[0][3] ~^ image[5][8] + kernel[0][4] ~^ image[5][9] + kernel[1][0] ~^ image[6][5] + kernel[1][1] ~^ image[6][6] + kernel[1][2] ~^ image[6][7] + kernel[1][3] ~^ image[6][8] + kernel[1][4] ~^ image[6][9] + kernel[2][0] ~^ image[7][5] + kernel[2][1] ~^ image[7][6] + kernel[2][2] ~^ image[7][7] + kernel[2][3] ~^ image[7][8] + kernel[2][4] ~^ image[7][9] + kernel[3][0] ~^ image[8][5] + kernel[3][1] ~^ image[8][6] + kernel[3][2] ~^ image[8][7] + kernel[3][3] ~^ image[8][8] + kernel[3][4] ~^ image[8][9] + kernel[4][0] ~^ image[9][5] + kernel[4][1] ~^ image[9][6] + kernel[4][2] ~^ image[9][7] + kernel[4][3] ~^ image[9][8] + kernel[4][4] ~^ image[9][9];
assign xor_sum[5][6] = kernel[0][0] ~^ image[5][6] + kernel[0][1] ~^ image[5][7] + kernel[0][2] ~^ image[5][8] + kernel[0][3] ~^ image[5][9] + kernel[0][4] ~^ image[5][10] + kernel[1][0] ~^ image[6][6] + kernel[1][1] ~^ image[6][7] + kernel[1][2] ~^ image[6][8] + kernel[1][3] ~^ image[6][9] + kernel[1][4] ~^ image[6][10] + kernel[2][0] ~^ image[7][6] + kernel[2][1] ~^ image[7][7] + kernel[2][2] ~^ image[7][8] + kernel[2][3] ~^ image[7][9] + kernel[2][4] ~^ image[7][10] + kernel[3][0] ~^ image[8][6] + kernel[3][1] ~^ image[8][7] + kernel[3][2] ~^ image[8][8] + kernel[3][3] ~^ image[8][9] + kernel[3][4] ~^ image[8][10] + kernel[4][0] ~^ image[9][6] + kernel[4][1] ~^ image[9][7] + kernel[4][2] ~^ image[9][8] + kernel[4][3] ~^ image[9][9] + kernel[4][4] ~^ image[9][10];
assign xor_sum[5][7] = kernel[0][0] ~^ image[5][7] + kernel[0][1] ~^ image[5][8] + kernel[0][2] ~^ image[5][9] + kernel[0][3] ~^ image[5][10] + kernel[0][4] ~^ image[5][11] + kernel[1][0] ~^ image[6][7] + kernel[1][1] ~^ image[6][8] + kernel[1][2] ~^ image[6][9] + kernel[1][3] ~^ image[6][10] + kernel[1][4] ~^ image[6][11] + kernel[2][0] ~^ image[7][7] + kernel[2][1] ~^ image[7][8] + kernel[2][2] ~^ image[7][9] + kernel[2][3] ~^ image[7][10] + kernel[2][4] ~^ image[7][11] + kernel[3][0] ~^ image[8][7] + kernel[3][1] ~^ image[8][8] + kernel[3][2] ~^ image[8][9] + kernel[3][3] ~^ image[8][10] + kernel[3][4] ~^ image[8][11] + kernel[4][0] ~^ image[9][7] + kernel[4][1] ~^ image[9][8] + kernel[4][2] ~^ image[9][9] + kernel[4][3] ~^ image[9][10] + kernel[4][4] ~^ image[9][11];
assign xor_sum[6][0] = kernel[0][0] ~^ image[6][0] + kernel[0][1] ~^ image[6][1] + kernel[0][2] ~^ image[6][2] + kernel[0][3] ~^ image[6][3] + kernel[0][4] ~^ image[6][4] + kernel[1][0] ~^ image[7][0] + kernel[1][1] ~^ image[7][1] + kernel[1][2] ~^ image[7][2] + kernel[1][3] ~^ image[7][3] + kernel[1][4] ~^ image[7][4] + kernel[2][0] ~^ image[8][0] + kernel[2][1] ~^ image[8][1] + kernel[2][2] ~^ image[8][2] + kernel[2][3] ~^ image[8][3] + kernel[2][4] ~^ image[8][4] + kernel[3][0] ~^ image[9][0] + kernel[3][1] ~^ image[9][1] + kernel[3][2] ~^ image[9][2] + kernel[3][3] ~^ image[9][3] + kernel[3][4] ~^ image[9][4] + kernel[4][0] ~^ image[10][0] + kernel[4][1] ~^ image[10][1] + kernel[4][2] ~^ image[10][2] + kernel[4][3] ~^ image[10][3] + kernel[4][4] ~^ image[10][4];
assign xor_sum[6][1] = kernel[0][0] ~^ image[6][1] + kernel[0][1] ~^ image[6][2] + kernel[0][2] ~^ image[6][3] + kernel[0][3] ~^ image[6][4] + kernel[0][4] ~^ image[6][5] + kernel[1][0] ~^ image[7][1] + kernel[1][1] ~^ image[7][2] + kernel[1][2] ~^ image[7][3] + kernel[1][3] ~^ image[7][4] + kernel[1][4] ~^ image[7][5] + kernel[2][0] ~^ image[8][1] + kernel[2][1] ~^ image[8][2] + kernel[2][2] ~^ image[8][3] + kernel[2][3] ~^ image[8][4] + kernel[2][4] ~^ image[8][5] + kernel[3][0] ~^ image[9][1] + kernel[3][1] ~^ image[9][2] + kernel[3][2] ~^ image[9][3] + kernel[3][3] ~^ image[9][4] + kernel[3][4] ~^ image[9][5] + kernel[4][0] ~^ image[10][1] + kernel[4][1] ~^ image[10][2] + kernel[4][2] ~^ image[10][3] + kernel[4][3] ~^ image[10][4] + kernel[4][4] ~^ image[10][5];
assign xor_sum[6][2] = kernel[0][0] ~^ image[6][2] + kernel[0][1] ~^ image[6][3] + kernel[0][2] ~^ image[6][4] + kernel[0][3] ~^ image[6][5] + kernel[0][4] ~^ image[6][6] + kernel[1][0] ~^ image[7][2] + kernel[1][1] ~^ image[7][3] + kernel[1][2] ~^ image[7][4] + kernel[1][3] ~^ image[7][5] + kernel[1][4] ~^ image[7][6] + kernel[2][0] ~^ image[8][2] + kernel[2][1] ~^ image[8][3] + kernel[2][2] ~^ image[8][4] + kernel[2][3] ~^ image[8][5] + kernel[2][4] ~^ image[8][6] + kernel[3][0] ~^ image[9][2] + kernel[3][1] ~^ image[9][3] + kernel[3][2] ~^ image[9][4] + kernel[3][3] ~^ image[9][5] + kernel[3][4] ~^ image[9][6] + kernel[4][0] ~^ image[10][2] + kernel[4][1] ~^ image[10][3] + kernel[4][2] ~^ image[10][4] + kernel[4][3] ~^ image[10][5] + kernel[4][4] ~^ image[10][6];
assign xor_sum[6][3] = kernel[0][0] ~^ image[6][3] + kernel[0][1] ~^ image[6][4] + kernel[0][2] ~^ image[6][5] + kernel[0][3] ~^ image[6][6] + kernel[0][4] ~^ image[6][7] + kernel[1][0] ~^ image[7][3] + kernel[1][1] ~^ image[7][4] + kernel[1][2] ~^ image[7][5] + kernel[1][3] ~^ image[7][6] + kernel[1][4] ~^ image[7][7] + kernel[2][0] ~^ image[8][3] + kernel[2][1] ~^ image[8][4] + kernel[2][2] ~^ image[8][5] + kernel[2][3] ~^ image[8][6] + kernel[2][4] ~^ image[8][7] + kernel[3][0] ~^ image[9][3] + kernel[3][1] ~^ image[9][4] + kernel[3][2] ~^ image[9][5] + kernel[3][3] ~^ image[9][6] + kernel[3][4] ~^ image[9][7] + kernel[4][0] ~^ image[10][3] + kernel[4][1] ~^ image[10][4] + kernel[4][2] ~^ image[10][5] + kernel[4][3] ~^ image[10][6] + kernel[4][4] ~^ image[10][7];
assign xor_sum[6][4] = kernel[0][0] ~^ image[6][4] + kernel[0][1] ~^ image[6][5] + kernel[0][2] ~^ image[6][6] + kernel[0][3] ~^ image[6][7] + kernel[0][4] ~^ image[6][8] + kernel[1][0] ~^ image[7][4] + kernel[1][1] ~^ image[7][5] + kernel[1][2] ~^ image[7][6] + kernel[1][3] ~^ image[7][7] + kernel[1][4] ~^ image[7][8] + kernel[2][0] ~^ image[8][4] + kernel[2][1] ~^ image[8][5] + kernel[2][2] ~^ image[8][6] + kernel[2][3] ~^ image[8][7] + kernel[2][4] ~^ image[8][8] + kernel[3][0] ~^ image[9][4] + kernel[3][1] ~^ image[9][5] + kernel[3][2] ~^ image[9][6] + kernel[3][3] ~^ image[9][7] + kernel[3][4] ~^ image[9][8] + kernel[4][0] ~^ image[10][4] + kernel[4][1] ~^ image[10][5] + kernel[4][2] ~^ image[10][6] + kernel[4][3] ~^ image[10][7] + kernel[4][4] ~^ image[10][8];
assign xor_sum[6][5] = kernel[0][0] ~^ image[6][5] + kernel[0][1] ~^ image[6][6] + kernel[0][2] ~^ image[6][7] + kernel[0][3] ~^ image[6][8] + kernel[0][4] ~^ image[6][9] + kernel[1][0] ~^ image[7][5] + kernel[1][1] ~^ image[7][6] + kernel[1][2] ~^ image[7][7] + kernel[1][3] ~^ image[7][8] + kernel[1][4] ~^ image[7][9] + kernel[2][0] ~^ image[8][5] + kernel[2][1] ~^ image[8][6] + kernel[2][2] ~^ image[8][7] + kernel[2][3] ~^ image[8][8] + kernel[2][4] ~^ image[8][9] + kernel[3][0] ~^ image[9][5] + kernel[3][1] ~^ image[9][6] + kernel[3][2] ~^ image[9][7] + kernel[3][3] ~^ image[9][8] + kernel[3][4] ~^ image[9][9] + kernel[4][0] ~^ image[10][5] + kernel[4][1] ~^ image[10][6] + kernel[4][2] ~^ image[10][7] + kernel[4][3] ~^ image[10][8] + kernel[4][4] ~^ image[10][9];
assign xor_sum[6][6] = kernel[0][0] ~^ image[6][6] + kernel[0][1] ~^ image[6][7] + kernel[0][2] ~^ image[6][8] + kernel[0][3] ~^ image[6][9] + kernel[0][4] ~^ image[6][10] + kernel[1][0] ~^ image[7][6] + kernel[1][1] ~^ image[7][7] + kernel[1][2] ~^ image[7][8] + kernel[1][3] ~^ image[7][9] + kernel[1][4] ~^ image[7][10] + kernel[2][0] ~^ image[8][6] + kernel[2][1] ~^ image[8][7] + kernel[2][2] ~^ image[8][8] + kernel[2][3] ~^ image[8][9] + kernel[2][4] ~^ image[8][10] + kernel[3][0] ~^ image[9][6] + kernel[3][1] ~^ image[9][7] + kernel[3][2] ~^ image[9][8] + kernel[3][3] ~^ image[9][9] + kernel[3][4] ~^ image[9][10] + kernel[4][0] ~^ image[10][6] + kernel[4][1] ~^ image[10][7] + kernel[4][2] ~^ image[10][8] + kernel[4][3] ~^ image[10][9] + kernel[4][4] ~^ image[10][10];
assign xor_sum[6][7] = kernel[0][0] ~^ image[6][7] + kernel[0][1] ~^ image[6][8] + kernel[0][2] ~^ image[6][9] + kernel[0][3] ~^ image[6][10] + kernel[0][4] ~^ image[6][11] + kernel[1][0] ~^ image[7][7] + kernel[1][1] ~^ image[7][8] + kernel[1][2] ~^ image[7][9] + kernel[1][3] ~^ image[7][10] + kernel[1][4] ~^ image[7][11] + kernel[2][0] ~^ image[8][7] + kernel[2][1] ~^ image[8][8] + kernel[2][2] ~^ image[8][9] + kernel[2][3] ~^ image[8][10] + kernel[2][4] ~^ image[8][11] + kernel[3][0] ~^ image[9][7] + kernel[3][1] ~^ image[9][8] + kernel[3][2] ~^ image[9][9] + kernel[3][3] ~^ image[9][10] + kernel[3][4] ~^ image[9][11] + kernel[4][0] ~^ image[10][7] + kernel[4][1] ~^ image[10][8] + kernel[4][2] ~^ image[10][9] + kernel[4][3] ~^ image[10][10] + kernel[4][4] ~^ image[10][11];
assign xor_sum[7][0] = kernel[0][0] ~^ image[7][0] + kernel[0][1] ~^ image[7][1] + kernel[0][2] ~^ image[7][2] + kernel[0][3] ~^ image[7][3] + kernel[0][4] ~^ image[7][4] + kernel[1][0] ~^ image[8][0] + kernel[1][1] ~^ image[8][1] + kernel[1][2] ~^ image[8][2] + kernel[1][3] ~^ image[8][3] + kernel[1][4] ~^ image[8][4] + kernel[2][0] ~^ image[9][0] + kernel[2][1] ~^ image[9][1] + kernel[2][2] ~^ image[9][2] + kernel[2][3] ~^ image[9][3] + kernel[2][4] ~^ image[9][4] + kernel[3][0] ~^ image[10][0] + kernel[3][1] ~^ image[10][1] + kernel[3][2] ~^ image[10][2] + kernel[3][3] ~^ image[10][3] + kernel[3][4] ~^ image[10][4] + kernel[4][0] ~^ image[11][0] + kernel[4][1] ~^ image[11][1] + kernel[4][2] ~^ image[11][2] + kernel[4][3] ~^ image[11][3] + kernel[4][4] ~^ image[11][4];
assign xor_sum[7][1] = kernel[0][0] ~^ image[7][1] + kernel[0][1] ~^ image[7][2] + kernel[0][2] ~^ image[7][3] + kernel[0][3] ~^ image[7][4] + kernel[0][4] ~^ image[7][5] + kernel[1][0] ~^ image[8][1] + kernel[1][1] ~^ image[8][2] + kernel[1][2] ~^ image[8][3] + kernel[1][3] ~^ image[8][4] + kernel[1][4] ~^ image[8][5] + kernel[2][0] ~^ image[9][1] + kernel[2][1] ~^ image[9][2] + kernel[2][2] ~^ image[9][3] + kernel[2][3] ~^ image[9][4] + kernel[2][4] ~^ image[9][5] + kernel[3][0] ~^ image[10][1] + kernel[3][1] ~^ image[10][2] + kernel[3][2] ~^ image[10][3] + kernel[3][3] ~^ image[10][4] + kernel[3][4] ~^ image[10][5] + kernel[4][0] ~^ image[11][1] + kernel[4][1] ~^ image[11][2] + kernel[4][2] ~^ image[11][3] + kernel[4][3] ~^ image[11][4] + kernel[4][4] ~^ image[11][5];
assign xor_sum[7][2] = kernel[0][0] ~^ image[7][2] + kernel[0][1] ~^ image[7][3] + kernel[0][2] ~^ image[7][4] + kernel[0][3] ~^ image[7][5] + kernel[0][4] ~^ image[7][6] + kernel[1][0] ~^ image[8][2] + kernel[1][1] ~^ image[8][3] + kernel[1][2] ~^ image[8][4] + kernel[1][3] ~^ image[8][5] + kernel[1][4] ~^ image[8][6] + kernel[2][0] ~^ image[9][2] + kernel[2][1] ~^ image[9][3] + kernel[2][2] ~^ image[9][4] + kernel[2][3] ~^ image[9][5] + kernel[2][4] ~^ image[9][6] + kernel[3][0] ~^ image[10][2] + kernel[3][1] ~^ image[10][3] + kernel[3][2] ~^ image[10][4] + kernel[3][3] ~^ image[10][5] + kernel[3][4] ~^ image[10][6] + kernel[4][0] ~^ image[11][2] + kernel[4][1] ~^ image[11][3] + kernel[4][2] ~^ image[11][4] + kernel[4][3] ~^ image[11][5] + kernel[4][4] ~^ image[11][6];
assign xor_sum[7][3] = kernel[0][0] ~^ image[7][3] + kernel[0][1] ~^ image[7][4] + kernel[0][2] ~^ image[7][5] + kernel[0][3] ~^ image[7][6] + kernel[0][4] ~^ image[7][7] + kernel[1][0] ~^ image[8][3] + kernel[1][1] ~^ image[8][4] + kernel[1][2] ~^ image[8][5] + kernel[1][3] ~^ image[8][6] + kernel[1][4] ~^ image[8][7] + kernel[2][0] ~^ image[9][3] + kernel[2][1] ~^ image[9][4] + kernel[2][2] ~^ image[9][5] + kernel[2][3] ~^ image[9][6] + kernel[2][4] ~^ image[9][7] + kernel[3][0] ~^ image[10][3] + kernel[3][1] ~^ image[10][4] + kernel[3][2] ~^ image[10][5] + kernel[3][3] ~^ image[10][6] + kernel[3][4] ~^ image[10][7] + kernel[4][0] ~^ image[11][3] + kernel[4][1] ~^ image[11][4] + kernel[4][2] ~^ image[11][5] + kernel[4][3] ~^ image[11][6] + kernel[4][4] ~^ image[11][7];
assign xor_sum[7][4] = kernel[0][0] ~^ image[7][4] + kernel[0][1] ~^ image[7][5] + kernel[0][2] ~^ image[7][6] + kernel[0][3] ~^ image[7][7] + kernel[0][4] ~^ image[7][8] + kernel[1][0] ~^ image[8][4] + kernel[1][1] ~^ image[8][5] + kernel[1][2] ~^ image[8][6] + kernel[1][3] ~^ image[8][7] + kernel[1][4] ~^ image[8][8] + kernel[2][0] ~^ image[9][4] + kernel[2][1] ~^ image[9][5] + kernel[2][2] ~^ image[9][6] + kernel[2][3] ~^ image[9][7] + kernel[2][4] ~^ image[9][8] + kernel[3][0] ~^ image[10][4] + kernel[3][1] ~^ image[10][5] + kernel[3][2] ~^ image[10][6] + kernel[3][3] ~^ image[10][7] + kernel[3][4] ~^ image[10][8] + kernel[4][0] ~^ image[11][4] + kernel[4][1] ~^ image[11][5] + kernel[4][2] ~^ image[11][6] + kernel[4][3] ~^ image[11][7] + kernel[4][4] ~^ image[11][8];
assign xor_sum[7][5] = kernel[0][0] ~^ image[7][5] + kernel[0][1] ~^ image[7][6] + kernel[0][2] ~^ image[7][7] + kernel[0][3] ~^ image[7][8] + kernel[0][4] ~^ image[7][9] + kernel[1][0] ~^ image[8][5] + kernel[1][1] ~^ image[8][6] + kernel[1][2] ~^ image[8][7] + kernel[1][3] ~^ image[8][8] + kernel[1][4] ~^ image[8][9] + kernel[2][0] ~^ image[9][5] + kernel[2][1] ~^ image[9][6] + kernel[2][2] ~^ image[9][7] + kernel[2][3] ~^ image[9][8] + kernel[2][4] ~^ image[9][9] + kernel[3][0] ~^ image[10][5] + kernel[3][1] ~^ image[10][6] + kernel[3][2] ~^ image[10][7] + kernel[3][3] ~^ image[10][8] + kernel[3][4] ~^ image[10][9] + kernel[4][0] ~^ image[11][5] + kernel[4][1] ~^ image[11][6] + kernel[4][2] ~^ image[11][7] + kernel[4][3] ~^ image[11][8] + kernel[4][4] ~^ image[11][9];
assign xor_sum[7][6] = kernel[0][0] ~^ image[7][6] + kernel[0][1] ~^ image[7][7] + kernel[0][2] ~^ image[7][8] + kernel[0][3] ~^ image[7][9] + kernel[0][4] ~^ image[7][10] + kernel[1][0] ~^ image[8][6] + kernel[1][1] ~^ image[8][7] + kernel[1][2] ~^ image[8][8] + kernel[1][3] ~^ image[8][9] + kernel[1][4] ~^ image[8][10] + kernel[2][0] ~^ image[9][6] + kernel[2][1] ~^ image[9][7] + kernel[2][2] ~^ image[9][8] + kernel[2][3] ~^ image[9][9] + kernel[2][4] ~^ image[9][10] + kernel[3][0] ~^ image[10][6] + kernel[3][1] ~^ image[10][7] + kernel[3][2] ~^ image[10][8] + kernel[3][3] ~^ image[10][9] + kernel[3][4] ~^ image[10][10] + kernel[4][0] ~^ image[11][6] + kernel[4][1] ~^ image[11][7] + kernel[4][2] ~^ image[11][8] + kernel[4][3] ~^ image[11][9] + kernel[4][4] ~^ image[11][10];
assign xor_sum[7][7] = kernel[0][0] ~^ image[7][7] + kernel[0][1] ~^ image[7][8] + kernel[0][2] ~^ image[7][9] + kernel[0][3] ~^ image[7][10] + kernel[0][4] ~^ image[7][11] + kernel[1][0] ~^ image[8][7] + kernel[1][1] ~^ image[8][8] + kernel[1][2] ~^ image[8][9] + kernel[1][3] ~^ image[8][10] + kernel[1][4] ~^ image[8][11] + kernel[2][0] ~^ image[9][7] + kernel[2][1] ~^ image[9][8] + kernel[2][2] ~^ image[9][9] + kernel[2][3] ~^ image[9][10] + kernel[2][4] ~^ image[9][11] + kernel[3][0] ~^ image[10][7] + kernel[3][1] ~^ image[10][8] + kernel[3][2] ~^ image[10][9] + kernel[3][3] ~^ image[10][10] + kernel[3][4] ~^ image[10][11] + kernel[4][0] ~^ image[11][7] + kernel[4][1] ~^ image[11][8] + kernel[4][2] ~^ image[11][9] + kernel[4][3] ~^ image[11][10] + kernel[4][4] ~^ image[11][11];


 // output just the sign bit 

assign out_fmap[0][0] = xor_sum[0][0][0];
assign out_fmap[0][1] = xor_sum[0][1][0];
assign out_fmap[0][2] = xor_sum[0][2][0];
assign out_fmap[0][3] = xor_sum[0][3][0];
assign out_fmap[0][4] = xor_sum[0][4][0];
assign out_fmap[0][5] = xor_sum[0][5][0];
assign out_fmap[0][6] = xor_sum[0][6][0];
assign out_fmap[0][7] = xor_sum[0][7][0];
assign out_fmap[0][8] = xor_sum[0][8][0];
assign out_fmap[0][9] = xor_sum[0][9][0];
assign out_fmap[0][10] = xor_sum[0][10][0];
assign out_fmap[0][11] = xor_sum[0][11][0];
assign out_fmap[0][12] = xor_sum[0][12][0];
assign out_fmap[0][13] = xor_sum[0][13][0];
assign out_fmap[0][14] = xor_sum[0][14][0];
assign out_fmap[0][15] = xor_sum[0][15][0];
assign out_fmap[0][16] = xor_sum[0][16][0];
assign out_fmap[0][17] = xor_sum[0][17][0];
assign out_fmap[0][18] = xor_sum[0][18][0];
assign out_fmap[0][19] = xor_sum[0][19][0];
assign out_fmap[0][20] = xor_sum[0][20][0];
assign out_fmap[0][21] = xor_sum[0][21][0];
assign out_fmap[0][22] = xor_sum[0][22][0];
assign out_fmap[0][23] = xor_sum[0][23][0];
assign out_fmap[1][0] = xor_sum[1][0][0];
assign out_fmap[1][1] = xor_sum[1][1][0];
assign out_fmap[1][2] = xor_sum[1][2][0];
assign out_fmap[1][3] = xor_sum[1][3][0];
assign out_fmap[1][4] = xor_sum[1][4][0];
assign out_fmap[1][5] = xor_sum[1][5][0];
assign out_fmap[1][6] = xor_sum[1][6][0];
assign out_fmap[1][7] = xor_sum[1][7][0];
assign out_fmap[1][8] = xor_sum[1][8][0];
assign out_fmap[1][9] = xor_sum[1][9][0];
assign out_fmap[1][10] = xor_sum[1][10][0];
assign out_fmap[1][11] = xor_sum[1][11][0];
assign out_fmap[1][12] = xor_sum[1][12][0];
assign out_fmap[1][13] = xor_sum[1][13][0];
assign out_fmap[1][14] = xor_sum[1][14][0];
assign out_fmap[1][15] = xor_sum[1][15][0];
assign out_fmap[1][16] = xor_sum[1][16][0];
assign out_fmap[1][17] = xor_sum[1][17][0];
assign out_fmap[1][18] = xor_sum[1][18][0];
assign out_fmap[1][19] = xor_sum[1][19][0];
assign out_fmap[1][20] = xor_sum[1][20][0];
assign out_fmap[1][21] = xor_sum[1][21][0];
assign out_fmap[1][22] = xor_sum[1][22][0];
assign out_fmap[1][23] = xor_sum[1][23][0];
assign out_fmap[2][0] = xor_sum[2][0][0];
assign out_fmap[2][1] = xor_sum[2][1][0];
assign out_fmap[2][2] = xor_sum[2][2][0];
assign out_fmap[2][3] = xor_sum[2][3][0];
assign out_fmap[2][4] = xor_sum[2][4][0];
assign out_fmap[2][5] = xor_sum[2][5][0];
assign out_fmap[2][6] = xor_sum[2][6][0];
assign out_fmap[2][7] = xor_sum[2][7][0];
assign out_fmap[2][8] = xor_sum[2][8][0];
assign out_fmap[2][9] = xor_sum[2][9][0];
assign out_fmap[2][10] = xor_sum[2][10][0];
assign out_fmap[2][11] = xor_sum[2][11][0];
assign out_fmap[2][12] = xor_sum[2][12][0];
assign out_fmap[2][13] = xor_sum[2][13][0];
assign out_fmap[2][14] = xor_sum[2][14][0];
assign out_fmap[2][15] = xor_sum[2][15][0];
assign out_fmap[2][16] = xor_sum[2][16][0];
assign out_fmap[2][17] = xor_sum[2][17][0];
assign out_fmap[2][18] = xor_sum[2][18][0];
assign out_fmap[2][19] = xor_sum[2][19][0];
assign out_fmap[2][20] = xor_sum[2][20][0];
assign out_fmap[2][21] = xor_sum[2][21][0];
assign out_fmap[2][22] = xor_sum[2][22][0];
assign out_fmap[2][23] = xor_sum[2][23][0];
assign out_fmap[3][0] = xor_sum[3][0][0];
assign out_fmap[3][1] = xor_sum[3][1][0];
assign out_fmap[3][2] = xor_sum[3][2][0];
assign out_fmap[3][3] = xor_sum[3][3][0];
assign out_fmap[3][4] = xor_sum[3][4][0];
assign out_fmap[3][5] = xor_sum[3][5][0];
assign out_fmap[3][6] = xor_sum[3][6][0];
assign out_fmap[3][7] = xor_sum[3][7][0];
assign out_fmap[3][8] = xor_sum[3][8][0];
assign out_fmap[3][9] = xor_sum[3][9][0];
assign out_fmap[3][10] = xor_sum[3][10][0];
assign out_fmap[3][11] = xor_sum[3][11][0];
assign out_fmap[3][12] = xor_sum[3][12][0];
assign out_fmap[3][13] = xor_sum[3][13][0];
assign out_fmap[3][14] = xor_sum[3][14][0];
assign out_fmap[3][15] = xor_sum[3][15][0];
assign out_fmap[3][16] = xor_sum[3][16][0];
assign out_fmap[3][17] = xor_sum[3][17][0];
assign out_fmap[3][18] = xor_sum[3][18][0];
assign out_fmap[3][19] = xor_sum[3][19][0];
assign out_fmap[3][20] = xor_sum[3][20][0];
assign out_fmap[3][21] = xor_sum[3][21][0];
assign out_fmap[3][22] = xor_sum[3][22][0];
assign out_fmap[3][23] = xor_sum[3][23][0];
assign out_fmap[4][0] = xor_sum[4][0][0];
assign out_fmap[4][1] = xor_sum[4][1][0];
assign out_fmap[4][2] = xor_sum[4][2][0];
assign out_fmap[4][3] = xor_sum[4][3][0];
assign out_fmap[4][4] = xor_sum[4][4][0];
assign out_fmap[4][5] = xor_sum[4][5][0];
assign out_fmap[4][6] = xor_sum[4][6][0];
assign out_fmap[4][7] = xor_sum[4][7][0];
assign out_fmap[4][8] = xor_sum[4][8][0];
assign out_fmap[4][9] = xor_sum[4][9][0];
assign out_fmap[4][10] = xor_sum[4][10][0];
assign out_fmap[4][11] = xor_sum[4][11][0];
assign out_fmap[4][12] = xor_sum[4][12][0];
assign out_fmap[4][13] = xor_sum[4][13][0];
assign out_fmap[4][14] = xor_sum[4][14][0];
assign out_fmap[4][15] = xor_sum[4][15][0];
assign out_fmap[4][16] = xor_sum[4][16][0];
assign out_fmap[4][17] = xor_sum[4][17][0];
assign out_fmap[4][18] = xor_sum[4][18][0];
assign out_fmap[4][19] = xor_sum[4][19][0];
assign out_fmap[4][20] = xor_sum[4][20][0];
assign out_fmap[4][21] = xor_sum[4][21][0];
assign out_fmap[4][22] = xor_sum[4][22][0];
assign out_fmap[4][23] = xor_sum[4][23][0];
assign out_fmap[5][0] = xor_sum[5][0][0];
assign out_fmap[5][1] = xor_sum[5][1][0];
assign out_fmap[5][2] = xor_sum[5][2][0];
assign out_fmap[5][3] = xor_sum[5][3][0];
assign out_fmap[5][4] = xor_sum[5][4][0];
assign out_fmap[5][5] = xor_sum[5][5][0];
assign out_fmap[5][6] = xor_sum[5][6][0];
assign out_fmap[5][7] = xor_sum[5][7][0];
assign out_fmap[5][8] = xor_sum[5][8][0];
assign out_fmap[5][9] = xor_sum[5][9][0];
assign out_fmap[5][10] = xor_sum[5][10][0];
assign out_fmap[5][11] = xor_sum[5][11][0];
assign out_fmap[5][12] = xor_sum[5][12][0];
assign out_fmap[5][13] = xor_sum[5][13][0];
assign out_fmap[5][14] = xor_sum[5][14][0];
assign out_fmap[5][15] = xor_sum[5][15][0];
assign out_fmap[5][16] = xor_sum[5][16][0];
assign out_fmap[5][17] = xor_sum[5][17][0];
assign out_fmap[5][18] = xor_sum[5][18][0];
assign out_fmap[5][19] = xor_sum[5][19][0];
assign out_fmap[5][20] = xor_sum[5][20][0];
assign out_fmap[5][21] = xor_sum[5][21][0];
assign out_fmap[5][22] = xor_sum[5][22][0];
assign out_fmap[5][23] = xor_sum[5][23][0];
assign out_fmap[6][0] = xor_sum[6][0][0];
assign out_fmap[6][1] = xor_sum[6][1][0];
assign out_fmap[6][2] = xor_sum[6][2][0];
assign out_fmap[6][3] = xor_sum[6][3][0];
assign out_fmap[6][4] = xor_sum[6][4][0];
assign out_fmap[6][5] = xor_sum[6][5][0];
assign out_fmap[6][6] = xor_sum[6][6][0];
assign out_fmap[6][7] = xor_sum[6][7][0];
assign out_fmap[6][8] = xor_sum[6][8][0];
assign out_fmap[6][9] = xor_sum[6][9][0];
assign out_fmap[6][10] = xor_sum[6][10][0];
assign out_fmap[6][11] = xor_sum[6][11][0];
assign out_fmap[6][12] = xor_sum[6][12][0];
assign out_fmap[6][13] = xor_sum[6][13][0];
assign out_fmap[6][14] = xor_sum[6][14][0];
assign out_fmap[6][15] = xor_sum[6][15][0];
assign out_fmap[6][16] = xor_sum[6][16][0];
assign out_fmap[6][17] = xor_sum[6][17][0];
assign out_fmap[6][18] = xor_sum[6][18][0];
assign out_fmap[6][19] = xor_sum[6][19][0];
assign out_fmap[6][20] = xor_sum[6][20][0];
assign out_fmap[6][21] = xor_sum[6][21][0];
assign out_fmap[6][22] = xor_sum[6][22][0];
assign out_fmap[6][23] = xor_sum[6][23][0];
assign out_fmap[7][0] = xor_sum[7][0][0];
assign out_fmap[7][1] = xor_sum[7][1][0];
assign out_fmap[7][2] = xor_sum[7][2][0];
assign out_fmap[7][3] = xor_sum[7][3][0];
assign out_fmap[7][4] = xor_sum[7][4][0];
assign out_fmap[7][5] = xor_sum[7][5][0];
assign out_fmap[7][6] = xor_sum[7][6][0];
assign out_fmap[7][7] = xor_sum[7][7][0];
assign out_fmap[7][8] = xor_sum[7][8][0];
assign out_fmap[7][9] = xor_sum[7][9][0];
assign out_fmap[7][10] = xor_sum[7][10][0];
assign out_fmap[7][11] = xor_sum[7][11][0];
assign out_fmap[7][12] = xor_sum[7][12][0];
assign out_fmap[7][13] = xor_sum[7][13][0];
assign out_fmap[7][14] = xor_sum[7][14][0];
assign out_fmap[7][15] = xor_sum[7][15][0];
assign out_fmap[7][16] = xor_sum[7][16][0];
assign out_fmap[7][17] = xor_sum[7][17][0];
assign out_fmap[7][18] = xor_sum[7][18][0];
assign out_fmap[7][19] = xor_sum[7][19][0];
assign out_fmap[7][20] = xor_sum[7][20][0];
assign out_fmap[7][21] = xor_sum[7][21][0];
assign out_fmap[7][22] = xor_sum[7][22][0];
assign out_fmap[7][23] = xor_sum[7][23][0];
assign out_fmap[8][0] = xor_sum[8][0][0];
assign out_fmap[8][1] = xor_sum[8][1][0];
assign out_fmap[8][2] = xor_sum[8][2][0];
assign out_fmap[8][3] = xor_sum[8][3][0];
assign out_fmap[8][4] = xor_sum[8][4][0];
assign out_fmap[8][5] = xor_sum[8][5][0];
assign out_fmap[8][6] = xor_sum[8][6][0];
assign out_fmap[8][7] = xor_sum[8][7][0];
assign out_fmap[8][8] = xor_sum[8][8][0];
assign out_fmap[8][9] = xor_sum[8][9][0];
assign out_fmap[8][10] = xor_sum[8][10][0];
assign out_fmap[8][11] = xor_sum[8][11][0];
assign out_fmap[8][12] = xor_sum[8][12][0];
assign out_fmap[8][13] = xor_sum[8][13][0];
assign out_fmap[8][14] = xor_sum[8][14][0];
assign out_fmap[8][15] = xor_sum[8][15][0];
assign out_fmap[8][16] = xor_sum[8][16][0];
assign out_fmap[8][17] = xor_sum[8][17][0];
assign out_fmap[8][18] = xor_sum[8][18][0];
assign out_fmap[8][19] = xor_sum[8][19][0];
assign out_fmap[8][20] = xor_sum[8][20][0];
assign out_fmap[8][21] = xor_sum[8][21][0];
assign out_fmap[8][22] = xor_sum[8][22][0];
assign out_fmap[8][23] = xor_sum[8][23][0];
assign out_fmap[9][0] = xor_sum[9][0][0];
assign out_fmap[9][1] = xor_sum[9][1][0];
assign out_fmap[9][2] = xor_sum[9][2][0];
assign out_fmap[9][3] = xor_sum[9][3][0];
assign out_fmap[9][4] = xor_sum[9][4][0];
assign out_fmap[9][5] = xor_sum[9][5][0];
assign out_fmap[9][6] = xor_sum[9][6][0];
assign out_fmap[9][7] = xor_sum[9][7][0];
assign out_fmap[9][8] = xor_sum[9][8][0];
assign out_fmap[9][9] = xor_sum[9][9][0];
assign out_fmap[9][10] = xor_sum[9][10][0];
assign out_fmap[9][11] = xor_sum[9][11][0];
assign out_fmap[9][12] = xor_sum[9][12][0];
assign out_fmap[9][13] = xor_sum[9][13][0];
assign out_fmap[9][14] = xor_sum[9][14][0];
assign out_fmap[9][15] = xor_sum[9][15][0];
assign out_fmap[9][16] = xor_sum[9][16][0];
assign out_fmap[9][17] = xor_sum[9][17][0];
assign out_fmap[9][18] = xor_sum[9][18][0];
assign out_fmap[9][19] = xor_sum[9][19][0];
assign out_fmap[9][20] = xor_sum[9][20][0];
assign out_fmap[9][21] = xor_sum[9][21][0];
assign out_fmap[9][22] = xor_sum[9][22][0];
assign out_fmap[9][23] = xor_sum[9][23][0];
assign out_fmap[10][0] = xor_sum[10][0][0];
assign out_fmap[10][1] = xor_sum[10][1][0];
assign out_fmap[10][2] = xor_sum[10][2][0];
assign out_fmap[10][3] = xor_sum[10][3][0];
assign out_fmap[10][4] = xor_sum[10][4][0];
assign out_fmap[10][5] = xor_sum[10][5][0];
assign out_fmap[10][6] = xor_sum[10][6][0];
assign out_fmap[10][7] = xor_sum[10][7][0];
assign out_fmap[10][8] = xor_sum[10][8][0];
assign out_fmap[10][9] = xor_sum[10][9][0];
assign out_fmap[10][10] = xor_sum[10][10][0];
assign out_fmap[10][11] = xor_sum[10][11][0];
assign out_fmap[10][12] = xor_sum[10][12][0];
assign out_fmap[10][13] = xor_sum[10][13][0];
assign out_fmap[10][14] = xor_sum[10][14][0];
assign out_fmap[10][15] = xor_sum[10][15][0];
assign out_fmap[10][16] = xor_sum[10][16][0];
assign out_fmap[10][17] = xor_sum[10][17][0];
assign out_fmap[10][18] = xor_sum[10][18][0];
assign out_fmap[10][19] = xor_sum[10][19][0];
assign out_fmap[10][20] = xor_sum[10][20][0];
assign out_fmap[10][21] = xor_sum[10][21][0];
assign out_fmap[10][22] = xor_sum[10][22][0];
assign out_fmap[10][23] = xor_sum[10][23][0];
assign out_fmap[11][0] = xor_sum[11][0][0];
assign out_fmap[11][1] = xor_sum[11][1][0];
assign out_fmap[11][2] = xor_sum[11][2][0];
assign out_fmap[11][3] = xor_sum[11][3][0];
assign out_fmap[11][4] = xor_sum[11][4][0];
assign out_fmap[11][5] = xor_sum[11][5][0];
assign out_fmap[11][6] = xor_sum[11][6][0];
assign out_fmap[11][7] = xor_sum[11][7][0];
assign out_fmap[11][8] = xor_sum[11][8][0];
assign out_fmap[11][9] = xor_sum[11][9][0];
assign out_fmap[11][10] = xor_sum[11][10][0];
assign out_fmap[11][11] = xor_sum[11][11][0];
assign out_fmap[11][12] = xor_sum[11][12][0];
assign out_fmap[11][13] = xor_sum[11][13][0];
assign out_fmap[11][14] = xor_sum[11][14][0];
assign out_fmap[11][15] = xor_sum[11][15][0];
assign out_fmap[11][16] = xor_sum[11][16][0];
assign out_fmap[11][17] = xor_sum[11][17][0];
assign out_fmap[11][18] = xor_sum[11][18][0];
assign out_fmap[11][19] = xor_sum[11][19][0];
assign out_fmap[11][20] = xor_sum[11][20][0];
assign out_fmap[11][21] = xor_sum[11][21][0];
assign out_fmap[11][22] = xor_sum[11][22][0];
assign out_fmap[11][23] = xor_sum[11][23][0];
assign out_fmap[12][0] = xor_sum[12][0][0];
assign out_fmap[12][1] = xor_sum[12][1][0];
assign out_fmap[12][2] = xor_sum[12][2][0];
assign out_fmap[12][3] = xor_sum[12][3][0];
assign out_fmap[12][4] = xor_sum[12][4][0];
assign out_fmap[12][5] = xor_sum[12][5][0];
assign out_fmap[12][6] = xor_sum[12][6][0];
assign out_fmap[12][7] = xor_sum[12][7][0];
assign out_fmap[12][8] = xor_sum[12][8][0];
assign out_fmap[12][9] = xor_sum[12][9][0];
assign out_fmap[12][10] = xor_sum[12][10][0];
assign out_fmap[12][11] = xor_sum[12][11][0];
assign out_fmap[12][12] = xor_sum[12][12][0];
assign out_fmap[12][13] = xor_sum[12][13][0];
assign out_fmap[12][14] = xor_sum[12][14][0];
assign out_fmap[12][15] = xor_sum[12][15][0];
assign out_fmap[12][16] = xor_sum[12][16][0];
assign out_fmap[12][17] = xor_sum[12][17][0];
assign out_fmap[12][18] = xor_sum[12][18][0];
assign out_fmap[12][19] = xor_sum[12][19][0];
assign out_fmap[12][20] = xor_sum[12][20][0];
assign out_fmap[12][21] = xor_sum[12][21][0];
assign out_fmap[12][22] = xor_sum[12][22][0];
assign out_fmap[12][23] = xor_sum[12][23][0];
assign out_fmap[13][0] = xor_sum[13][0][0];
assign out_fmap[13][1] = xor_sum[13][1][0];
assign out_fmap[13][2] = xor_sum[13][2][0];
assign out_fmap[13][3] = xor_sum[13][3][0];
assign out_fmap[13][4] = xor_sum[13][4][0];
assign out_fmap[13][5] = xor_sum[13][5][0];
assign out_fmap[13][6] = xor_sum[13][6][0];
assign out_fmap[13][7] = xor_sum[13][7][0];
assign out_fmap[13][8] = xor_sum[13][8][0];
assign out_fmap[13][9] = xor_sum[13][9][0];
assign out_fmap[13][10] = xor_sum[13][10][0];
assign out_fmap[13][11] = xor_sum[13][11][0];
assign out_fmap[13][12] = xor_sum[13][12][0];
assign out_fmap[13][13] = xor_sum[13][13][0];
assign out_fmap[13][14] = xor_sum[13][14][0];
assign out_fmap[13][15] = xor_sum[13][15][0];
assign out_fmap[13][16] = xor_sum[13][16][0];
assign out_fmap[13][17] = xor_sum[13][17][0];
assign out_fmap[13][18] = xor_sum[13][18][0];
assign out_fmap[13][19] = xor_sum[13][19][0];
assign out_fmap[13][20] = xor_sum[13][20][0];
assign out_fmap[13][21] = xor_sum[13][21][0];
assign out_fmap[13][22] = xor_sum[13][22][0];
assign out_fmap[13][23] = xor_sum[13][23][0];
assign out_fmap[14][0] = xor_sum[14][0][0];
assign out_fmap[14][1] = xor_sum[14][1][0];
assign out_fmap[14][2] = xor_sum[14][2][0];
assign out_fmap[14][3] = xor_sum[14][3][0];
assign out_fmap[14][4] = xor_sum[14][4][0];
assign out_fmap[14][5] = xor_sum[14][5][0];
assign out_fmap[14][6] = xor_sum[14][6][0];
assign out_fmap[14][7] = xor_sum[14][7][0];
assign out_fmap[14][8] = xor_sum[14][8][0];
assign out_fmap[14][9] = xor_sum[14][9][0];
assign out_fmap[14][10] = xor_sum[14][10][0];
assign out_fmap[14][11] = xor_sum[14][11][0];
assign out_fmap[14][12] = xor_sum[14][12][0];
assign out_fmap[14][13] = xor_sum[14][13][0];
assign out_fmap[14][14] = xor_sum[14][14][0];
assign out_fmap[14][15] = xor_sum[14][15][0];
assign out_fmap[14][16] = xor_sum[14][16][0];
assign out_fmap[14][17] = xor_sum[14][17][0];
assign out_fmap[14][18] = xor_sum[14][18][0];
assign out_fmap[14][19] = xor_sum[14][19][0];
assign out_fmap[14][20] = xor_sum[14][20][0];
assign out_fmap[14][21] = xor_sum[14][21][0];
assign out_fmap[14][22] = xor_sum[14][22][0];
assign out_fmap[14][23] = xor_sum[14][23][0];
assign out_fmap[15][0] = xor_sum[15][0][0];
assign out_fmap[15][1] = xor_sum[15][1][0];
assign out_fmap[15][2] = xor_sum[15][2][0];
assign out_fmap[15][3] = xor_sum[15][3][0];
assign out_fmap[15][4] = xor_sum[15][4][0];
assign out_fmap[15][5] = xor_sum[15][5][0];
assign out_fmap[15][6] = xor_sum[15][6][0];
assign out_fmap[15][7] = xor_sum[15][7][0];
assign out_fmap[15][8] = xor_sum[15][8][0];
assign out_fmap[15][9] = xor_sum[15][9][0];
assign out_fmap[15][10] = xor_sum[15][10][0];
assign out_fmap[15][11] = xor_sum[15][11][0];
assign out_fmap[15][12] = xor_sum[15][12][0];
assign out_fmap[15][13] = xor_sum[15][13][0];
assign out_fmap[15][14] = xor_sum[15][14][0];
assign out_fmap[15][15] = xor_sum[15][15][0];
assign out_fmap[15][16] = xor_sum[15][16][0];
assign out_fmap[15][17] = xor_sum[15][17][0];
assign out_fmap[15][18] = xor_sum[15][18][0];
assign out_fmap[15][19] = xor_sum[15][19][0];
assign out_fmap[15][20] = xor_sum[15][20][0];
assign out_fmap[15][21] = xor_sum[15][21][0];
assign out_fmap[15][22] = xor_sum[15][22][0];
assign out_fmap[15][23] = xor_sum[15][23][0];
assign out_fmap[16][0] = xor_sum[16][0][0];
assign out_fmap[16][1] = xor_sum[16][1][0];
assign out_fmap[16][2] = xor_sum[16][2][0];
assign out_fmap[16][3] = xor_sum[16][3][0];
assign out_fmap[16][4] = xor_sum[16][4][0];
assign out_fmap[16][5] = xor_sum[16][5][0];
assign out_fmap[16][6] = xor_sum[16][6][0];
assign out_fmap[16][7] = xor_sum[16][7][0];
assign out_fmap[16][8] = xor_sum[16][8][0];
assign out_fmap[16][9] = xor_sum[16][9][0];
assign out_fmap[16][10] = xor_sum[16][10][0];
assign out_fmap[16][11] = xor_sum[16][11][0];
assign out_fmap[16][12] = xor_sum[16][12][0];
assign out_fmap[16][13] = xor_sum[16][13][0];
assign out_fmap[16][14] = xor_sum[16][14][0];
assign out_fmap[16][15] = xor_sum[16][15][0];
assign out_fmap[16][16] = xor_sum[16][16][0];
assign out_fmap[16][17] = xor_sum[16][17][0];
assign out_fmap[16][18] = xor_sum[16][18][0];
assign out_fmap[16][19] = xor_sum[16][19][0];
assign out_fmap[16][20] = xor_sum[16][20][0];
assign out_fmap[16][21] = xor_sum[16][21][0];
assign out_fmap[16][22] = xor_sum[16][22][0];
assign out_fmap[16][23] = xor_sum[16][23][0];
assign out_fmap[17][0] = xor_sum[17][0][0];
assign out_fmap[17][1] = xor_sum[17][1][0];
assign out_fmap[17][2] = xor_sum[17][2][0];
assign out_fmap[17][3] = xor_sum[17][3][0];
assign out_fmap[17][4] = xor_sum[17][4][0];
assign out_fmap[17][5] = xor_sum[17][5][0];
assign out_fmap[17][6] = xor_sum[17][6][0];
assign out_fmap[17][7] = xor_sum[17][7][0];
assign out_fmap[17][8] = xor_sum[17][8][0];
assign out_fmap[17][9] = xor_sum[17][9][0];
assign out_fmap[17][10] = xor_sum[17][10][0];
assign out_fmap[17][11] = xor_sum[17][11][0];
assign out_fmap[17][12] = xor_sum[17][12][0];
assign out_fmap[17][13] = xor_sum[17][13][0];
assign out_fmap[17][14] = xor_sum[17][14][0];
assign out_fmap[17][15] = xor_sum[17][15][0];
assign out_fmap[17][16] = xor_sum[17][16][0];
assign out_fmap[17][17] = xor_sum[17][17][0];
assign out_fmap[17][18] = xor_sum[17][18][0];
assign out_fmap[17][19] = xor_sum[17][19][0];
assign out_fmap[17][20] = xor_sum[17][20][0];
assign out_fmap[17][21] = xor_sum[17][21][0];
assign out_fmap[17][22] = xor_sum[17][22][0];
assign out_fmap[17][23] = xor_sum[17][23][0];
assign out_fmap[18][0] = xor_sum[18][0][0];
assign out_fmap[18][1] = xor_sum[18][1][0];
assign out_fmap[18][2] = xor_sum[18][2][0];
assign out_fmap[18][3] = xor_sum[18][3][0];
assign out_fmap[18][4] = xor_sum[18][4][0];
assign out_fmap[18][5] = xor_sum[18][5][0];
assign out_fmap[18][6] = xor_sum[18][6][0];
assign out_fmap[18][7] = xor_sum[18][7][0];
assign out_fmap[18][8] = xor_sum[18][8][0];
assign out_fmap[18][9] = xor_sum[18][9][0];
assign out_fmap[18][10] = xor_sum[18][10][0];
assign out_fmap[18][11] = xor_sum[18][11][0];
assign out_fmap[18][12] = xor_sum[18][12][0];
assign out_fmap[18][13] = xor_sum[18][13][0];
assign out_fmap[18][14] = xor_sum[18][14][0];
assign out_fmap[18][15] = xor_sum[18][15][0];
assign out_fmap[18][16] = xor_sum[18][16][0];
assign out_fmap[18][17] = xor_sum[18][17][0];
assign out_fmap[18][18] = xor_sum[18][18][0];
assign out_fmap[18][19] = xor_sum[18][19][0];
assign out_fmap[18][20] = xor_sum[18][20][0];
assign out_fmap[18][21] = xor_sum[18][21][0];
assign out_fmap[18][22] = xor_sum[18][22][0];
assign out_fmap[18][23] = xor_sum[18][23][0];
assign out_fmap[19][0] = xor_sum[19][0][0];
assign out_fmap[19][1] = xor_sum[19][1][0];
assign out_fmap[19][2] = xor_sum[19][2][0];
assign out_fmap[19][3] = xor_sum[19][3][0];
assign out_fmap[19][4] = xor_sum[19][4][0];
assign out_fmap[19][5] = xor_sum[19][5][0];
assign out_fmap[19][6] = xor_sum[19][6][0];
assign out_fmap[19][7] = xor_sum[19][7][0];
assign out_fmap[19][8] = xor_sum[19][8][0];
assign out_fmap[19][9] = xor_sum[19][9][0];
assign out_fmap[19][10] = xor_sum[19][10][0];
assign out_fmap[19][11] = xor_sum[19][11][0];
assign out_fmap[19][12] = xor_sum[19][12][0];
assign out_fmap[19][13] = xor_sum[19][13][0];
assign out_fmap[19][14] = xor_sum[19][14][0];
assign out_fmap[19][15] = xor_sum[19][15][0];
assign out_fmap[19][16] = xor_sum[19][16][0];
assign out_fmap[19][17] = xor_sum[19][17][0];
assign out_fmap[19][18] = xor_sum[19][18][0];
assign out_fmap[19][19] = xor_sum[19][19][0];
assign out_fmap[19][20] = xor_sum[19][20][0];
assign out_fmap[19][21] = xor_sum[19][21][0];
assign out_fmap[19][22] = xor_sum[19][22][0];
assign out_fmap[19][23] = xor_sum[19][23][0];
assign out_fmap[20][0] = xor_sum[20][0][0];
assign out_fmap[20][1] = xor_sum[20][1][0];
assign out_fmap[20][2] = xor_sum[20][2][0];
assign out_fmap[20][3] = xor_sum[20][3][0];
assign out_fmap[20][4] = xor_sum[20][4][0];
assign out_fmap[20][5] = xor_sum[20][5][0];
assign out_fmap[20][6] = xor_sum[20][6][0];
assign out_fmap[20][7] = xor_sum[20][7][0];
assign out_fmap[20][8] = xor_sum[20][8][0];
assign out_fmap[20][9] = xor_sum[20][9][0];
assign out_fmap[20][10] = xor_sum[20][10][0];
assign out_fmap[20][11] = xor_sum[20][11][0];
assign out_fmap[20][12] = xor_sum[20][12][0];
assign out_fmap[20][13] = xor_sum[20][13][0];
assign out_fmap[20][14] = xor_sum[20][14][0];
assign out_fmap[20][15] = xor_sum[20][15][0];
assign out_fmap[20][16] = xor_sum[20][16][0];
assign out_fmap[20][17] = xor_sum[20][17][0];
assign out_fmap[20][18] = xor_sum[20][18][0];
assign out_fmap[20][19] = xor_sum[20][19][0];
assign out_fmap[20][20] = xor_sum[20][20][0];
assign out_fmap[20][21] = xor_sum[20][21][0];
assign out_fmap[20][22] = xor_sum[20][22][0];
assign out_fmap[20][23] = xor_sum[20][23][0];
assign out_fmap[21][0] = xor_sum[21][0][0];
assign out_fmap[21][1] = xor_sum[21][1][0];
assign out_fmap[21][2] = xor_sum[21][2][0];
assign out_fmap[21][3] = xor_sum[21][3][0];
assign out_fmap[21][4] = xor_sum[21][4][0];
assign out_fmap[21][5] = xor_sum[21][5][0];
assign out_fmap[21][6] = xor_sum[21][6][0];
assign out_fmap[21][7] = xor_sum[21][7][0];
assign out_fmap[21][8] = xor_sum[21][8][0];
assign out_fmap[21][9] = xor_sum[21][9][0];
assign out_fmap[21][10] = xor_sum[21][10][0];
assign out_fmap[21][11] = xor_sum[21][11][0];
assign out_fmap[21][12] = xor_sum[21][12][0];
assign out_fmap[21][13] = xor_sum[21][13][0];
assign out_fmap[21][14] = xor_sum[21][14][0];
assign out_fmap[21][15] = xor_sum[21][15][0];
assign out_fmap[21][16] = xor_sum[21][16][0];
assign out_fmap[21][17] = xor_sum[21][17][0];
assign out_fmap[21][18] = xor_sum[21][18][0];
assign out_fmap[21][19] = xor_sum[21][19][0];
assign out_fmap[21][20] = xor_sum[21][20][0];
assign out_fmap[21][21] = xor_sum[21][21][0];
assign out_fmap[21][22] = xor_sum[21][22][0];
assign out_fmap[21][23] = xor_sum[21][23][0];
assign out_fmap[22][0] = xor_sum[22][0][0];
assign out_fmap[22][1] = xor_sum[22][1][0];
assign out_fmap[22][2] = xor_sum[22][2][0];
assign out_fmap[22][3] = xor_sum[22][3][0];
assign out_fmap[22][4] = xor_sum[22][4][0];
assign out_fmap[22][5] = xor_sum[22][5][0];
assign out_fmap[22][6] = xor_sum[22][6][0];
assign out_fmap[22][7] = xor_sum[22][7][0];
assign out_fmap[22][8] = xor_sum[22][8][0];
assign out_fmap[22][9] = xor_sum[22][9][0];
assign out_fmap[22][10] = xor_sum[22][10][0];
assign out_fmap[22][11] = xor_sum[22][11][0];
assign out_fmap[22][12] = xor_sum[22][12][0];
assign out_fmap[22][13] = xor_sum[22][13][0];
assign out_fmap[22][14] = xor_sum[22][14][0];
assign out_fmap[22][15] = xor_sum[22][15][0];
assign out_fmap[22][16] = xor_sum[22][16][0];
assign out_fmap[22][17] = xor_sum[22][17][0];
assign out_fmap[22][18] = xor_sum[22][18][0];
assign out_fmap[22][19] = xor_sum[22][19][0];
assign out_fmap[22][20] = xor_sum[22][20][0];
assign out_fmap[22][21] = xor_sum[22][21][0];
assign out_fmap[22][22] = xor_sum[22][22][0];
assign out_fmap[22][23] = xor_sum[22][23][0];
assign out_fmap[23][0] = xor_sum[23][0][0];
assign out_fmap[23][1] = xor_sum[23][1][0];
assign out_fmap[23][2] = xor_sum[23][2][0];
assign out_fmap[23][3] = xor_sum[23][3][0];
assign out_fmap[23][4] = xor_sum[23][4][0];
assign out_fmap[23][5] = xor_sum[23][5][0];
assign out_fmap[23][6] = xor_sum[23][6][0];
assign out_fmap[23][7] = xor_sum[23][7][0];
assign out_fmap[23][8] = xor_sum[23][8][0];
assign out_fmap[23][9] = xor_sum[23][9][0];
assign out_fmap[23][10] = xor_sum[23][10][0];
assign out_fmap[23][11] = xor_sum[23][11][0];
assign out_fmap[23][12] = xor_sum[23][12][0];
assign out_fmap[23][13] = xor_sum[23][13][0];
assign out_fmap[23][14] = xor_sum[23][14][0];
assign out_fmap[23][15] = xor_sum[23][15][0];
assign out_fmap[23][16] = xor_sum[23][16][0];
assign out_fmap[23][17] = xor_sum[23][17][0];
assign out_fmap[23][18] = xor_sum[23][18][0];
assign out_fmap[23][19] = xor_sum[23][19][0];
assign out_fmap[23][20] = xor_sum[23][20][0];
assign out_fmap[23][21] = xor_sum[23][21][0];
assign out_fmap[23][22] = xor_sum[23][22][0];
assign out_fmap[23][23] = xor_sum[23][23][0];

endmodule