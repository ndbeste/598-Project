module convchan1 
    #( parameter bW = 8 )
    ( 
    input  logic          image     [0:27][0:27],
    input  logic          kernel    [0:4] [0:4],
    output logic [bW-1:0] out_fmap  [0:23][0:23]
    );

assign xor_sum[0][0] = kernel[0][0] ~^ image[0][0] + kernel[0][1] ~^ image[0][1] + kernel[0][2] ~^ image[0][2] + kernel[0][3] ~^ image[0][3] + kernel[0][4] ~^ image[0][4] + kernel[1][0] ~^ image[1][0] + kernel[1][1] ~^ image[1][1] + kernel[1][2] ~^ image[1][2] + kernel[1][3] ~^ image[1][3] + kernel[1][4] ~^ image[1][4] + kernel[2][0] ~^ image[2][0] + kernel[2][1] ~^ image[2][1] + kernel[2][2] ~^ image[2][2] + kernel[2][3] ~^ image[2][3] + kernel[2][4] ~^ image[2][4] + kernel[3][0] ~^ image[3][0] + kernel[3][1] ~^ image[3][1] + kernel[3][2] ~^ image[3][2] + kernel[3][3] ~^ image[3][3] + kernel[3][4] ~^ image[3][4] + kernel[4][0] ~^ image[4][0] + kernel[4][1] ~^ image[4][1] + kernel[4][2] ~^ image[4][2] + kernel[4][3] ~^ image[4][3] + kernel[4][4] ~^ image[4][4];
assign xor_sum[0][1] = kernel[0][0] ~^ image[0][1] + kernel[0][1] ~^ image[0][2] + kernel[0][2] ~^ image[0][3] + kernel[0][3] ~^ image[0][4] + kernel[0][4] ~^ image[0][5] + kernel[1][0] ~^ image[1][1] + kernel[1][1] ~^ image[1][2] + kernel[1][2] ~^ image[1][3] + kernel[1][3] ~^ image[1][4] + kernel[1][4] ~^ image[1][5] + kernel[2][0] ~^ image[2][1] + kernel[2][1] ~^ image[2][2] + kernel[2][2] ~^ image[2][3] + kernel[2][3] ~^ image[2][4] + kernel[2][4] ~^ image[2][5] + kernel[3][0] ~^ image[3][1] + kernel[3][1] ~^ image[3][2] + kernel[3][2] ~^ image[3][3] + kernel[3][3] ~^ image[3][4] + kernel[3][4] ~^ image[3][5] + kernel[4][0] ~^ image[4][1] + kernel[4][1] ~^ image[4][2] + kernel[4][2] ~^ image[4][3] + kernel[4][3] ~^ image[4][4] + kernel[4][4] ~^ image[4][5];
assign xor_sum[0][2] = kernel[0][0] ~^ image[0][2] + kernel[0][1] ~^ image[0][3] + kernel[0][2] ~^ image[0][4] + kernel[0][3] ~^ image[0][5] + kernel[0][4] ~^ image[0][6] + kernel[1][0] ~^ image[1][2] + kernel[1][1] ~^ image[1][3] + kernel[1][2] ~^ image[1][4] + kernel[1][3] ~^ image[1][5] + kernel[1][4] ~^ image[1][6] + kernel[2][0] ~^ image[2][2] + kernel[2][1] ~^ image[2][3] + kernel[2][2] ~^ image[2][4] + kernel[2][3] ~^ image[2][5] + kernel[2][4] ~^ image[2][6] + kernel[3][0] ~^ image[3][2] + kernel[3][1] ~^ image[3][3] + kernel[3][2] ~^ image[3][4] + kernel[3][3] ~^ image[3][5] + kernel[3][4] ~^ image[3][6] + kernel[4][0] ~^ image[4][2] + kernel[4][1] ~^ image[4][3] + kernel[4][2] ~^ image[4][4] + kernel[4][3] ~^ image[4][5] + kernel[4][4] ~^ image[4][6];
assign xor_sum[0][3] = kernel[0][0] ~^ image[0][3] + kernel[0][1] ~^ image[0][4] + kernel[0][2] ~^ image[0][5] + kernel[0][3] ~^ image[0][6] + kernel[0][4] ~^ image[0][7] + kernel[1][0] ~^ image[1][3] + kernel[1][1] ~^ image[1][4] + kernel[1][2] ~^ image[1][5] + kernel[1][3] ~^ image[1][6] + kernel[1][4] ~^ image[1][7] + kernel[2][0] ~^ image[2][3] + kernel[2][1] ~^ image[2][4] + kernel[2][2] ~^ image[2][5] + kernel[2][3] ~^ image[2][6] + kernel[2][4] ~^ image[2][7] + kernel[3][0] ~^ image[3][3] + kernel[3][1] ~^ image[3][4] + kernel[3][2] ~^ image[3][5] + kernel[3][3] ~^ image[3][6] + kernel[3][4] ~^ image[3][7] + kernel[4][0] ~^ image[4][3] + kernel[4][1] ~^ image[4][4] + kernel[4][2] ~^ image[4][5] + kernel[4][3] ~^ image[4][6] + kernel[4][4] ~^ image[4][7];
assign xor_sum[0][4] = kernel[0][0] ~^ image[0][4] + kernel[0][1] ~^ image[0][5] + kernel[0][2] ~^ image[0][6] + kernel[0][3] ~^ image[0][7] + kernel[0][4] ~^ image[0][8] + kernel[1][0] ~^ image[1][4] + kernel[1][1] ~^ image[1][5] + kernel[1][2] ~^ image[1][6] + kernel[1][3] ~^ image[1][7] + kernel[1][4] ~^ image[1][8] + kernel[2][0] ~^ image[2][4] + kernel[2][1] ~^ image[2][5] + kernel[2][2] ~^ image[2][6] + kernel[2][3] ~^ image[2][7] + kernel[2][4] ~^ image[2][8] + kernel[3][0] ~^ image[3][4] + kernel[3][1] ~^ image[3][5] + kernel[3][2] ~^ image[3][6] + kernel[3][3] ~^ image[3][7] + kernel[3][4] ~^ image[3][8] + kernel[4][0] ~^ image[4][4] + kernel[4][1] ~^ image[4][5] + kernel[4][2] ~^ image[4][6] + kernel[4][3] ~^ image[4][7] + kernel[4][4] ~^ image[4][8];
assign xor_sum[0][5] = kernel[0][0] ~^ image[0][5] + kernel[0][1] ~^ image[0][6] + kernel[0][2] ~^ image[0][7] + kernel[0][3] ~^ image[0][8] + kernel[0][4] ~^ image[0][9] + kernel[1][0] ~^ image[1][5] + kernel[1][1] ~^ image[1][6] + kernel[1][2] ~^ image[1][7] + kernel[1][3] ~^ image[1][8] + kernel[1][4] ~^ image[1][9] + kernel[2][0] ~^ image[2][5] + kernel[2][1] ~^ image[2][6] + kernel[2][2] ~^ image[2][7] + kernel[2][3] ~^ image[2][8] + kernel[2][4] ~^ image[2][9] + kernel[3][0] ~^ image[3][5] + kernel[3][1] ~^ image[3][6] + kernel[3][2] ~^ image[3][7] + kernel[3][3] ~^ image[3][8] + kernel[3][4] ~^ image[3][9] + kernel[4][0] ~^ image[4][5] + kernel[4][1] ~^ image[4][6] + kernel[4][2] ~^ image[4][7] + kernel[4][3] ~^ image[4][8] + kernel[4][4] ~^ image[4][9];
assign xor_sum[0][6] = kernel[0][0] ~^ image[0][6] + kernel[0][1] ~^ image[0][7] + kernel[0][2] ~^ image[0][8] + kernel[0][3] ~^ image[0][9] + kernel[0][4] ~^ image[0][10] + kernel[1][0] ~^ image[1][6] + kernel[1][1] ~^ image[1][7] + kernel[1][2] ~^ image[1][8] + kernel[1][3] ~^ image[1][9] + kernel[1][4] ~^ image[1][10] + kernel[2][0] ~^ image[2][6] + kernel[2][1] ~^ image[2][7] + kernel[2][2] ~^ image[2][8] + kernel[2][3] ~^ image[2][9] + kernel[2][4] ~^ image[2][10] + kernel[3][0] ~^ image[3][6] + kernel[3][1] ~^ image[3][7] + kernel[3][2] ~^ image[3][8] + kernel[3][3] ~^ image[3][9] + kernel[3][4] ~^ image[3][10] + kernel[4][0] ~^ image[4][6] + kernel[4][1] ~^ image[4][7] + kernel[4][2] ~^ image[4][8] + kernel[4][3] ~^ image[4][9] + kernel[4][4] ~^ image[4][10];
assign xor_sum[0][7] = kernel[0][0] ~^ image[0][7] + kernel[0][1] ~^ image[0][8] + kernel[0][2] ~^ image[0][9] + kernel[0][3] ~^ image[0][10] + kernel[0][4] ~^ image[0][11] + kernel[1][0] ~^ image[1][7] + kernel[1][1] ~^ image[1][8] + kernel[1][2] ~^ image[1][9] + kernel[1][3] ~^ image[1][10] + kernel[1][4] ~^ image[1][11] + kernel[2][0] ~^ image[2][7] + kernel[2][1] ~^ image[2][8] + kernel[2][2] ~^ image[2][9] + kernel[2][3] ~^ image[2][10] + kernel[2][4] ~^ image[2][11] + kernel[3][0] ~^ image[3][7] + kernel[3][1] ~^ image[3][8] + kernel[3][2] ~^ image[3][9] + kernel[3][3] ~^ image[3][10] + kernel[3][4] ~^ image[3][11] + kernel[4][0] ~^ image[4][7] + kernel[4][1] ~^ image[4][8] + kernel[4][2] ~^ image[4][9] + kernel[4][3] ~^ image[4][10] + kernel[4][4] ~^ image[4][11];
assign xor_sum[0][8] = kernel[0][0] ~^ image[0][8] + kernel[0][1] ~^ image[0][9] + kernel[0][2] ~^ image[0][10] + kernel[0][3] ~^ image[0][11] + kernel[0][4] ~^ image[0][12] + kernel[1][0] ~^ image[1][8] + kernel[1][1] ~^ image[1][9] + kernel[1][2] ~^ image[1][10] + kernel[1][3] ~^ image[1][11] + kernel[1][4] ~^ image[1][12] + kernel[2][0] ~^ image[2][8] + kernel[2][1] ~^ image[2][9] + kernel[2][2] ~^ image[2][10] + kernel[2][3] ~^ image[2][11] + kernel[2][4] ~^ image[2][12] + kernel[3][0] ~^ image[3][8] + kernel[3][1] ~^ image[3][9] + kernel[3][2] ~^ image[3][10] + kernel[3][3] ~^ image[3][11] + kernel[3][4] ~^ image[3][12] + kernel[4][0] ~^ image[4][8] + kernel[4][1] ~^ image[4][9] + kernel[4][2] ~^ image[4][10] + kernel[4][3] ~^ image[4][11] + kernel[4][4] ~^ image[4][12];
assign xor_sum[0][9] = kernel[0][0] ~^ image[0][9] + kernel[0][1] ~^ image[0][10] + kernel[0][2] ~^ image[0][11] + kernel[0][3] ~^ image[0][12] + kernel[0][4] ~^ image[0][13] + kernel[1][0] ~^ image[1][9] + kernel[1][1] ~^ image[1][10] + kernel[1][2] ~^ image[1][11] + kernel[1][3] ~^ image[1][12] + kernel[1][4] ~^ image[1][13] + kernel[2][0] ~^ image[2][9] + kernel[2][1] ~^ image[2][10] + kernel[2][2] ~^ image[2][11] + kernel[2][3] ~^ image[2][12] + kernel[2][4] ~^ image[2][13] + kernel[3][0] ~^ image[3][9] + kernel[3][1] ~^ image[3][10] + kernel[3][2] ~^ image[3][11] + kernel[3][3] ~^ image[3][12] + kernel[3][4] ~^ image[3][13] + kernel[4][0] ~^ image[4][9] + kernel[4][1] ~^ image[4][10] + kernel[4][2] ~^ image[4][11] + kernel[4][3] ~^ image[4][12] + kernel[4][4] ~^ image[4][13];
assign xor_sum[0][10] = kernel[0][0] ~^ image[0][10] + kernel[0][1] ~^ image[0][11] + kernel[0][2] ~^ image[0][12] + kernel[0][3] ~^ image[0][13] + kernel[0][4] ~^ image[0][14] + kernel[1][0] ~^ image[1][10] + kernel[1][1] ~^ image[1][11] + kernel[1][2] ~^ image[1][12] + kernel[1][3] ~^ image[1][13] + kernel[1][4] ~^ image[1][14] + kernel[2][0] ~^ image[2][10] + kernel[2][1] ~^ image[2][11] + kernel[2][2] ~^ image[2][12] + kernel[2][3] ~^ image[2][13] + kernel[2][4] ~^ image[2][14] + kernel[3][0] ~^ image[3][10] + kernel[3][1] ~^ image[3][11] + kernel[3][2] ~^ image[3][12] + kernel[3][3] ~^ image[3][13] + kernel[3][4] ~^ image[3][14] + kernel[4][0] ~^ image[4][10] + kernel[4][1] ~^ image[4][11] + kernel[4][2] ~^ image[4][12] + kernel[4][3] ~^ image[4][13] + kernel[4][4] ~^ image[4][14];
assign xor_sum[0][11] = kernel[0][0] ~^ image[0][11] + kernel[0][1] ~^ image[0][12] + kernel[0][2] ~^ image[0][13] + kernel[0][3] ~^ image[0][14] + kernel[0][4] ~^ image[0][15] + kernel[1][0] ~^ image[1][11] + kernel[1][1] ~^ image[1][12] + kernel[1][2] ~^ image[1][13] + kernel[1][3] ~^ image[1][14] + kernel[1][4] ~^ image[1][15] + kernel[2][0] ~^ image[2][11] + kernel[2][1] ~^ image[2][12] + kernel[2][2] ~^ image[2][13] + kernel[2][3] ~^ image[2][14] + kernel[2][4] ~^ image[2][15] + kernel[3][0] ~^ image[3][11] + kernel[3][1] ~^ image[3][12] + kernel[3][2] ~^ image[3][13] + kernel[3][3] ~^ image[3][14] + kernel[3][4] ~^ image[3][15] + kernel[4][0] ~^ image[4][11] + kernel[4][1] ~^ image[4][12] + kernel[4][2] ~^ image[4][13] + kernel[4][3] ~^ image[4][14] + kernel[4][4] ~^ image[4][15];
assign xor_sum[0][12] = kernel[0][0] ~^ image[0][12] + kernel[0][1] ~^ image[0][13] + kernel[0][2] ~^ image[0][14] + kernel[0][3] ~^ image[0][15] + kernel[0][4] ~^ image[0][16] + kernel[1][0] ~^ image[1][12] + kernel[1][1] ~^ image[1][13] + kernel[1][2] ~^ image[1][14] + kernel[1][3] ~^ image[1][15] + kernel[1][4] ~^ image[1][16] + kernel[2][0] ~^ image[2][12] + kernel[2][1] ~^ image[2][13] + kernel[2][2] ~^ image[2][14] + kernel[2][3] ~^ image[2][15] + kernel[2][4] ~^ image[2][16] + kernel[3][0] ~^ image[3][12] + kernel[3][1] ~^ image[3][13] + kernel[3][2] ~^ image[3][14] + kernel[3][3] ~^ image[3][15] + kernel[3][4] ~^ image[3][16] + kernel[4][0] ~^ image[4][12] + kernel[4][1] ~^ image[4][13] + kernel[4][2] ~^ image[4][14] + kernel[4][3] ~^ image[4][15] + kernel[4][4] ~^ image[4][16];
assign xor_sum[0][13] = kernel[0][0] ~^ image[0][13] + kernel[0][1] ~^ image[0][14] + kernel[0][2] ~^ image[0][15] + kernel[0][3] ~^ image[0][16] + kernel[0][4] ~^ image[0][17] + kernel[1][0] ~^ image[1][13] + kernel[1][1] ~^ image[1][14] + kernel[1][2] ~^ image[1][15] + kernel[1][3] ~^ image[1][16] + kernel[1][4] ~^ image[1][17] + kernel[2][0] ~^ image[2][13] + kernel[2][1] ~^ image[2][14] + kernel[2][2] ~^ image[2][15] + kernel[2][3] ~^ image[2][16] + kernel[2][4] ~^ image[2][17] + kernel[3][0] ~^ image[3][13] + kernel[3][1] ~^ image[3][14] + kernel[3][2] ~^ image[3][15] + kernel[3][3] ~^ image[3][16] + kernel[3][4] ~^ image[3][17] + kernel[4][0] ~^ image[4][13] + kernel[4][1] ~^ image[4][14] + kernel[4][2] ~^ image[4][15] + kernel[4][3] ~^ image[4][16] + kernel[4][4] ~^ image[4][17];
assign xor_sum[0][14] = kernel[0][0] ~^ image[0][14] + kernel[0][1] ~^ image[0][15] + kernel[0][2] ~^ image[0][16] + kernel[0][3] ~^ image[0][17] + kernel[0][4] ~^ image[0][18] + kernel[1][0] ~^ image[1][14] + kernel[1][1] ~^ image[1][15] + kernel[1][2] ~^ image[1][16] + kernel[1][3] ~^ image[1][17] + kernel[1][4] ~^ image[1][18] + kernel[2][0] ~^ image[2][14] + kernel[2][1] ~^ image[2][15] + kernel[2][2] ~^ image[2][16] + kernel[2][3] ~^ image[2][17] + kernel[2][4] ~^ image[2][18] + kernel[3][0] ~^ image[3][14] + kernel[3][1] ~^ image[3][15] + kernel[3][2] ~^ image[3][16] + kernel[3][3] ~^ image[3][17] + kernel[3][4] ~^ image[3][18] + kernel[4][0] ~^ image[4][14] + kernel[4][1] ~^ image[4][15] + kernel[4][2] ~^ image[4][16] + kernel[4][3] ~^ image[4][17] + kernel[4][4] ~^ image[4][18];
assign xor_sum[0][15] = kernel[0][0] ~^ image[0][15] + kernel[0][1] ~^ image[0][16] + kernel[0][2] ~^ image[0][17] + kernel[0][3] ~^ image[0][18] + kernel[0][4] ~^ image[0][19] + kernel[1][0] ~^ image[1][15] + kernel[1][1] ~^ image[1][16] + kernel[1][2] ~^ image[1][17] + kernel[1][3] ~^ image[1][18] + kernel[1][4] ~^ image[1][19] + kernel[2][0] ~^ image[2][15] + kernel[2][1] ~^ image[2][16] + kernel[2][2] ~^ image[2][17] + kernel[2][3] ~^ image[2][18] + kernel[2][4] ~^ image[2][19] + kernel[3][0] ~^ image[3][15] + kernel[3][1] ~^ image[3][16] + kernel[3][2] ~^ image[3][17] + kernel[3][3] ~^ image[3][18] + kernel[3][4] ~^ image[3][19] + kernel[4][0] ~^ image[4][15] + kernel[4][1] ~^ image[4][16] + kernel[4][2] ~^ image[4][17] + kernel[4][3] ~^ image[4][18] + kernel[4][4] ~^ image[4][19];
assign xor_sum[0][16] = kernel[0][0] ~^ image[0][16] + kernel[0][1] ~^ image[0][17] + kernel[0][2] ~^ image[0][18] + kernel[0][3] ~^ image[0][19] + kernel[0][4] ~^ image[0][20] + kernel[1][0] ~^ image[1][16] + kernel[1][1] ~^ image[1][17] + kernel[1][2] ~^ image[1][18] + kernel[1][3] ~^ image[1][19] + kernel[1][4] ~^ image[1][20] + kernel[2][0] ~^ image[2][16] + kernel[2][1] ~^ image[2][17] + kernel[2][2] ~^ image[2][18] + kernel[2][3] ~^ image[2][19] + kernel[2][4] ~^ image[2][20] + kernel[3][0] ~^ image[3][16] + kernel[3][1] ~^ image[3][17] + kernel[3][2] ~^ image[3][18] + kernel[3][3] ~^ image[3][19] + kernel[3][4] ~^ image[3][20] + kernel[4][0] ~^ image[4][16] + kernel[4][1] ~^ image[4][17] + kernel[4][2] ~^ image[4][18] + kernel[4][3] ~^ image[4][19] + kernel[4][4] ~^ image[4][20];
assign xor_sum[0][17] = kernel[0][0] ~^ image[0][17] + kernel[0][1] ~^ image[0][18] + kernel[0][2] ~^ image[0][19] + kernel[0][3] ~^ image[0][20] + kernel[0][4] ~^ image[0][21] + kernel[1][0] ~^ image[1][17] + kernel[1][1] ~^ image[1][18] + kernel[1][2] ~^ image[1][19] + kernel[1][3] ~^ image[1][20] + kernel[1][4] ~^ image[1][21] + kernel[2][0] ~^ image[2][17] + kernel[2][1] ~^ image[2][18] + kernel[2][2] ~^ image[2][19] + kernel[2][3] ~^ image[2][20] + kernel[2][4] ~^ image[2][21] + kernel[3][0] ~^ image[3][17] + kernel[3][1] ~^ image[3][18] + kernel[3][2] ~^ image[3][19] + kernel[3][3] ~^ image[3][20] + kernel[3][4] ~^ image[3][21] + kernel[4][0] ~^ image[4][17] + kernel[4][1] ~^ image[4][18] + kernel[4][2] ~^ image[4][19] + kernel[4][3] ~^ image[4][20] + kernel[4][4] ~^ image[4][21];
assign xor_sum[0][18] = kernel[0][0] ~^ image[0][18] + kernel[0][1] ~^ image[0][19] + kernel[0][2] ~^ image[0][20] + kernel[0][3] ~^ image[0][21] + kernel[0][4] ~^ image[0][22] + kernel[1][0] ~^ image[1][18] + kernel[1][1] ~^ image[1][19] + kernel[1][2] ~^ image[1][20] + kernel[1][3] ~^ image[1][21] + kernel[1][4] ~^ image[1][22] + kernel[2][0] ~^ image[2][18] + kernel[2][1] ~^ image[2][19] + kernel[2][2] ~^ image[2][20] + kernel[2][3] ~^ image[2][21] + kernel[2][4] ~^ image[2][22] + kernel[3][0] ~^ image[3][18] + kernel[3][1] ~^ image[3][19] + kernel[3][2] ~^ image[3][20] + kernel[3][3] ~^ image[3][21] + kernel[3][4] ~^ image[3][22] + kernel[4][0] ~^ image[4][18] + kernel[4][1] ~^ image[4][19] + kernel[4][2] ~^ image[4][20] + kernel[4][3] ~^ image[4][21] + kernel[4][4] ~^ image[4][22];
assign xor_sum[0][19] = kernel[0][0] ~^ image[0][19] + kernel[0][1] ~^ image[0][20] + kernel[0][2] ~^ image[0][21] + kernel[0][3] ~^ image[0][22] + kernel[0][4] ~^ image[0][23] + kernel[1][0] ~^ image[1][19] + kernel[1][1] ~^ image[1][20] + kernel[1][2] ~^ image[1][21] + kernel[1][3] ~^ image[1][22] + kernel[1][4] ~^ image[1][23] + kernel[2][0] ~^ image[2][19] + kernel[2][1] ~^ image[2][20] + kernel[2][2] ~^ image[2][21] + kernel[2][3] ~^ image[2][22] + kernel[2][4] ~^ image[2][23] + kernel[3][0] ~^ image[3][19] + kernel[3][1] ~^ image[3][20] + kernel[3][2] ~^ image[3][21] + kernel[3][3] ~^ image[3][22] + kernel[3][4] ~^ image[3][23] + kernel[4][0] ~^ image[4][19] + kernel[4][1] ~^ image[4][20] + kernel[4][2] ~^ image[4][21] + kernel[4][3] ~^ image[4][22] + kernel[4][4] ~^ image[4][23];
assign xor_sum[0][20] = kernel[0][0] ~^ image[0][20] + kernel[0][1] ~^ image[0][21] + kernel[0][2] ~^ image[0][22] + kernel[0][3] ~^ image[0][23] + kernel[0][4] ~^ image[0][24] + kernel[1][0] ~^ image[1][20] + kernel[1][1] ~^ image[1][21] + kernel[1][2] ~^ image[1][22] + kernel[1][3] ~^ image[1][23] + kernel[1][4] ~^ image[1][24] + kernel[2][0] ~^ image[2][20] + kernel[2][1] ~^ image[2][21] + kernel[2][2] ~^ image[2][22] + kernel[2][3] ~^ image[2][23] + kernel[2][4] ~^ image[2][24] + kernel[3][0] ~^ image[3][20] + kernel[3][1] ~^ image[3][21] + kernel[3][2] ~^ image[3][22] + kernel[3][3] ~^ image[3][23] + kernel[3][4] ~^ image[3][24] + kernel[4][0] ~^ image[4][20] + kernel[4][1] ~^ image[4][21] + kernel[4][2] ~^ image[4][22] + kernel[4][3] ~^ image[4][23] + kernel[4][4] ~^ image[4][24];
assign xor_sum[0][21] = kernel[0][0] ~^ image[0][21] + kernel[0][1] ~^ image[0][22] + kernel[0][2] ~^ image[0][23] + kernel[0][3] ~^ image[0][24] + kernel[0][4] ~^ image[0][25] + kernel[1][0] ~^ image[1][21] + kernel[1][1] ~^ image[1][22] + kernel[1][2] ~^ image[1][23] + kernel[1][3] ~^ image[1][24] + kernel[1][4] ~^ image[1][25] + kernel[2][0] ~^ image[2][21] + kernel[2][1] ~^ image[2][22] + kernel[2][2] ~^ image[2][23] + kernel[2][3] ~^ image[2][24] + kernel[2][4] ~^ image[2][25] + kernel[3][0] ~^ image[3][21] + kernel[3][1] ~^ image[3][22] + kernel[3][2] ~^ image[3][23] + kernel[3][3] ~^ image[3][24] + kernel[3][4] ~^ image[3][25] + kernel[4][0] ~^ image[4][21] + kernel[4][1] ~^ image[4][22] + kernel[4][2] ~^ image[4][23] + kernel[4][3] ~^ image[4][24] + kernel[4][4] ~^ image[4][25];
assign xor_sum[0][22] = kernel[0][0] ~^ image[0][22] + kernel[0][1] ~^ image[0][23] + kernel[0][2] ~^ image[0][24] + kernel[0][3] ~^ image[0][25] + kernel[0][4] ~^ image[0][26] + kernel[1][0] ~^ image[1][22] + kernel[1][1] ~^ image[1][23] + kernel[1][2] ~^ image[1][24] + kernel[1][3] ~^ image[1][25] + kernel[1][4] ~^ image[1][26] + kernel[2][0] ~^ image[2][22] + kernel[2][1] ~^ image[2][23] + kernel[2][2] ~^ image[2][24] + kernel[2][3] ~^ image[2][25] + kernel[2][4] ~^ image[2][26] + kernel[3][0] ~^ image[3][22] + kernel[3][1] ~^ image[3][23] + kernel[3][2] ~^ image[3][24] + kernel[3][3] ~^ image[3][25] + kernel[3][4] ~^ image[3][26] + kernel[4][0] ~^ image[4][22] + kernel[4][1] ~^ image[4][23] + kernel[4][2] ~^ image[4][24] + kernel[4][3] ~^ image[4][25] + kernel[4][4] ~^ image[4][26];
assign xor_sum[0][23] = kernel[0][0] ~^ image[0][23] + kernel[0][1] ~^ image[0][24] + kernel[0][2] ~^ image[0][25] + kernel[0][3] ~^ image[0][26] + kernel[0][4] ~^ image[0][27] + kernel[1][0] ~^ image[1][23] + kernel[1][1] ~^ image[1][24] + kernel[1][2] ~^ image[1][25] + kernel[1][3] ~^ image[1][26] + kernel[1][4] ~^ image[1][27] + kernel[2][0] ~^ image[2][23] + kernel[2][1] ~^ image[2][24] + kernel[2][2] ~^ image[2][25] + kernel[2][3] ~^ image[2][26] + kernel[2][4] ~^ image[2][27] + kernel[3][0] ~^ image[3][23] + kernel[3][1] ~^ image[3][24] + kernel[3][2] ~^ image[3][25] + kernel[3][3] ~^ image[3][26] + kernel[3][4] ~^ image[3][27] + kernel[4][0] ~^ image[4][23] + kernel[4][1] ~^ image[4][24] + kernel[4][2] ~^ image[4][25] + kernel[4][3] ~^ image[4][26] + kernel[4][4] ~^ image[4][27];
assign xor_sum[1][0] = kernel[0][0] ~^ image[1][0] + kernel[0][1] ~^ image[1][1] + kernel[0][2] ~^ image[1][2] + kernel[0][3] ~^ image[1][3] + kernel[0][4] ~^ image[1][4] + kernel[1][0] ~^ image[2][0] + kernel[1][1] ~^ image[2][1] + kernel[1][2] ~^ image[2][2] + kernel[1][3] ~^ image[2][3] + kernel[1][4] ~^ image[2][4] + kernel[2][0] ~^ image[3][0] + kernel[2][1] ~^ image[3][1] + kernel[2][2] ~^ image[3][2] + kernel[2][3] ~^ image[3][3] + kernel[2][4] ~^ image[3][4] + kernel[3][0] ~^ image[4][0] + kernel[3][1] ~^ image[4][1] + kernel[3][2] ~^ image[4][2] + kernel[3][3] ~^ image[4][3] + kernel[3][4] ~^ image[4][4] + kernel[4][0] ~^ image[5][0] + kernel[4][1] ~^ image[5][1] + kernel[4][2] ~^ image[5][2] + kernel[4][3] ~^ image[5][3] + kernel[4][4] ~^ image[5][4];
assign xor_sum[1][1] = kernel[0][0] ~^ image[1][1] + kernel[0][1] ~^ image[1][2] + kernel[0][2] ~^ image[1][3] + kernel[0][3] ~^ image[1][4] + kernel[0][4] ~^ image[1][5] + kernel[1][0] ~^ image[2][1] + kernel[1][1] ~^ image[2][2] + kernel[1][2] ~^ image[2][3] + kernel[1][3] ~^ image[2][4] + kernel[1][4] ~^ image[2][5] + kernel[2][0] ~^ image[3][1] + kernel[2][1] ~^ image[3][2] + kernel[2][2] ~^ image[3][3] + kernel[2][3] ~^ image[3][4] + kernel[2][4] ~^ image[3][5] + kernel[3][0] ~^ image[4][1] + kernel[3][1] ~^ image[4][2] + kernel[3][2] ~^ image[4][3] + kernel[3][3] ~^ image[4][4] + kernel[3][4] ~^ image[4][5] + kernel[4][0] ~^ image[5][1] + kernel[4][1] ~^ image[5][2] + kernel[4][2] ~^ image[5][3] + kernel[4][3] ~^ image[5][4] + kernel[4][4] ~^ image[5][5];
assign xor_sum[1][2] = kernel[0][0] ~^ image[1][2] + kernel[0][1] ~^ image[1][3] + kernel[0][2] ~^ image[1][4] + kernel[0][3] ~^ image[1][5] + kernel[0][4] ~^ image[1][6] + kernel[1][0] ~^ image[2][2] + kernel[1][1] ~^ image[2][3] + kernel[1][2] ~^ image[2][4] + kernel[1][3] ~^ image[2][5] + kernel[1][4] ~^ image[2][6] + kernel[2][0] ~^ image[3][2] + kernel[2][1] ~^ image[3][3] + kernel[2][2] ~^ image[3][4] + kernel[2][3] ~^ image[3][5] + kernel[2][4] ~^ image[3][6] + kernel[3][0] ~^ image[4][2] + kernel[3][1] ~^ image[4][3] + kernel[3][2] ~^ image[4][4] + kernel[3][3] ~^ image[4][5] + kernel[3][4] ~^ image[4][6] + kernel[4][0] ~^ image[5][2] + kernel[4][1] ~^ image[5][3] + kernel[4][2] ~^ image[5][4] + kernel[4][3] ~^ image[5][5] + kernel[4][4] ~^ image[5][6];
assign xor_sum[1][3] = kernel[0][0] ~^ image[1][3] + kernel[0][1] ~^ image[1][4] + kernel[0][2] ~^ image[1][5] + kernel[0][3] ~^ image[1][6] + kernel[0][4] ~^ image[1][7] + kernel[1][0] ~^ image[2][3] + kernel[1][1] ~^ image[2][4] + kernel[1][2] ~^ image[2][5] + kernel[1][3] ~^ image[2][6] + kernel[1][4] ~^ image[2][7] + kernel[2][0] ~^ image[3][3] + kernel[2][1] ~^ image[3][4] + kernel[2][2] ~^ image[3][5] + kernel[2][3] ~^ image[3][6] + kernel[2][4] ~^ image[3][7] + kernel[3][0] ~^ image[4][3] + kernel[3][1] ~^ image[4][4] + kernel[3][2] ~^ image[4][5] + kernel[3][3] ~^ image[4][6] + kernel[3][4] ~^ image[4][7] + kernel[4][0] ~^ image[5][3] + kernel[4][1] ~^ image[5][4] + kernel[4][2] ~^ image[5][5] + kernel[4][3] ~^ image[5][6] + kernel[4][4] ~^ image[5][7];
assign xor_sum[1][4] = kernel[0][0] ~^ image[1][4] + kernel[0][1] ~^ image[1][5] + kernel[0][2] ~^ image[1][6] + kernel[0][3] ~^ image[1][7] + kernel[0][4] ~^ image[1][8] + kernel[1][0] ~^ image[2][4] + kernel[1][1] ~^ image[2][5] + kernel[1][2] ~^ image[2][6] + kernel[1][3] ~^ image[2][7] + kernel[1][4] ~^ image[2][8] + kernel[2][0] ~^ image[3][4] + kernel[2][1] ~^ image[3][5] + kernel[2][2] ~^ image[3][6] + kernel[2][3] ~^ image[3][7] + kernel[2][4] ~^ image[3][8] + kernel[3][0] ~^ image[4][4] + kernel[3][1] ~^ image[4][5] + kernel[3][2] ~^ image[4][6] + kernel[3][3] ~^ image[4][7] + kernel[3][4] ~^ image[4][8] + kernel[4][0] ~^ image[5][4] + kernel[4][1] ~^ image[5][5] + kernel[4][2] ~^ image[5][6] + kernel[4][3] ~^ image[5][7] + kernel[4][4] ~^ image[5][8];
assign xor_sum[1][5] = kernel[0][0] ~^ image[1][5] + kernel[0][1] ~^ image[1][6] + kernel[0][2] ~^ image[1][7] + kernel[0][3] ~^ image[1][8] + kernel[0][4] ~^ image[1][9] + kernel[1][0] ~^ image[2][5] + kernel[1][1] ~^ image[2][6] + kernel[1][2] ~^ image[2][7] + kernel[1][3] ~^ image[2][8] + kernel[1][4] ~^ image[2][9] + kernel[2][0] ~^ image[3][5] + kernel[2][1] ~^ image[3][6] + kernel[2][2] ~^ image[3][7] + kernel[2][3] ~^ image[3][8] + kernel[2][4] ~^ image[3][9] + kernel[3][0] ~^ image[4][5] + kernel[3][1] ~^ image[4][6] + kernel[3][2] ~^ image[4][7] + kernel[3][3] ~^ image[4][8] + kernel[3][4] ~^ image[4][9] + kernel[4][0] ~^ image[5][5] + kernel[4][1] ~^ image[5][6] + kernel[4][2] ~^ image[5][7] + kernel[4][3] ~^ image[5][8] + kernel[4][4] ~^ image[5][9];
assign xor_sum[1][6] = kernel[0][0] ~^ image[1][6] + kernel[0][1] ~^ image[1][7] + kernel[0][2] ~^ image[1][8] + kernel[0][3] ~^ image[1][9] + kernel[0][4] ~^ image[1][10] + kernel[1][0] ~^ image[2][6] + kernel[1][1] ~^ image[2][7] + kernel[1][2] ~^ image[2][8] + kernel[1][3] ~^ image[2][9] + kernel[1][4] ~^ image[2][10] + kernel[2][0] ~^ image[3][6] + kernel[2][1] ~^ image[3][7] + kernel[2][2] ~^ image[3][8] + kernel[2][3] ~^ image[3][9] + kernel[2][4] ~^ image[3][10] + kernel[3][0] ~^ image[4][6] + kernel[3][1] ~^ image[4][7] + kernel[3][2] ~^ image[4][8] + kernel[3][3] ~^ image[4][9] + kernel[3][4] ~^ image[4][10] + kernel[4][0] ~^ image[5][6] + kernel[4][1] ~^ image[5][7] + kernel[4][2] ~^ image[5][8] + kernel[4][3] ~^ image[5][9] + kernel[4][4] ~^ image[5][10];
assign xor_sum[1][7] = kernel[0][0] ~^ image[1][7] + kernel[0][1] ~^ image[1][8] + kernel[0][2] ~^ image[1][9] + kernel[0][3] ~^ image[1][10] + kernel[0][4] ~^ image[1][11] + kernel[1][0] ~^ image[2][7] + kernel[1][1] ~^ image[2][8] + kernel[1][2] ~^ image[2][9] + kernel[1][3] ~^ image[2][10] + kernel[1][4] ~^ image[2][11] + kernel[2][0] ~^ image[3][7] + kernel[2][1] ~^ image[3][8] + kernel[2][2] ~^ image[3][9] + kernel[2][3] ~^ image[3][10] + kernel[2][4] ~^ image[3][11] + kernel[3][0] ~^ image[4][7] + kernel[3][1] ~^ image[4][8] + kernel[3][2] ~^ image[4][9] + kernel[3][3] ~^ image[4][10] + kernel[3][4] ~^ image[4][11] + kernel[4][0] ~^ image[5][7] + kernel[4][1] ~^ image[5][8] + kernel[4][2] ~^ image[5][9] + kernel[4][3] ~^ image[5][10] + kernel[4][4] ~^ image[5][11];
assign xor_sum[1][8] = kernel[0][0] ~^ image[1][8] + kernel[0][1] ~^ image[1][9] + kernel[0][2] ~^ image[1][10] + kernel[0][3] ~^ image[1][11] + kernel[0][4] ~^ image[1][12] + kernel[1][0] ~^ image[2][8] + kernel[1][1] ~^ image[2][9] + kernel[1][2] ~^ image[2][10] + kernel[1][3] ~^ image[2][11] + kernel[1][4] ~^ image[2][12] + kernel[2][0] ~^ image[3][8] + kernel[2][1] ~^ image[3][9] + kernel[2][2] ~^ image[3][10] + kernel[2][3] ~^ image[3][11] + kernel[2][4] ~^ image[3][12] + kernel[3][0] ~^ image[4][8] + kernel[3][1] ~^ image[4][9] + kernel[3][2] ~^ image[4][10] + kernel[3][3] ~^ image[4][11] + kernel[3][4] ~^ image[4][12] + kernel[4][0] ~^ image[5][8] + kernel[4][1] ~^ image[5][9] + kernel[4][2] ~^ image[5][10] + kernel[4][3] ~^ image[5][11] + kernel[4][4] ~^ image[5][12];
assign xor_sum[1][9] = kernel[0][0] ~^ image[1][9] + kernel[0][1] ~^ image[1][10] + kernel[0][2] ~^ image[1][11] + kernel[0][3] ~^ image[1][12] + kernel[0][4] ~^ image[1][13] + kernel[1][0] ~^ image[2][9] + kernel[1][1] ~^ image[2][10] + kernel[1][2] ~^ image[2][11] + kernel[1][3] ~^ image[2][12] + kernel[1][4] ~^ image[2][13] + kernel[2][0] ~^ image[3][9] + kernel[2][1] ~^ image[3][10] + kernel[2][2] ~^ image[3][11] + kernel[2][3] ~^ image[3][12] + kernel[2][4] ~^ image[3][13] + kernel[3][0] ~^ image[4][9] + kernel[3][1] ~^ image[4][10] + kernel[3][2] ~^ image[4][11] + kernel[3][3] ~^ image[4][12] + kernel[3][4] ~^ image[4][13] + kernel[4][0] ~^ image[5][9] + kernel[4][1] ~^ image[5][10] + kernel[4][2] ~^ image[5][11] + kernel[4][3] ~^ image[5][12] + kernel[4][4] ~^ image[5][13];
assign xor_sum[1][10] = kernel[0][0] ~^ image[1][10] + kernel[0][1] ~^ image[1][11] + kernel[0][2] ~^ image[1][12] + kernel[0][3] ~^ image[1][13] + kernel[0][4] ~^ image[1][14] + kernel[1][0] ~^ image[2][10] + kernel[1][1] ~^ image[2][11] + kernel[1][2] ~^ image[2][12] + kernel[1][3] ~^ image[2][13] + kernel[1][4] ~^ image[2][14] + kernel[2][0] ~^ image[3][10] + kernel[2][1] ~^ image[3][11] + kernel[2][2] ~^ image[3][12] + kernel[2][3] ~^ image[3][13] + kernel[2][4] ~^ image[3][14] + kernel[3][0] ~^ image[4][10] + kernel[3][1] ~^ image[4][11] + kernel[3][2] ~^ image[4][12] + kernel[3][3] ~^ image[4][13] + kernel[3][4] ~^ image[4][14] + kernel[4][0] ~^ image[5][10] + kernel[4][1] ~^ image[5][11] + kernel[4][2] ~^ image[5][12] + kernel[4][3] ~^ image[5][13] + kernel[4][4] ~^ image[5][14];
assign xor_sum[1][11] = kernel[0][0] ~^ image[1][11] + kernel[0][1] ~^ image[1][12] + kernel[0][2] ~^ image[1][13] + kernel[0][3] ~^ image[1][14] + kernel[0][4] ~^ image[1][15] + kernel[1][0] ~^ image[2][11] + kernel[1][1] ~^ image[2][12] + kernel[1][2] ~^ image[2][13] + kernel[1][3] ~^ image[2][14] + kernel[1][4] ~^ image[2][15] + kernel[2][0] ~^ image[3][11] + kernel[2][1] ~^ image[3][12] + kernel[2][2] ~^ image[3][13] + kernel[2][3] ~^ image[3][14] + kernel[2][4] ~^ image[3][15] + kernel[3][0] ~^ image[4][11] + kernel[3][1] ~^ image[4][12] + kernel[3][2] ~^ image[4][13] + kernel[3][3] ~^ image[4][14] + kernel[3][4] ~^ image[4][15] + kernel[4][0] ~^ image[5][11] + kernel[4][1] ~^ image[5][12] + kernel[4][2] ~^ image[5][13] + kernel[4][3] ~^ image[5][14] + kernel[4][4] ~^ image[5][15];
assign xor_sum[1][12] = kernel[0][0] ~^ image[1][12] + kernel[0][1] ~^ image[1][13] + kernel[0][2] ~^ image[1][14] + kernel[0][3] ~^ image[1][15] + kernel[0][4] ~^ image[1][16] + kernel[1][0] ~^ image[2][12] + kernel[1][1] ~^ image[2][13] + kernel[1][2] ~^ image[2][14] + kernel[1][3] ~^ image[2][15] + kernel[1][4] ~^ image[2][16] + kernel[2][0] ~^ image[3][12] + kernel[2][1] ~^ image[3][13] + kernel[2][2] ~^ image[3][14] + kernel[2][3] ~^ image[3][15] + kernel[2][4] ~^ image[3][16] + kernel[3][0] ~^ image[4][12] + kernel[3][1] ~^ image[4][13] + kernel[3][2] ~^ image[4][14] + kernel[3][3] ~^ image[4][15] + kernel[3][4] ~^ image[4][16] + kernel[4][0] ~^ image[5][12] + kernel[4][1] ~^ image[5][13] + kernel[4][2] ~^ image[5][14] + kernel[4][3] ~^ image[5][15] + kernel[4][4] ~^ image[5][16];
assign xor_sum[1][13] = kernel[0][0] ~^ image[1][13] + kernel[0][1] ~^ image[1][14] + kernel[0][2] ~^ image[1][15] + kernel[0][3] ~^ image[1][16] + kernel[0][4] ~^ image[1][17] + kernel[1][0] ~^ image[2][13] + kernel[1][1] ~^ image[2][14] + kernel[1][2] ~^ image[2][15] + kernel[1][3] ~^ image[2][16] + kernel[1][4] ~^ image[2][17] + kernel[2][0] ~^ image[3][13] + kernel[2][1] ~^ image[3][14] + kernel[2][2] ~^ image[3][15] + kernel[2][3] ~^ image[3][16] + kernel[2][4] ~^ image[3][17] + kernel[3][0] ~^ image[4][13] + kernel[3][1] ~^ image[4][14] + kernel[3][2] ~^ image[4][15] + kernel[3][3] ~^ image[4][16] + kernel[3][4] ~^ image[4][17] + kernel[4][0] ~^ image[5][13] + kernel[4][1] ~^ image[5][14] + kernel[4][2] ~^ image[5][15] + kernel[4][3] ~^ image[5][16] + kernel[4][4] ~^ image[5][17];
assign xor_sum[1][14] = kernel[0][0] ~^ image[1][14] + kernel[0][1] ~^ image[1][15] + kernel[0][2] ~^ image[1][16] + kernel[0][3] ~^ image[1][17] + kernel[0][4] ~^ image[1][18] + kernel[1][0] ~^ image[2][14] + kernel[1][1] ~^ image[2][15] + kernel[1][2] ~^ image[2][16] + kernel[1][3] ~^ image[2][17] + kernel[1][4] ~^ image[2][18] + kernel[2][0] ~^ image[3][14] + kernel[2][1] ~^ image[3][15] + kernel[2][2] ~^ image[3][16] + kernel[2][3] ~^ image[3][17] + kernel[2][4] ~^ image[3][18] + kernel[3][0] ~^ image[4][14] + kernel[3][1] ~^ image[4][15] + kernel[3][2] ~^ image[4][16] + kernel[3][3] ~^ image[4][17] + kernel[3][4] ~^ image[4][18] + kernel[4][0] ~^ image[5][14] + kernel[4][1] ~^ image[5][15] + kernel[4][2] ~^ image[5][16] + kernel[4][3] ~^ image[5][17] + kernel[4][4] ~^ image[5][18];
assign xor_sum[1][15] = kernel[0][0] ~^ image[1][15] + kernel[0][1] ~^ image[1][16] + kernel[0][2] ~^ image[1][17] + kernel[0][3] ~^ image[1][18] + kernel[0][4] ~^ image[1][19] + kernel[1][0] ~^ image[2][15] + kernel[1][1] ~^ image[2][16] + kernel[1][2] ~^ image[2][17] + kernel[1][3] ~^ image[2][18] + kernel[1][4] ~^ image[2][19] + kernel[2][0] ~^ image[3][15] + kernel[2][1] ~^ image[3][16] + kernel[2][2] ~^ image[3][17] + kernel[2][3] ~^ image[3][18] + kernel[2][4] ~^ image[3][19] + kernel[3][0] ~^ image[4][15] + kernel[3][1] ~^ image[4][16] + kernel[3][2] ~^ image[4][17] + kernel[3][3] ~^ image[4][18] + kernel[3][4] ~^ image[4][19] + kernel[4][0] ~^ image[5][15] + kernel[4][1] ~^ image[5][16] + kernel[4][2] ~^ image[5][17] + kernel[4][3] ~^ image[5][18] + kernel[4][4] ~^ image[5][19];
assign xor_sum[1][16] = kernel[0][0] ~^ image[1][16] + kernel[0][1] ~^ image[1][17] + kernel[0][2] ~^ image[1][18] + kernel[0][3] ~^ image[1][19] + kernel[0][4] ~^ image[1][20] + kernel[1][0] ~^ image[2][16] + kernel[1][1] ~^ image[2][17] + kernel[1][2] ~^ image[2][18] + kernel[1][3] ~^ image[2][19] + kernel[1][4] ~^ image[2][20] + kernel[2][0] ~^ image[3][16] + kernel[2][1] ~^ image[3][17] + kernel[2][2] ~^ image[3][18] + kernel[2][3] ~^ image[3][19] + kernel[2][4] ~^ image[3][20] + kernel[3][0] ~^ image[4][16] + kernel[3][1] ~^ image[4][17] + kernel[3][2] ~^ image[4][18] + kernel[3][3] ~^ image[4][19] + kernel[3][4] ~^ image[4][20] + kernel[4][0] ~^ image[5][16] + kernel[4][1] ~^ image[5][17] + kernel[4][2] ~^ image[5][18] + kernel[4][3] ~^ image[5][19] + kernel[4][4] ~^ image[5][20];
assign xor_sum[1][17] = kernel[0][0] ~^ image[1][17] + kernel[0][1] ~^ image[1][18] + kernel[0][2] ~^ image[1][19] + kernel[0][3] ~^ image[1][20] + kernel[0][4] ~^ image[1][21] + kernel[1][0] ~^ image[2][17] + kernel[1][1] ~^ image[2][18] + kernel[1][2] ~^ image[2][19] + kernel[1][3] ~^ image[2][20] + kernel[1][4] ~^ image[2][21] + kernel[2][0] ~^ image[3][17] + kernel[2][1] ~^ image[3][18] + kernel[2][2] ~^ image[3][19] + kernel[2][3] ~^ image[3][20] + kernel[2][4] ~^ image[3][21] + kernel[3][0] ~^ image[4][17] + kernel[3][1] ~^ image[4][18] + kernel[3][2] ~^ image[4][19] + kernel[3][3] ~^ image[4][20] + kernel[3][4] ~^ image[4][21] + kernel[4][0] ~^ image[5][17] + kernel[4][1] ~^ image[5][18] + kernel[4][2] ~^ image[5][19] + kernel[4][3] ~^ image[5][20] + kernel[4][4] ~^ image[5][21];
assign xor_sum[1][18] = kernel[0][0] ~^ image[1][18] + kernel[0][1] ~^ image[1][19] + kernel[0][2] ~^ image[1][20] + kernel[0][3] ~^ image[1][21] + kernel[0][4] ~^ image[1][22] + kernel[1][0] ~^ image[2][18] + kernel[1][1] ~^ image[2][19] + kernel[1][2] ~^ image[2][20] + kernel[1][3] ~^ image[2][21] + kernel[1][4] ~^ image[2][22] + kernel[2][0] ~^ image[3][18] + kernel[2][1] ~^ image[3][19] + kernel[2][2] ~^ image[3][20] + kernel[2][3] ~^ image[3][21] + kernel[2][4] ~^ image[3][22] + kernel[3][0] ~^ image[4][18] + kernel[3][1] ~^ image[4][19] + kernel[3][2] ~^ image[4][20] + kernel[3][3] ~^ image[4][21] + kernel[3][4] ~^ image[4][22] + kernel[4][0] ~^ image[5][18] + kernel[4][1] ~^ image[5][19] + kernel[4][2] ~^ image[5][20] + kernel[4][3] ~^ image[5][21] + kernel[4][4] ~^ image[5][22];
assign xor_sum[1][19] = kernel[0][0] ~^ image[1][19] + kernel[0][1] ~^ image[1][20] + kernel[0][2] ~^ image[1][21] + kernel[0][3] ~^ image[1][22] + kernel[0][4] ~^ image[1][23] + kernel[1][0] ~^ image[2][19] + kernel[1][1] ~^ image[2][20] + kernel[1][2] ~^ image[2][21] + kernel[1][3] ~^ image[2][22] + kernel[1][4] ~^ image[2][23] + kernel[2][0] ~^ image[3][19] + kernel[2][1] ~^ image[3][20] + kernel[2][2] ~^ image[3][21] + kernel[2][3] ~^ image[3][22] + kernel[2][4] ~^ image[3][23] + kernel[3][0] ~^ image[4][19] + kernel[3][1] ~^ image[4][20] + kernel[3][2] ~^ image[4][21] + kernel[3][3] ~^ image[4][22] + kernel[3][4] ~^ image[4][23] + kernel[4][0] ~^ image[5][19] + kernel[4][1] ~^ image[5][20] + kernel[4][2] ~^ image[5][21] + kernel[4][3] ~^ image[5][22] + kernel[4][4] ~^ image[5][23];
assign xor_sum[1][20] = kernel[0][0] ~^ image[1][20] + kernel[0][1] ~^ image[1][21] + kernel[0][2] ~^ image[1][22] + kernel[0][3] ~^ image[1][23] + kernel[0][4] ~^ image[1][24] + kernel[1][0] ~^ image[2][20] + kernel[1][1] ~^ image[2][21] + kernel[1][2] ~^ image[2][22] + kernel[1][3] ~^ image[2][23] + kernel[1][4] ~^ image[2][24] + kernel[2][0] ~^ image[3][20] + kernel[2][1] ~^ image[3][21] + kernel[2][2] ~^ image[3][22] + kernel[2][3] ~^ image[3][23] + kernel[2][4] ~^ image[3][24] + kernel[3][0] ~^ image[4][20] + kernel[3][1] ~^ image[4][21] + kernel[3][2] ~^ image[4][22] + kernel[3][3] ~^ image[4][23] + kernel[3][4] ~^ image[4][24] + kernel[4][0] ~^ image[5][20] + kernel[4][1] ~^ image[5][21] + kernel[4][2] ~^ image[5][22] + kernel[4][3] ~^ image[5][23] + kernel[4][4] ~^ image[5][24];
assign xor_sum[1][21] = kernel[0][0] ~^ image[1][21] + kernel[0][1] ~^ image[1][22] + kernel[0][2] ~^ image[1][23] + kernel[0][3] ~^ image[1][24] + kernel[0][4] ~^ image[1][25] + kernel[1][0] ~^ image[2][21] + kernel[1][1] ~^ image[2][22] + kernel[1][2] ~^ image[2][23] + kernel[1][3] ~^ image[2][24] + kernel[1][4] ~^ image[2][25] + kernel[2][0] ~^ image[3][21] + kernel[2][1] ~^ image[3][22] + kernel[2][2] ~^ image[3][23] + kernel[2][3] ~^ image[3][24] + kernel[2][4] ~^ image[3][25] + kernel[3][0] ~^ image[4][21] + kernel[3][1] ~^ image[4][22] + kernel[3][2] ~^ image[4][23] + kernel[3][3] ~^ image[4][24] + kernel[3][4] ~^ image[4][25] + kernel[4][0] ~^ image[5][21] + kernel[4][1] ~^ image[5][22] + kernel[4][2] ~^ image[5][23] + kernel[4][3] ~^ image[5][24] + kernel[4][4] ~^ image[5][25];
assign xor_sum[1][22] = kernel[0][0] ~^ image[1][22] + kernel[0][1] ~^ image[1][23] + kernel[0][2] ~^ image[1][24] + kernel[0][3] ~^ image[1][25] + kernel[0][4] ~^ image[1][26] + kernel[1][0] ~^ image[2][22] + kernel[1][1] ~^ image[2][23] + kernel[1][2] ~^ image[2][24] + kernel[1][3] ~^ image[2][25] + kernel[1][4] ~^ image[2][26] + kernel[2][0] ~^ image[3][22] + kernel[2][1] ~^ image[3][23] + kernel[2][2] ~^ image[3][24] + kernel[2][3] ~^ image[3][25] + kernel[2][4] ~^ image[3][26] + kernel[3][0] ~^ image[4][22] + kernel[3][1] ~^ image[4][23] + kernel[3][2] ~^ image[4][24] + kernel[3][3] ~^ image[4][25] + kernel[3][4] ~^ image[4][26] + kernel[4][0] ~^ image[5][22] + kernel[4][1] ~^ image[5][23] + kernel[4][2] ~^ image[5][24] + kernel[4][3] ~^ image[5][25] + kernel[4][4] ~^ image[5][26];
assign xor_sum[1][23] = kernel[0][0] ~^ image[1][23] + kernel[0][1] ~^ image[1][24] + kernel[0][2] ~^ image[1][25] + kernel[0][3] ~^ image[1][26] + kernel[0][4] ~^ image[1][27] + kernel[1][0] ~^ image[2][23] + kernel[1][1] ~^ image[2][24] + kernel[1][2] ~^ image[2][25] + kernel[1][3] ~^ image[2][26] + kernel[1][4] ~^ image[2][27] + kernel[2][0] ~^ image[3][23] + kernel[2][1] ~^ image[3][24] + kernel[2][2] ~^ image[3][25] + kernel[2][3] ~^ image[3][26] + kernel[2][4] ~^ image[3][27] + kernel[3][0] ~^ image[4][23] + kernel[3][1] ~^ image[4][24] + kernel[3][2] ~^ image[4][25] + kernel[3][3] ~^ image[4][26] + kernel[3][4] ~^ image[4][27] + kernel[4][0] ~^ image[5][23] + kernel[4][1] ~^ image[5][24] + kernel[4][2] ~^ image[5][25] + kernel[4][3] ~^ image[5][26] + kernel[4][4] ~^ image[5][27];
assign xor_sum[2][0] = kernel[0][0] ~^ image[2][0] + kernel[0][1] ~^ image[2][1] + kernel[0][2] ~^ image[2][2] + kernel[0][3] ~^ image[2][3] + kernel[0][4] ~^ image[2][4] + kernel[1][0] ~^ image[3][0] + kernel[1][1] ~^ image[3][1] + kernel[1][2] ~^ image[3][2] + kernel[1][3] ~^ image[3][3] + kernel[1][4] ~^ image[3][4] + kernel[2][0] ~^ image[4][0] + kernel[2][1] ~^ image[4][1] + kernel[2][2] ~^ image[4][2] + kernel[2][3] ~^ image[4][3] + kernel[2][4] ~^ image[4][4] + kernel[3][0] ~^ image[5][0] + kernel[3][1] ~^ image[5][1] + kernel[3][2] ~^ image[5][2] + kernel[3][3] ~^ image[5][3] + kernel[3][4] ~^ image[5][4] + kernel[4][0] ~^ image[6][0] + kernel[4][1] ~^ image[6][1] + kernel[4][2] ~^ image[6][2] + kernel[4][3] ~^ image[6][3] + kernel[4][4] ~^ image[6][4];
assign xor_sum[2][1] = kernel[0][0] ~^ image[2][1] + kernel[0][1] ~^ image[2][2] + kernel[0][2] ~^ image[2][3] + kernel[0][3] ~^ image[2][4] + kernel[0][4] ~^ image[2][5] + kernel[1][0] ~^ image[3][1] + kernel[1][1] ~^ image[3][2] + kernel[1][2] ~^ image[3][3] + kernel[1][3] ~^ image[3][4] + kernel[1][4] ~^ image[3][5] + kernel[2][0] ~^ image[4][1] + kernel[2][1] ~^ image[4][2] + kernel[2][2] ~^ image[4][3] + kernel[2][3] ~^ image[4][4] + kernel[2][4] ~^ image[4][5] + kernel[3][0] ~^ image[5][1] + kernel[3][1] ~^ image[5][2] + kernel[3][2] ~^ image[5][3] + kernel[3][3] ~^ image[5][4] + kernel[3][4] ~^ image[5][5] + kernel[4][0] ~^ image[6][1] + kernel[4][1] ~^ image[6][2] + kernel[4][2] ~^ image[6][3] + kernel[4][3] ~^ image[6][4] + kernel[4][4] ~^ image[6][5];
assign xor_sum[2][2] = kernel[0][0] ~^ image[2][2] + kernel[0][1] ~^ image[2][3] + kernel[0][2] ~^ image[2][4] + kernel[0][3] ~^ image[2][5] + kernel[0][4] ~^ image[2][6] + kernel[1][0] ~^ image[3][2] + kernel[1][1] ~^ image[3][3] + kernel[1][2] ~^ image[3][4] + kernel[1][3] ~^ image[3][5] + kernel[1][4] ~^ image[3][6] + kernel[2][0] ~^ image[4][2] + kernel[2][1] ~^ image[4][3] + kernel[2][2] ~^ image[4][4] + kernel[2][3] ~^ image[4][5] + kernel[2][4] ~^ image[4][6] + kernel[3][0] ~^ image[5][2] + kernel[3][1] ~^ image[5][3] + kernel[3][2] ~^ image[5][4] + kernel[3][3] ~^ image[5][5] + kernel[3][4] ~^ image[5][6] + kernel[4][0] ~^ image[6][2] + kernel[4][1] ~^ image[6][3] + kernel[4][2] ~^ image[6][4] + kernel[4][3] ~^ image[6][5] + kernel[4][4] ~^ image[6][6];
assign xor_sum[2][3] = kernel[0][0] ~^ image[2][3] + kernel[0][1] ~^ image[2][4] + kernel[0][2] ~^ image[2][5] + kernel[0][3] ~^ image[2][6] + kernel[0][4] ~^ image[2][7] + kernel[1][0] ~^ image[3][3] + kernel[1][1] ~^ image[3][4] + kernel[1][2] ~^ image[3][5] + kernel[1][3] ~^ image[3][6] + kernel[1][4] ~^ image[3][7] + kernel[2][0] ~^ image[4][3] + kernel[2][1] ~^ image[4][4] + kernel[2][2] ~^ image[4][5] + kernel[2][3] ~^ image[4][6] + kernel[2][4] ~^ image[4][7] + kernel[3][0] ~^ image[5][3] + kernel[3][1] ~^ image[5][4] + kernel[3][2] ~^ image[5][5] + kernel[3][3] ~^ image[5][6] + kernel[3][4] ~^ image[5][7] + kernel[4][0] ~^ image[6][3] + kernel[4][1] ~^ image[6][4] + kernel[4][2] ~^ image[6][5] + kernel[4][3] ~^ image[6][6] + kernel[4][4] ~^ image[6][7];
assign xor_sum[2][4] = kernel[0][0] ~^ image[2][4] + kernel[0][1] ~^ image[2][5] + kernel[0][2] ~^ image[2][6] + kernel[0][3] ~^ image[2][7] + kernel[0][4] ~^ image[2][8] + kernel[1][0] ~^ image[3][4] + kernel[1][1] ~^ image[3][5] + kernel[1][2] ~^ image[3][6] + kernel[1][3] ~^ image[3][7] + kernel[1][4] ~^ image[3][8] + kernel[2][0] ~^ image[4][4] + kernel[2][1] ~^ image[4][5] + kernel[2][2] ~^ image[4][6] + kernel[2][3] ~^ image[4][7] + kernel[2][4] ~^ image[4][8] + kernel[3][0] ~^ image[5][4] + kernel[3][1] ~^ image[5][5] + kernel[3][2] ~^ image[5][6] + kernel[3][3] ~^ image[5][7] + kernel[3][4] ~^ image[5][8] + kernel[4][0] ~^ image[6][4] + kernel[4][1] ~^ image[6][5] + kernel[4][2] ~^ image[6][6] + kernel[4][3] ~^ image[6][7] + kernel[4][4] ~^ image[6][8];
assign xor_sum[2][5] = kernel[0][0] ~^ image[2][5] + kernel[0][1] ~^ image[2][6] + kernel[0][2] ~^ image[2][7] + kernel[0][3] ~^ image[2][8] + kernel[0][4] ~^ image[2][9] + kernel[1][0] ~^ image[3][5] + kernel[1][1] ~^ image[3][6] + kernel[1][2] ~^ image[3][7] + kernel[1][3] ~^ image[3][8] + kernel[1][4] ~^ image[3][9] + kernel[2][0] ~^ image[4][5] + kernel[2][1] ~^ image[4][6] + kernel[2][2] ~^ image[4][7] + kernel[2][3] ~^ image[4][8] + kernel[2][4] ~^ image[4][9] + kernel[3][0] ~^ image[5][5] + kernel[3][1] ~^ image[5][6] + kernel[3][2] ~^ image[5][7] + kernel[3][3] ~^ image[5][8] + kernel[3][4] ~^ image[5][9] + kernel[4][0] ~^ image[6][5] + kernel[4][1] ~^ image[6][6] + kernel[4][2] ~^ image[6][7] + kernel[4][3] ~^ image[6][8] + kernel[4][4] ~^ image[6][9];
assign xor_sum[2][6] = kernel[0][0] ~^ image[2][6] + kernel[0][1] ~^ image[2][7] + kernel[0][2] ~^ image[2][8] + kernel[0][3] ~^ image[2][9] + kernel[0][4] ~^ image[2][10] + kernel[1][0] ~^ image[3][6] + kernel[1][1] ~^ image[3][7] + kernel[1][2] ~^ image[3][8] + kernel[1][3] ~^ image[3][9] + kernel[1][4] ~^ image[3][10] + kernel[2][0] ~^ image[4][6] + kernel[2][1] ~^ image[4][7] + kernel[2][2] ~^ image[4][8] + kernel[2][3] ~^ image[4][9] + kernel[2][4] ~^ image[4][10] + kernel[3][0] ~^ image[5][6] + kernel[3][1] ~^ image[5][7] + kernel[3][2] ~^ image[5][8] + kernel[3][3] ~^ image[5][9] + kernel[3][4] ~^ image[5][10] + kernel[4][0] ~^ image[6][6] + kernel[4][1] ~^ image[6][7] + kernel[4][2] ~^ image[6][8] + kernel[4][3] ~^ image[6][9] + kernel[4][4] ~^ image[6][10];
assign xor_sum[2][7] = kernel[0][0] ~^ image[2][7] + kernel[0][1] ~^ image[2][8] + kernel[0][2] ~^ image[2][9] + kernel[0][3] ~^ image[2][10] + kernel[0][4] ~^ image[2][11] + kernel[1][0] ~^ image[3][7] + kernel[1][1] ~^ image[3][8] + kernel[1][2] ~^ image[3][9] + kernel[1][3] ~^ image[3][10] + kernel[1][4] ~^ image[3][11] + kernel[2][0] ~^ image[4][7] + kernel[2][1] ~^ image[4][8] + kernel[2][2] ~^ image[4][9] + kernel[2][3] ~^ image[4][10] + kernel[2][4] ~^ image[4][11] + kernel[3][0] ~^ image[5][7] + kernel[3][1] ~^ image[5][8] + kernel[3][2] ~^ image[5][9] + kernel[3][3] ~^ image[5][10] + kernel[3][4] ~^ image[5][11] + kernel[4][0] ~^ image[6][7] + kernel[4][1] ~^ image[6][8] + kernel[4][2] ~^ image[6][9] + kernel[4][3] ~^ image[6][10] + kernel[4][4] ~^ image[6][11];
assign xor_sum[2][8] = kernel[0][0] ~^ image[2][8] + kernel[0][1] ~^ image[2][9] + kernel[0][2] ~^ image[2][10] + kernel[0][3] ~^ image[2][11] + kernel[0][4] ~^ image[2][12] + kernel[1][0] ~^ image[3][8] + kernel[1][1] ~^ image[3][9] + kernel[1][2] ~^ image[3][10] + kernel[1][3] ~^ image[3][11] + kernel[1][4] ~^ image[3][12] + kernel[2][0] ~^ image[4][8] + kernel[2][1] ~^ image[4][9] + kernel[2][2] ~^ image[4][10] + kernel[2][3] ~^ image[4][11] + kernel[2][4] ~^ image[4][12] + kernel[3][0] ~^ image[5][8] + kernel[3][1] ~^ image[5][9] + kernel[3][2] ~^ image[5][10] + kernel[3][3] ~^ image[5][11] + kernel[3][4] ~^ image[5][12] + kernel[4][0] ~^ image[6][8] + kernel[4][1] ~^ image[6][9] + kernel[4][2] ~^ image[6][10] + kernel[4][3] ~^ image[6][11] + kernel[4][4] ~^ image[6][12];
assign xor_sum[2][9] = kernel[0][0] ~^ image[2][9] + kernel[0][1] ~^ image[2][10] + kernel[0][2] ~^ image[2][11] + kernel[0][3] ~^ image[2][12] + kernel[0][4] ~^ image[2][13] + kernel[1][0] ~^ image[3][9] + kernel[1][1] ~^ image[3][10] + kernel[1][2] ~^ image[3][11] + kernel[1][3] ~^ image[3][12] + kernel[1][4] ~^ image[3][13] + kernel[2][0] ~^ image[4][9] + kernel[2][1] ~^ image[4][10] + kernel[2][2] ~^ image[4][11] + kernel[2][3] ~^ image[4][12] + kernel[2][4] ~^ image[4][13] + kernel[3][0] ~^ image[5][9] + kernel[3][1] ~^ image[5][10] + kernel[3][2] ~^ image[5][11] + kernel[3][3] ~^ image[5][12] + kernel[3][4] ~^ image[5][13] + kernel[4][0] ~^ image[6][9] + kernel[4][1] ~^ image[6][10] + kernel[4][2] ~^ image[6][11] + kernel[4][3] ~^ image[6][12] + kernel[4][4] ~^ image[6][13];
assign xor_sum[2][10] = kernel[0][0] ~^ image[2][10] + kernel[0][1] ~^ image[2][11] + kernel[0][2] ~^ image[2][12] + kernel[0][3] ~^ image[2][13] + kernel[0][4] ~^ image[2][14] + kernel[1][0] ~^ image[3][10] + kernel[1][1] ~^ image[3][11] + kernel[1][2] ~^ image[3][12] + kernel[1][3] ~^ image[3][13] + kernel[1][4] ~^ image[3][14] + kernel[2][0] ~^ image[4][10] + kernel[2][1] ~^ image[4][11] + kernel[2][2] ~^ image[4][12] + kernel[2][3] ~^ image[4][13] + kernel[2][4] ~^ image[4][14] + kernel[3][0] ~^ image[5][10] + kernel[3][1] ~^ image[5][11] + kernel[3][2] ~^ image[5][12] + kernel[3][3] ~^ image[5][13] + kernel[3][4] ~^ image[5][14] + kernel[4][0] ~^ image[6][10] + kernel[4][1] ~^ image[6][11] + kernel[4][2] ~^ image[6][12] + kernel[4][3] ~^ image[6][13] + kernel[4][4] ~^ image[6][14];
assign xor_sum[2][11] = kernel[0][0] ~^ image[2][11] + kernel[0][1] ~^ image[2][12] + kernel[0][2] ~^ image[2][13] + kernel[0][3] ~^ image[2][14] + kernel[0][4] ~^ image[2][15] + kernel[1][0] ~^ image[3][11] + kernel[1][1] ~^ image[3][12] + kernel[1][2] ~^ image[3][13] + kernel[1][3] ~^ image[3][14] + kernel[1][4] ~^ image[3][15] + kernel[2][0] ~^ image[4][11] + kernel[2][1] ~^ image[4][12] + kernel[2][2] ~^ image[4][13] + kernel[2][3] ~^ image[4][14] + kernel[2][4] ~^ image[4][15] + kernel[3][0] ~^ image[5][11] + kernel[3][1] ~^ image[5][12] + kernel[3][2] ~^ image[5][13] + kernel[3][3] ~^ image[5][14] + kernel[3][4] ~^ image[5][15] + kernel[4][0] ~^ image[6][11] + kernel[4][1] ~^ image[6][12] + kernel[4][2] ~^ image[6][13] + kernel[4][3] ~^ image[6][14] + kernel[4][4] ~^ image[6][15];
assign xor_sum[2][12] = kernel[0][0] ~^ image[2][12] + kernel[0][1] ~^ image[2][13] + kernel[0][2] ~^ image[2][14] + kernel[0][3] ~^ image[2][15] + kernel[0][4] ~^ image[2][16] + kernel[1][0] ~^ image[3][12] + kernel[1][1] ~^ image[3][13] + kernel[1][2] ~^ image[3][14] + kernel[1][3] ~^ image[3][15] + kernel[1][4] ~^ image[3][16] + kernel[2][0] ~^ image[4][12] + kernel[2][1] ~^ image[4][13] + kernel[2][2] ~^ image[4][14] + kernel[2][3] ~^ image[4][15] + kernel[2][4] ~^ image[4][16] + kernel[3][0] ~^ image[5][12] + kernel[3][1] ~^ image[5][13] + kernel[3][2] ~^ image[5][14] + kernel[3][3] ~^ image[5][15] + kernel[3][4] ~^ image[5][16] + kernel[4][0] ~^ image[6][12] + kernel[4][1] ~^ image[6][13] + kernel[4][2] ~^ image[6][14] + kernel[4][3] ~^ image[6][15] + kernel[4][4] ~^ image[6][16];
assign xor_sum[2][13] = kernel[0][0] ~^ image[2][13] + kernel[0][1] ~^ image[2][14] + kernel[0][2] ~^ image[2][15] + kernel[0][3] ~^ image[2][16] + kernel[0][4] ~^ image[2][17] + kernel[1][0] ~^ image[3][13] + kernel[1][1] ~^ image[3][14] + kernel[1][2] ~^ image[3][15] + kernel[1][3] ~^ image[3][16] + kernel[1][4] ~^ image[3][17] + kernel[2][0] ~^ image[4][13] + kernel[2][1] ~^ image[4][14] + kernel[2][2] ~^ image[4][15] + kernel[2][3] ~^ image[4][16] + kernel[2][4] ~^ image[4][17] + kernel[3][0] ~^ image[5][13] + kernel[3][1] ~^ image[5][14] + kernel[3][2] ~^ image[5][15] + kernel[3][3] ~^ image[5][16] + kernel[3][4] ~^ image[5][17] + kernel[4][0] ~^ image[6][13] + kernel[4][1] ~^ image[6][14] + kernel[4][2] ~^ image[6][15] + kernel[4][3] ~^ image[6][16] + kernel[4][4] ~^ image[6][17];
assign xor_sum[2][14] = kernel[0][0] ~^ image[2][14] + kernel[0][1] ~^ image[2][15] + kernel[0][2] ~^ image[2][16] + kernel[0][3] ~^ image[2][17] + kernel[0][4] ~^ image[2][18] + kernel[1][0] ~^ image[3][14] + kernel[1][1] ~^ image[3][15] + kernel[1][2] ~^ image[3][16] + kernel[1][3] ~^ image[3][17] + kernel[1][4] ~^ image[3][18] + kernel[2][0] ~^ image[4][14] + kernel[2][1] ~^ image[4][15] + kernel[2][2] ~^ image[4][16] + kernel[2][3] ~^ image[4][17] + kernel[2][4] ~^ image[4][18] + kernel[3][0] ~^ image[5][14] + kernel[3][1] ~^ image[5][15] + kernel[3][2] ~^ image[5][16] + kernel[3][3] ~^ image[5][17] + kernel[3][4] ~^ image[5][18] + kernel[4][0] ~^ image[6][14] + kernel[4][1] ~^ image[6][15] + kernel[4][2] ~^ image[6][16] + kernel[4][3] ~^ image[6][17] + kernel[4][4] ~^ image[6][18];
assign xor_sum[2][15] = kernel[0][0] ~^ image[2][15] + kernel[0][1] ~^ image[2][16] + kernel[0][2] ~^ image[2][17] + kernel[0][3] ~^ image[2][18] + kernel[0][4] ~^ image[2][19] + kernel[1][0] ~^ image[3][15] + kernel[1][1] ~^ image[3][16] + kernel[1][2] ~^ image[3][17] + kernel[1][3] ~^ image[3][18] + kernel[1][4] ~^ image[3][19] + kernel[2][0] ~^ image[4][15] + kernel[2][1] ~^ image[4][16] + kernel[2][2] ~^ image[4][17] + kernel[2][3] ~^ image[4][18] + kernel[2][4] ~^ image[4][19] + kernel[3][0] ~^ image[5][15] + kernel[3][1] ~^ image[5][16] + kernel[3][2] ~^ image[5][17] + kernel[3][3] ~^ image[5][18] + kernel[3][4] ~^ image[5][19] + kernel[4][0] ~^ image[6][15] + kernel[4][1] ~^ image[6][16] + kernel[4][2] ~^ image[6][17] + kernel[4][3] ~^ image[6][18] + kernel[4][4] ~^ image[6][19];
assign xor_sum[2][16] = kernel[0][0] ~^ image[2][16] + kernel[0][1] ~^ image[2][17] + kernel[0][2] ~^ image[2][18] + kernel[0][3] ~^ image[2][19] + kernel[0][4] ~^ image[2][20] + kernel[1][0] ~^ image[3][16] + kernel[1][1] ~^ image[3][17] + kernel[1][2] ~^ image[3][18] + kernel[1][3] ~^ image[3][19] + kernel[1][4] ~^ image[3][20] + kernel[2][0] ~^ image[4][16] + kernel[2][1] ~^ image[4][17] + kernel[2][2] ~^ image[4][18] + kernel[2][3] ~^ image[4][19] + kernel[2][4] ~^ image[4][20] + kernel[3][0] ~^ image[5][16] + kernel[3][1] ~^ image[5][17] + kernel[3][2] ~^ image[5][18] + kernel[3][3] ~^ image[5][19] + kernel[3][4] ~^ image[5][20] + kernel[4][0] ~^ image[6][16] + kernel[4][1] ~^ image[6][17] + kernel[4][2] ~^ image[6][18] + kernel[4][3] ~^ image[6][19] + kernel[4][4] ~^ image[6][20];
assign xor_sum[2][17] = kernel[0][0] ~^ image[2][17] + kernel[0][1] ~^ image[2][18] + kernel[0][2] ~^ image[2][19] + kernel[0][3] ~^ image[2][20] + kernel[0][4] ~^ image[2][21] + kernel[1][0] ~^ image[3][17] + kernel[1][1] ~^ image[3][18] + kernel[1][2] ~^ image[3][19] + kernel[1][3] ~^ image[3][20] + kernel[1][4] ~^ image[3][21] + kernel[2][0] ~^ image[4][17] + kernel[2][1] ~^ image[4][18] + kernel[2][2] ~^ image[4][19] + kernel[2][3] ~^ image[4][20] + kernel[2][4] ~^ image[4][21] + kernel[3][0] ~^ image[5][17] + kernel[3][1] ~^ image[5][18] + kernel[3][2] ~^ image[5][19] + kernel[3][3] ~^ image[5][20] + kernel[3][4] ~^ image[5][21] + kernel[4][0] ~^ image[6][17] + kernel[4][1] ~^ image[6][18] + kernel[4][2] ~^ image[6][19] + kernel[4][3] ~^ image[6][20] + kernel[4][4] ~^ image[6][21];
assign xor_sum[2][18] = kernel[0][0] ~^ image[2][18] + kernel[0][1] ~^ image[2][19] + kernel[0][2] ~^ image[2][20] + kernel[0][3] ~^ image[2][21] + kernel[0][4] ~^ image[2][22] + kernel[1][0] ~^ image[3][18] + kernel[1][1] ~^ image[3][19] + kernel[1][2] ~^ image[3][20] + kernel[1][3] ~^ image[3][21] + kernel[1][4] ~^ image[3][22] + kernel[2][0] ~^ image[4][18] + kernel[2][1] ~^ image[4][19] + kernel[2][2] ~^ image[4][20] + kernel[2][3] ~^ image[4][21] + kernel[2][4] ~^ image[4][22] + kernel[3][0] ~^ image[5][18] + kernel[3][1] ~^ image[5][19] + kernel[3][2] ~^ image[5][20] + kernel[3][3] ~^ image[5][21] + kernel[3][4] ~^ image[5][22] + kernel[4][0] ~^ image[6][18] + kernel[4][1] ~^ image[6][19] + kernel[4][2] ~^ image[6][20] + kernel[4][3] ~^ image[6][21] + kernel[4][4] ~^ image[6][22];
assign xor_sum[2][19] = kernel[0][0] ~^ image[2][19] + kernel[0][1] ~^ image[2][20] + kernel[0][2] ~^ image[2][21] + kernel[0][3] ~^ image[2][22] + kernel[0][4] ~^ image[2][23] + kernel[1][0] ~^ image[3][19] + kernel[1][1] ~^ image[3][20] + kernel[1][2] ~^ image[3][21] + kernel[1][3] ~^ image[3][22] + kernel[1][4] ~^ image[3][23] + kernel[2][0] ~^ image[4][19] + kernel[2][1] ~^ image[4][20] + kernel[2][2] ~^ image[4][21] + kernel[2][3] ~^ image[4][22] + kernel[2][4] ~^ image[4][23] + kernel[3][0] ~^ image[5][19] + kernel[3][1] ~^ image[5][20] + kernel[3][2] ~^ image[5][21] + kernel[3][3] ~^ image[5][22] + kernel[3][4] ~^ image[5][23] + kernel[4][0] ~^ image[6][19] + kernel[4][1] ~^ image[6][20] + kernel[4][2] ~^ image[6][21] + kernel[4][3] ~^ image[6][22] + kernel[4][4] ~^ image[6][23];
assign xor_sum[2][20] = kernel[0][0] ~^ image[2][20] + kernel[0][1] ~^ image[2][21] + kernel[0][2] ~^ image[2][22] + kernel[0][3] ~^ image[2][23] + kernel[0][4] ~^ image[2][24] + kernel[1][0] ~^ image[3][20] + kernel[1][1] ~^ image[3][21] + kernel[1][2] ~^ image[3][22] + kernel[1][3] ~^ image[3][23] + kernel[1][4] ~^ image[3][24] + kernel[2][0] ~^ image[4][20] + kernel[2][1] ~^ image[4][21] + kernel[2][2] ~^ image[4][22] + kernel[2][3] ~^ image[4][23] + kernel[2][4] ~^ image[4][24] + kernel[3][0] ~^ image[5][20] + kernel[3][1] ~^ image[5][21] + kernel[3][2] ~^ image[5][22] + kernel[3][3] ~^ image[5][23] + kernel[3][4] ~^ image[5][24] + kernel[4][0] ~^ image[6][20] + kernel[4][1] ~^ image[6][21] + kernel[4][2] ~^ image[6][22] + kernel[4][3] ~^ image[6][23] + kernel[4][4] ~^ image[6][24];
assign xor_sum[2][21] = kernel[0][0] ~^ image[2][21] + kernel[0][1] ~^ image[2][22] + kernel[0][2] ~^ image[2][23] + kernel[0][3] ~^ image[2][24] + kernel[0][4] ~^ image[2][25] + kernel[1][0] ~^ image[3][21] + kernel[1][1] ~^ image[3][22] + kernel[1][2] ~^ image[3][23] + kernel[1][3] ~^ image[3][24] + kernel[1][4] ~^ image[3][25] + kernel[2][0] ~^ image[4][21] + kernel[2][1] ~^ image[4][22] + kernel[2][2] ~^ image[4][23] + kernel[2][3] ~^ image[4][24] + kernel[2][4] ~^ image[4][25] + kernel[3][0] ~^ image[5][21] + kernel[3][1] ~^ image[5][22] + kernel[3][2] ~^ image[5][23] + kernel[3][3] ~^ image[5][24] + kernel[3][4] ~^ image[5][25] + kernel[4][0] ~^ image[6][21] + kernel[4][1] ~^ image[6][22] + kernel[4][2] ~^ image[6][23] + kernel[4][3] ~^ image[6][24] + kernel[4][4] ~^ image[6][25];
assign xor_sum[2][22] = kernel[0][0] ~^ image[2][22] + kernel[0][1] ~^ image[2][23] + kernel[0][2] ~^ image[2][24] + kernel[0][3] ~^ image[2][25] + kernel[0][4] ~^ image[2][26] + kernel[1][0] ~^ image[3][22] + kernel[1][1] ~^ image[3][23] + kernel[1][2] ~^ image[3][24] + kernel[1][3] ~^ image[3][25] + kernel[1][4] ~^ image[3][26] + kernel[2][0] ~^ image[4][22] + kernel[2][1] ~^ image[4][23] + kernel[2][2] ~^ image[4][24] + kernel[2][3] ~^ image[4][25] + kernel[2][4] ~^ image[4][26] + kernel[3][0] ~^ image[5][22] + kernel[3][1] ~^ image[5][23] + kernel[3][2] ~^ image[5][24] + kernel[3][3] ~^ image[5][25] + kernel[3][4] ~^ image[5][26] + kernel[4][0] ~^ image[6][22] + kernel[4][1] ~^ image[6][23] + kernel[4][2] ~^ image[6][24] + kernel[4][3] ~^ image[6][25] + kernel[4][4] ~^ image[6][26];
assign xor_sum[2][23] = kernel[0][0] ~^ image[2][23] + kernel[0][1] ~^ image[2][24] + kernel[0][2] ~^ image[2][25] + kernel[0][3] ~^ image[2][26] + kernel[0][4] ~^ image[2][27] + kernel[1][0] ~^ image[3][23] + kernel[1][1] ~^ image[3][24] + kernel[1][2] ~^ image[3][25] + kernel[1][3] ~^ image[3][26] + kernel[1][4] ~^ image[3][27] + kernel[2][0] ~^ image[4][23] + kernel[2][1] ~^ image[4][24] + kernel[2][2] ~^ image[4][25] + kernel[2][3] ~^ image[4][26] + kernel[2][4] ~^ image[4][27] + kernel[3][0] ~^ image[5][23] + kernel[3][1] ~^ image[5][24] + kernel[3][2] ~^ image[5][25] + kernel[3][3] ~^ image[5][26] + kernel[3][4] ~^ image[5][27] + kernel[4][0] ~^ image[6][23] + kernel[4][1] ~^ image[6][24] + kernel[4][2] ~^ image[6][25] + kernel[4][3] ~^ image[6][26] + kernel[4][4] ~^ image[6][27];
assign xor_sum[3][0] = kernel[0][0] ~^ image[3][0] + kernel[0][1] ~^ image[3][1] + kernel[0][2] ~^ image[3][2] + kernel[0][3] ~^ image[3][3] + kernel[0][4] ~^ image[3][4] + kernel[1][0] ~^ image[4][0] + kernel[1][1] ~^ image[4][1] + kernel[1][2] ~^ image[4][2] + kernel[1][3] ~^ image[4][3] + kernel[1][4] ~^ image[4][4] + kernel[2][0] ~^ image[5][0] + kernel[2][1] ~^ image[5][1] + kernel[2][2] ~^ image[5][2] + kernel[2][3] ~^ image[5][3] + kernel[2][4] ~^ image[5][4] + kernel[3][0] ~^ image[6][0] + kernel[3][1] ~^ image[6][1] + kernel[3][2] ~^ image[6][2] + kernel[3][3] ~^ image[6][3] + kernel[3][4] ~^ image[6][4] + kernel[4][0] ~^ image[7][0] + kernel[4][1] ~^ image[7][1] + kernel[4][2] ~^ image[7][2] + kernel[4][3] ~^ image[7][3] + kernel[4][4] ~^ image[7][4];
assign xor_sum[3][1] = kernel[0][0] ~^ image[3][1] + kernel[0][1] ~^ image[3][2] + kernel[0][2] ~^ image[3][3] + kernel[0][3] ~^ image[3][4] + kernel[0][4] ~^ image[3][5] + kernel[1][0] ~^ image[4][1] + kernel[1][1] ~^ image[4][2] + kernel[1][2] ~^ image[4][3] + kernel[1][3] ~^ image[4][4] + kernel[1][4] ~^ image[4][5] + kernel[2][0] ~^ image[5][1] + kernel[2][1] ~^ image[5][2] + kernel[2][2] ~^ image[5][3] + kernel[2][3] ~^ image[5][4] + kernel[2][4] ~^ image[5][5] + kernel[3][0] ~^ image[6][1] + kernel[3][1] ~^ image[6][2] + kernel[3][2] ~^ image[6][3] + kernel[3][3] ~^ image[6][4] + kernel[3][4] ~^ image[6][5] + kernel[4][0] ~^ image[7][1] + kernel[4][1] ~^ image[7][2] + kernel[4][2] ~^ image[7][3] + kernel[4][3] ~^ image[7][4] + kernel[4][4] ~^ image[7][5];
assign xor_sum[3][2] = kernel[0][0] ~^ image[3][2] + kernel[0][1] ~^ image[3][3] + kernel[0][2] ~^ image[3][4] + kernel[0][3] ~^ image[3][5] + kernel[0][4] ~^ image[3][6] + kernel[1][0] ~^ image[4][2] + kernel[1][1] ~^ image[4][3] + kernel[1][2] ~^ image[4][4] + kernel[1][3] ~^ image[4][5] + kernel[1][4] ~^ image[4][6] + kernel[2][0] ~^ image[5][2] + kernel[2][1] ~^ image[5][3] + kernel[2][2] ~^ image[5][4] + kernel[2][3] ~^ image[5][5] + kernel[2][4] ~^ image[5][6] + kernel[3][0] ~^ image[6][2] + kernel[3][1] ~^ image[6][3] + kernel[3][2] ~^ image[6][4] + kernel[3][3] ~^ image[6][5] + kernel[3][4] ~^ image[6][6] + kernel[4][0] ~^ image[7][2] + kernel[4][1] ~^ image[7][3] + kernel[4][2] ~^ image[7][4] + kernel[4][3] ~^ image[7][5] + kernel[4][4] ~^ image[7][6];
assign xor_sum[3][3] = kernel[0][0] ~^ image[3][3] + kernel[0][1] ~^ image[3][4] + kernel[0][2] ~^ image[3][5] + kernel[0][3] ~^ image[3][6] + kernel[0][4] ~^ image[3][7] + kernel[1][0] ~^ image[4][3] + kernel[1][1] ~^ image[4][4] + kernel[1][2] ~^ image[4][5] + kernel[1][3] ~^ image[4][6] + kernel[1][4] ~^ image[4][7] + kernel[2][0] ~^ image[5][3] + kernel[2][1] ~^ image[5][4] + kernel[2][2] ~^ image[5][5] + kernel[2][3] ~^ image[5][6] + kernel[2][4] ~^ image[5][7] + kernel[3][0] ~^ image[6][3] + kernel[3][1] ~^ image[6][4] + kernel[3][2] ~^ image[6][5] + kernel[3][3] ~^ image[6][6] + kernel[3][4] ~^ image[6][7] + kernel[4][0] ~^ image[7][3] + kernel[4][1] ~^ image[7][4] + kernel[4][2] ~^ image[7][5] + kernel[4][3] ~^ image[7][6] + kernel[4][4] ~^ image[7][7];
assign xor_sum[3][4] = kernel[0][0] ~^ image[3][4] + kernel[0][1] ~^ image[3][5] + kernel[0][2] ~^ image[3][6] + kernel[0][3] ~^ image[3][7] + kernel[0][4] ~^ image[3][8] + kernel[1][0] ~^ image[4][4] + kernel[1][1] ~^ image[4][5] + kernel[1][2] ~^ image[4][6] + kernel[1][3] ~^ image[4][7] + kernel[1][4] ~^ image[4][8] + kernel[2][0] ~^ image[5][4] + kernel[2][1] ~^ image[5][5] + kernel[2][2] ~^ image[5][6] + kernel[2][3] ~^ image[5][7] + kernel[2][4] ~^ image[5][8] + kernel[3][0] ~^ image[6][4] + kernel[3][1] ~^ image[6][5] + kernel[3][2] ~^ image[6][6] + kernel[3][3] ~^ image[6][7] + kernel[3][4] ~^ image[6][8] + kernel[4][0] ~^ image[7][4] + kernel[4][1] ~^ image[7][5] + kernel[4][2] ~^ image[7][6] + kernel[4][3] ~^ image[7][7] + kernel[4][4] ~^ image[7][8];
assign xor_sum[3][5] = kernel[0][0] ~^ image[3][5] + kernel[0][1] ~^ image[3][6] + kernel[0][2] ~^ image[3][7] + kernel[0][3] ~^ image[3][8] + kernel[0][4] ~^ image[3][9] + kernel[1][0] ~^ image[4][5] + kernel[1][1] ~^ image[4][6] + kernel[1][2] ~^ image[4][7] + kernel[1][3] ~^ image[4][8] + kernel[1][4] ~^ image[4][9] + kernel[2][0] ~^ image[5][5] + kernel[2][1] ~^ image[5][6] + kernel[2][2] ~^ image[5][7] + kernel[2][3] ~^ image[5][8] + kernel[2][4] ~^ image[5][9] + kernel[3][0] ~^ image[6][5] + kernel[3][1] ~^ image[6][6] + kernel[3][2] ~^ image[6][7] + kernel[3][3] ~^ image[6][8] + kernel[3][4] ~^ image[6][9] + kernel[4][0] ~^ image[7][5] + kernel[4][1] ~^ image[7][6] + kernel[4][2] ~^ image[7][7] + kernel[4][3] ~^ image[7][8] + kernel[4][4] ~^ image[7][9];
assign xor_sum[3][6] = kernel[0][0] ~^ image[3][6] + kernel[0][1] ~^ image[3][7] + kernel[0][2] ~^ image[3][8] + kernel[0][3] ~^ image[3][9] + kernel[0][4] ~^ image[3][10] + kernel[1][0] ~^ image[4][6] + kernel[1][1] ~^ image[4][7] + kernel[1][2] ~^ image[4][8] + kernel[1][3] ~^ image[4][9] + kernel[1][4] ~^ image[4][10] + kernel[2][0] ~^ image[5][6] + kernel[2][1] ~^ image[5][7] + kernel[2][2] ~^ image[5][8] + kernel[2][3] ~^ image[5][9] + kernel[2][4] ~^ image[5][10] + kernel[3][0] ~^ image[6][6] + kernel[3][1] ~^ image[6][7] + kernel[3][2] ~^ image[6][8] + kernel[3][3] ~^ image[6][9] + kernel[3][4] ~^ image[6][10] + kernel[4][0] ~^ image[7][6] + kernel[4][1] ~^ image[7][7] + kernel[4][2] ~^ image[7][8] + kernel[4][3] ~^ image[7][9] + kernel[4][4] ~^ image[7][10];
assign xor_sum[3][7] = kernel[0][0] ~^ image[3][7] + kernel[0][1] ~^ image[3][8] + kernel[0][2] ~^ image[3][9] + kernel[0][3] ~^ image[3][10] + kernel[0][4] ~^ image[3][11] + kernel[1][0] ~^ image[4][7] + kernel[1][1] ~^ image[4][8] + kernel[1][2] ~^ image[4][9] + kernel[1][3] ~^ image[4][10] + kernel[1][4] ~^ image[4][11] + kernel[2][0] ~^ image[5][7] + kernel[2][1] ~^ image[5][8] + kernel[2][2] ~^ image[5][9] + kernel[2][3] ~^ image[5][10] + kernel[2][4] ~^ image[5][11] + kernel[3][0] ~^ image[6][7] + kernel[3][1] ~^ image[6][8] + kernel[3][2] ~^ image[6][9] + kernel[3][3] ~^ image[6][10] + kernel[3][4] ~^ image[6][11] + kernel[4][0] ~^ image[7][7] + kernel[4][1] ~^ image[7][8] + kernel[4][2] ~^ image[7][9] + kernel[4][3] ~^ image[7][10] + kernel[4][4] ~^ image[7][11];
assign xor_sum[3][8] = kernel[0][0] ~^ image[3][8] + kernel[0][1] ~^ image[3][9] + kernel[0][2] ~^ image[3][10] + kernel[0][3] ~^ image[3][11] + kernel[0][4] ~^ image[3][12] + kernel[1][0] ~^ image[4][8] + kernel[1][1] ~^ image[4][9] + kernel[1][2] ~^ image[4][10] + kernel[1][3] ~^ image[4][11] + kernel[1][4] ~^ image[4][12] + kernel[2][0] ~^ image[5][8] + kernel[2][1] ~^ image[5][9] + kernel[2][2] ~^ image[5][10] + kernel[2][3] ~^ image[5][11] + kernel[2][4] ~^ image[5][12] + kernel[3][0] ~^ image[6][8] + kernel[3][1] ~^ image[6][9] + kernel[3][2] ~^ image[6][10] + kernel[3][3] ~^ image[6][11] + kernel[3][4] ~^ image[6][12] + kernel[4][0] ~^ image[7][8] + kernel[4][1] ~^ image[7][9] + kernel[4][2] ~^ image[7][10] + kernel[4][3] ~^ image[7][11] + kernel[4][4] ~^ image[7][12];
assign xor_sum[3][9] = kernel[0][0] ~^ image[3][9] + kernel[0][1] ~^ image[3][10] + kernel[0][2] ~^ image[3][11] + kernel[0][3] ~^ image[3][12] + kernel[0][4] ~^ image[3][13] + kernel[1][0] ~^ image[4][9] + kernel[1][1] ~^ image[4][10] + kernel[1][2] ~^ image[4][11] + kernel[1][3] ~^ image[4][12] + kernel[1][4] ~^ image[4][13] + kernel[2][0] ~^ image[5][9] + kernel[2][1] ~^ image[5][10] + kernel[2][2] ~^ image[5][11] + kernel[2][3] ~^ image[5][12] + kernel[2][4] ~^ image[5][13] + kernel[3][0] ~^ image[6][9] + kernel[3][1] ~^ image[6][10] + kernel[3][2] ~^ image[6][11] + kernel[3][3] ~^ image[6][12] + kernel[3][4] ~^ image[6][13] + kernel[4][0] ~^ image[7][9] + kernel[4][1] ~^ image[7][10] + kernel[4][2] ~^ image[7][11] + kernel[4][3] ~^ image[7][12] + kernel[4][4] ~^ image[7][13];
assign xor_sum[3][10] = kernel[0][0] ~^ image[3][10] + kernel[0][1] ~^ image[3][11] + kernel[0][2] ~^ image[3][12] + kernel[0][3] ~^ image[3][13] + kernel[0][4] ~^ image[3][14] + kernel[1][0] ~^ image[4][10] + kernel[1][1] ~^ image[4][11] + kernel[1][2] ~^ image[4][12] + kernel[1][3] ~^ image[4][13] + kernel[1][4] ~^ image[4][14] + kernel[2][0] ~^ image[5][10] + kernel[2][1] ~^ image[5][11] + kernel[2][2] ~^ image[5][12] + kernel[2][3] ~^ image[5][13] + kernel[2][4] ~^ image[5][14] + kernel[3][0] ~^ image[6][10] + kernel[3][1] ~^ image[6][11] + kernel[3][2] ~^ image[6][12] + kernel[3][3] ~^ image[6][13] + kernel[3][4] ~^ image[6][14] + kernel[4][0] ~^ image[7][10] + kernel[4][1] ~^ image[7][11] + kernel[4][2] ~^ image[7][12] + kernel[4][3] ~^ image[7][13] + kernel[4][4] ~^ image[7][14];
assign xor_sum[3][11] = kernel[0][0] ~^ image[3][11] + kernel[0][1] ~^ image[3][12] + kernel[0][2] ~^ image[3][13] + kernel[0][3] ~^ image[3][14] + kernel[0][4] ~^ image[3][15] + kernel[1][0] ~^ image[4][11] + kernel[1][1] ~^ image[4][12] + kernel[1][2] ~^ image[4][13] + kernel[1][3] ~^ image[4][14] + kernel[1][4] ~^ image[4][15] + kernel[2][0] ~^ image[5][11] + kernel[2][1] ~^ image[5][12] + kernel[2][2] ~^ image[5][13] + kernel[2][3] ~^ image[5][14] + kernel[2][4] ~^ image[5][15] + kernel[3][0] ~^ image[6][11] + kernel[3][1] ~^ image[6][12] + kernel[3][2] ~^ image[6][13] + kernel[3][3] ~^ image[6][14] + kernel[3][4] ~^ image[6][15] + kernel[4][0] ~^ image[7][11] + kernel[4][1] ~^ image[7][12] + kernel[4][2] ~^ image[7][13] + kernel[4][3] ~^ image[7][14] + kernel[4][4] ~^ image[7][15];
assign xor_sum[3][12] = kernel[0][0] ~^ image[3][12] + kernel[0][1] ~^ image[3][13] + kernel[0][2] ~^ image[3][14] + kernel[0][3] ~^ image[3][15] + kernel[0][4] ~^ image[3][16] + kernel[1][0] ~^ image[4][12] + kernel[1][1] ~^ image[4][13] + kernel[1][2] ~^ image[4][14] + kernel[1][3] ~^ image[4][15] + kernel[1][4] ~^ image[4][16] + kernel[2][0] ~^ image[5][12] + kernel[2][1] ~^ image[5][13] + kernel[2][2] ~^ image[5][14] + kernel[2][3] ~^ image[5][15] + kernel[2][4] ~^ image[5][16] + kernel[3][0] ~^ image[6][12] + kernel[3][1] ~^ image[6][13] + kernel[3][2] ~^ image[6][14] + kernel[3][3] ~^ image[6][15] + kernel[3][4] ~^ image[6][16] + kernel[4][0] ~^ image[7][12] + kernel[4][1] ~^ image[7][13] + kernel[4][2] ~^ image[7][14] + kernel[4][3] ~^ image[7][15] + kernel[4][4] ~^ image[7][16];
assign xor_sum[3][13] = kernel[0][0] ~^ image[3][13] + kernel[0][1] ~^ image[3][14] + kernel[0][2] ~^ image[3][15] + kernel[0][3] ~^ image[3][16] + kernel[0][4] ~^ image[3][17] + kernel[1][0] ~^ image[4][13] + kernel[1][1] ~^ image[4][14] + kernel[1][2] ~^ image[4][15] + kernel[1][3] ~^ image[4][16] + kernel[1][4] ~^ image[4][17] + kernel[2][0] ~^ image[5][13] + kernel[2][1] ~^ image[5][14] + kernel[2][2] ~^ image[5][15] + kernel[2][3] ~^ image[5][16] + kernel[2][4] ~^ image[5][17] + kernel[3][0] ~^ image[6][13] + kernel[3][1] ~^ image[6][14] + kernel[3][2] ~^ image[6][15] + kernel[3][3] ~^ image[6][16] + kernel[3][4] ~^ image[6][17] + kernel[4][0] ~^ image[7][13] + kernel[4][1] ~^ image[7][14] + kernel[4][2] ~^ image[7][15] + kernel[4][3] ~^ image[7][16] + kernel[4][4] ~^ image[7][17];
assign xor_sum[3][14] = kernel[0][0] ~^ image[3][14] + kernel[0][1] ~^ image[3][15] + kernel[0][2] ~^ image[3][16] + kernel[0][3] ~^ image[3][17] + kernel[0][4] ~^ image[3][18] + kernel[1][0] ~^ image[4][14] + kernel[1][1] ~^ image[4][15] + kernel[1][2] ~^ image[4][16] + kernel[1][3] ~^ image[4][17] + kernel[1][4] ~^ image[4][18] + kernel[2][0] ~^ image[5][14] + kernel[2][1] ~^ image[5][15] + kernel[2][2] ~^ image[5][16] + kernel[2][3] ~^ image[5][17] + kernel[2][4] ~^ image[5][18] + kernel[3][0] ~^ image[6][14] + kernel[3][1] ~^ image[6][15] + kernel[3][2] ~^ image[6][16] + kernel[3][3] ~^ image[6][17] + kernel[3][4] ~^ image[6][18] + kernel[4][0] ~^ image[7][14] + kernel[4][1] ~^ image[7][15] + kernel[4][2] ~^ image[7][16] + kernel[4][3] ~^ image[7][17] + kernel[4][4] ~^ image[7][18];
assign xor_sum[3][15] = kernel[0][0] ~^ image[3][15] + kernel[0][1] ~^ image[3][16] + kernel[0][2] ~^ image[3][17] + kernel[0][3] ~^ image[3][18] + kernel[0][4] ~^ image[3][19] + kernel[1][0] ~^ image[4][15] + kernel[1][1] ~^ image[4][16] + kernel[1][2] ~^ image[4][17] + kernel[1][3] ~^ image[4][18] + kernel[1][4] ~^ image[4][19] + kernel[2][0] ~^ image[5][15] + kernel[2][1] ~^ image[5][16] + kernel[2][2] ~^ image[5][17] + kernel[2][3] ~^ image[5][18] + kernel[2][4] ~^ image[5][19] + kernel[3][0] ~^ image[6][15] + kernel[3][1] ~^ image[6][16] + kernel[3][2] ~^ image[6][17] + kernel[3][3] ~^ image[6][18] + kernel[3][4] ~^ image[6][19] + kernel[4][0] ~^ image[7][15] + kernel[4][1] ~^ image[7][16] + kernel[4][2] ~^ image[7][17] + kernel[4][3] ~^ image[7][18] + kernel[4][4] ~^ image[7][19];
assign xor_sum[3][16] = kernel[0][0] ~^ image[3][16] + kernel[0][1] ~^ image[3][17] + kernel[0][2] ~^ image[3][18] + kernel[0][3] ~^ image[3][19] + kernel[0][4] ~^ image[3][20] + kernel[1][0] ~^ image[4][16] + kernel[1][1] ~^ image[4][17] + kernel[1][2] ~^ image[4][18] + kernel[1][3] ~^ image[4][19] + kernel[1][4] ~^ image[4][20] + kernel[2][0] ~^ image[5][16] + kernel[2][1] ~^ image[5][17] + kernel[2][2] ~^ image[5][18] + kernel[2][3] ~^ image[5][19] + kernel[2][4] ~^ image[5][20] + kernel[3][0] ~^ image[6][16] + kernel[3][1] ~^ image[6][17] + kernel[3][2] ~^ image[6][18] + kernel[3][3] ~^ image[6][19] + kernel[3][4] ~^ image[6][20] + kernel[4][0] ~^ image[7][16] + kernel[4][1] ~^ image[7][17] + kernel[4][2] ~^ image[7][18] + kernel[4][3] ~^ image[7][19] + kernel[4][4] ~^ image[7][20];
assign xor_sum[3][17] = kernel[0][0] ~^ image[3][17] + kernel[0][1] ~^ image[3][18] + kernel[0][2] ~^ image[3][19] + kernel[0][3] ~^ image[3][20] + kernel[0][4] ~^ image[3][21] + kernel[1][0] ~^ image[4][17] + kernel[1][1] ~^ image[4][18] + kernel[1][2] ~^ image[4][19] + kernel[1][3] ~^ image[4][20] + kernel[1][4] ~^ image[4][21] + kernel[2][0] ~^ image[5][17] + kernel[2][1] ~^ image[5][18] + kernel[2][2] ~^ image[5][19] + kernel[2][3] ~^ image[5][20] + kernel[2][4] ~^ image[5][21] + kernel[3][0] ~^ image[6][17] + kernel[3][1] ~^ image[6][18] + kernel[3][2] ~^ image[6][19] + kernel[3][3] ~^ image[6][20] + kernel[3][4] ~^ image[6][21] + kernel[4][0] ~^ image[7][17] + kernel[4][1] ~^ image[7][18] + kernel[4][2] ~^ image[7][19] + kernel[4][3] ~^ image[7][20] + kernel[4][4] ~^ image[7][21];
assign xor_sum[3][18] = kernel[0][0] ~^ image[3][18] + kernel[0][1] ~^ image[3][19] + kernel[0][2] ~^ image[3][20] + kernel[0][3] ~^ image[3][21] + kernel[0][4] ~^ image[3][22] + kernel[1][0] ~^ image[4][18] + kernel[1][1] ~^ image[4][19] + kernel[1][2] ~^ image[4][20] + kernel[1][3] ~^ image[4][21] + kernel[1][4] ~^ image[4][22] + kernel[2][0] ~^ image[5][18] + kernel[2][1] ~^ image[5][19] + kernel[2][2] ~^ image[5][20] + kernel[2][3] ~^ image[5][21] + kernel[2][4] ~^ image[5][22] + kernel[3][0] ~^ image[6][18] + kernel[3][1] ~^ image[6][19] + kernel[3][2] ~^ image[6][20] + kernel[3][3] ~^ image[6][21] + kernel[3][4] ~^ image[6][22] + kernel[4][0] ~^ image[7][18] + kernel[4][1] ~^ image[7][19] + kernel[4][2] ~^ image[7][20] + kernel[4][3] ~^ image[7][21] + kernel[4][4] ~^ image[7][22];
assign xor_sum[3][19] = kernel[0][0] ~^ image[3][19] + kernel[0][1] ~^ image[3][20] + kernel[0][2] ~^ image[3][21] + kernel[0][3] ~^ image[3][22] + kernel[0][4] ~^ image[3][23] + kernel[1][0] ~^ image[4][19] + kernel[1][1] ~^ image[4][20] + kernel[1][2] ~^ image[4][21] + kernel[1][3] ~^ image[4][22] + kernel[1][4] ~^ image[4][23] + kernel[2][0] ~^ image[5][19] + kernel[2][1] ~^ image[5][20] + kernel[2][2] ~^ image[5][21] + kernel[2][3] ~^ image[5][22] + kernel[2][4] ~^ image[5][23] + kernel[3][0] ~^ image[6][19] + kernel[3][1] ~^ image[6][20] + kernel[3][2] ~^ image[6][21] + kernel[3][3] ~^ image[6][22] + kernel[3][4] ~^ image[6][23] + kernel[4][0] ~^ image[7][19] + kernel[4][1] ~^ image[7][20] + kernel[4][2] ~^ image[7][21] + kernel[4][3] ~^ image[7][22] + kernel[4][4] ~^ image[7][23];
assign xor_sum[3][20] = kernel[0][0] ~^ image[3][20] + kernel[0][1] ~^ image[3][21] + kernel[0][2] ~^ image[3][22] + kernel[0][3] ~^ image[3][23] + kernel[0][4] ~^ image[3][24] + kernel[1][0] ~^ image[4][20] + kernel[1][1] ~^ image[4][21] + kernel[1][2] ~^ image[4][22] + kernel[1][3] ~^ image[4][23] + kernel[1][4] ~^ image[4][24] + kernel[2][0] ~^ image[5][20] + kernel[2][1] ~^ image[5][21] + kernel[2][2] ~^ image[5][22] + kernel[2][3] ~^ image[5][23] + kernel[2][4] ~^ image[5][24] + kernel[3][0] ~^ image[6][20] + kernel[3][1] ~^ image[6][21] + kernel[3][2] ~^ image[6][22] + kernel[3][3] ~^ image[6][23] + kernel[3][4] ~^ image[6][24] + kernel[4][0] ~^ image[7][20] + kernel[4][1] ~^ image[7][21] + kernel[4][2] ~^ image[7][22] + kernel[4][3] ~^ image[7][23] + kernel[4][4] ~^ image[7][24];
assign xor_sum[3][21] = kernel[0][0] ~^ image[3][21] + kernel[0][1] ~^ image[3][22] + kernel[0][2] ~^ image[3][23] + kernel[0][3] ~^ image[3][24] + kernel[0][4] ~^ image[3][25] + kernel[1][0] ~^ image[4][21] + kernel[1][1] ~^ image[4][22] + kernel[1][2] ~^ image[4][23] + kernel[1][3] ~^ image[4][24] + kernel[1][4] ~^ image[4][25] + kernel[2][0] ~^ image[5][21] + kernel[2][1] ~^ image[5][22] + kernel[2][2] ~^ image[5][23] + kernel[2][3] ~^ image[5][24] + kernel[2][4] ~^ image[5][25] + kernel[3][0] ~^ image[6][21] + kernel[3][1] ~^ image[6][22] + kernel[3][2] ~^ image[6][23] + kernel[3][3] ~^ image[6][24] + kernel[3][4] ~^ image[6][25] + kernel[4][0] ~^ image[7][21] + kernel[4][1] ~^ image[7][22] + kernel[4][2] ~^ image[7][23] + kernel[4][3] ~^ image[7][24] + kernel[4][4] ~^ image[7][25];
assign xor_sum[3][22] = kernel[0][0] ~^ image[3][22] + kernel[0][1] ~^ image[3][23] + kernel[0][2] ~^ image[3][24] + kernel[0][3] ~^ image[3][25] + kernel[0][4] ~^ image[3][26] + kernel[1][0] ~^ image[4][22] + kernel[1][1] ~^ image[4][23] + kernel[1][2] ~^ image[4][24] + kernel[1][3] ~^ image[4][25] + kernel[1][4] ~^ image[4][26] + kernel[2][0] ~^ image[5][22] + kernel[2][1] ~^ image[5][23] + kernel[2][2] ~^ image[5][24] + kernel[2][3] ~^ image[5][25] + kernel[2][4] ~^ image[5][26] + kernel[3][0] ~^ image[6][22] + kernel[3][1] ~^ image[6][23] + kernel[3][2] ~^ image[6][24] + kernel[3][3] ~^ image[6][25] + kernel[3][4] ~^ image[6][26] + kernel[4][0] ~^ image[7][22] + kernel[4][1] ~^ image[7][23] + kernel[4][2] ~^ image[7][24] + kernel[4][3] ~^ image[7][25] + kernel[4][4] ~^ image[7][26];
assign xor_sum[3][23] = kernel[0][0] ~^ image[3][23] + kernel[0][1] ~^ image[3][24] + kernel[0][2] ~^ image[3][25] + kernel[0][3] ~^ image[3][26] + kernel[0][4] ~^ image[3][27] + kernel[1][0] ~^ image[4][23] + kernel[1][1] ~^ image[4][24] + kernel[1][2] ~^ image[4][25] + kernel[1][3] ~^ image[4][26] + kernel[1][4] ~^ image[4][27] + kernel[2][0] ~^ image[5][23] + kernel[2][1] ~^ image[5][24] + kernel[2][2] ~^ image[5][25] + kernel[2][3] ~^ image[5][26] + kernel[2][4] ~^ image[5][27] + kernel[3][0] ~^ image[6][23] + kernel[3][1] ~^ image[6][24] + kernel[3][2] ~^ image[6][25] + kernel[3][3] ~^ image[6][26] + kernel[3][4] ~^ image[6][27] + kernel[4][0] ~^ image[7][23] + kernel[4][1] ~^ image[7][24] + kernel[4][2] ~^ image[7][25] + kernel[4][3] ~^ image[7][26] + kernel[4][4] ~^ image[7][27];
assign xor_sum[4][0] = kernel[0][0] ~^ image[4][0] + kernel[0][1] ~^ image[4][1] + kernel[0][2] ~^ image[4][2] + kernel[0][3] ~^ image[4][3] + kernel[0][4] ~^ image[4][4] + kernel[1][0] ~^ image[5][0] + kernel[1][1] ~^ image[5][1] + kernel[1][2] ~^ image[5][2] + kernel[1][3] ~^ image[5][3] + kernel[1][4] ~^ image[5][4] + kernel[2][0] ~^ image[6][0] + kernel[2][1] ~^ image[6][1] + kernel[2][2] ~^ image[6][2] + kernel[2][3] ~^ image[6][3] + kernel[2][4] ~^ image[6][4] + kernel[3][0] ~^ image[7][0] + kernel[3][1] ~^ image[7][1] + kernel[3][2] ~^ image[7][2] + kernel[3][3] ~^ image[7][3] + kernel[3][4] ~^ image[7][4] + kernel[4][0] ~^ image[8][0] + kernel[4][1] ~^ image[8][1] + kernel[4][2] ~^ image[8][2] + kernel[4][3] ~^ image[8][3] + kernel[4][4] ~^ image[8][4];
assign xor_sum[4][1] = kernel[0][0] ~^ image[4][1] + kernel[0][1] ~^ image[4][2] + kernel[0][2] ~^ image[4][3] + kernel[0][3] ~^ image[4][4] + kernel[0][4] ~^ image[4][5] + kernel[1][0] ~^ image[5][1] + kernel[1][1] ~^ image[5][2] + kernel[1][2] ~^ image[5][3] + kernel[1][3] ~^ image[5][4] + kernel[1][4] ~^ image[5][5] + kernel[2][0] ~^ image[6][1] + kernel[2][1] ~^ image[6][2] + kernel[2][2] ~^ image[6][3] + kernel[2][3] ~^ image[6][4] + kernel[2][4] ~^ image[6][5] + kernel[3][0] ~^ image[7][1] + kernel[3][1] ~^ image[7][2] + kernel[3][2] ~^ image[7][3] + kernel[3][3] ~^ image[7][4] + kernel[3][4] ~^ image[7][5] + kernel[4][0] ~^ image[8][1] + kernel[4][1] ~^ image[8][2] + kernel[4][2] ~^ image[8][3] + kernel[4][3] ~^ image[8][4] + kernel[4][4] ~^ image[8][5];
assign xor_sum[4][2] = kernel[0][0] ~^ image[4][2] + kernel[0][1] ~^ image[4][3] + kernel[0][2] ~^ image[4][4] + kernel[0][3] ~^ image[4][5] + kernel[0][4] ~^ image[4][6] + kernel[1][0] ~^ image[5][2] + kernel[1][1] ~^ image[5][3] + kernel[1][2] ~^ image[5][4] + kernel[1][3] ~^ image[5][5] + kernel[1][4] ~^ image[5][6] + kernel[2][0] ~^ image[6][2] + kernel[2][1] ~^ image[6][3] + kernel[2][2] ~^ image[6][4] + kernel[2][3] ~^ image[6][5] + kernel[2][4] ~^ image[6][6] + kernel[3][0] ~^ image[7][2] + kernel[3][1] ~^ image[7][3] + kernel[3][2] ~^ image[7][4] + kernel[3][3] ~^ image[7][5] + kernel[3][4] ~^ image[7][6] + kernel[4][0] ~^ image[8][2] + kernel[4][1] ~^ image[8][3] + kernel[4][2] ~^ image[8][4] + kernel[4][3] ~^ image[8][5] + kernel[4][4] ~^ image[8][6];
assign xor_sum[4][3] = kernel[0][0] ~^ image[4][3] + kernel[0][1] ~^ image[4][4] + kernel[0][2] ~^ image[4][5] + kernel[0][3] ~^ image[4][6] + kernel[0][4] ~^ image[4][7] + kernel[1][0] ~^ image[5][3] + kernel[1][1] ~^ image[5][4] + kernel[1][2] ~^ image[5][5] + kernel[1][3] ~^ image[5][6] + kernel[1][4] ~^ image[5][7] + kernel[2][0] ~^ image[6][3] + kernel[2][1] ~^ image[6][4] + kernel[2][2] ~^ image[6][5] + kernel[2][3] ~^ image[6][6] + kernel[2][4] ~^ image[6][7] + kernel[3][0] ~^ image[7][3] + kernel[3][1] ~^ image[7][4] + kernel[3][2] ~^ image[7][5] + kernel[3][3] ~^ image[7][6] + kernel[3][4] ~^ image[7][7] + kernel[4][0] ~^ image[8][3] + kernel[4][1] ~^ image[8][4] + kernel[4][2] ~^ image[8][5] + kernel[4][3] ~^ image[8][6] + kernel[4][4] ~^ image[8][7];
assign xor_sum[4][4] = kernel[0][0] ~^ image[4][4] + kernel[0][1] ~^ image[4][5] + kernel[0][2] ~^ image[4][6] + kernel[0][3] ~^ image[4][7] + kernel[0][4] ~^ image[4][8] + kernel[1][0] ~^ image[5][4] + kernel[1][1] ~^ image[5][5] + kernel[1][2] ~^ image[5][6] + kernel[1][3] ~^ image[5][7] + kernel[1][4] ~^ image[5][8] + kernel[2][0] ~^ image[6][4] + kernel[2][1] ~^ image[6][5] + kernel[2][2] ~^ image[6][6] + kernel[2][3] ~^ image[6][7] + kernel[2][4] ~^ image[6][8] + kernel[3][0] ~^ image[7][4] + kernel[3][1] ~^ image[7][5] + kernel[3][2] ~^ image[7][6] + kernel[3][3] ~^ image[7][7] + kernel[3][4] ~^ image[7][8] + kernel[4][0] ~^ image[8][4] + kernel[4][1] ~^ image[8][5] + kernel[4][2] ~^ image[8][6] + kernel[4][3] ~^ image[8][7] + kernel[4][4] ~^ image[8][8];
assign xor_sum[4][5] = kernel[0][0] ~^ image[4][5] + kernel[0][1] ~^ image[4][6] + kernel[0][2] ~^ image[4][7] + kernel[0][3] ~^ image[4][8] + kernel[0][4] ~^ image[4][9] + kernel[1][0] ~^ image[5][5] + kernel[1][1] ~^ image[5][6] + kernel[1][2] ~^ image[5][7] + kernel[1][3] ~^ image[5][8] + kernel[1][4] ~^ image[5][9] + kernel[2][0] ~^ image[6][5] + kernel[2][1] ~^ image[6][6] + kernel[2][2] ~^ image[6][7] + kernel[2][3] ~^ image[6][8] + kernel[2][4] ~^ image[6][9] + kernel[3][0] ~^ image[7][5] + kernel[3][1] ~^ image[7][6] + kernel[3][2] ~^ image[7][7] + kernel[3][3] ~^ image[7][8] + kernel[3][4] ~^ image[7][9] + kernel[4][0] ~^ image[8][5] + kernel[4][1] ~^ image[8][6] + kernel[4][2] ~^ image[8][7] + kernel[4][3] ~^ image[8][8] + kernel[4][4] ~^ image[8][9];
assign xor_sum[4][6] = kernel[0][0] ~^ image[4][6] + kernel[0][1] ~^ image[4][7] + kernel[0][2] ~^ image[4][8] + kernel[0][3] ~^ image[4][9] + kernel[0][4] ~^ image[4][10] + kernel[1][0] ~^ image[5][6] + kernel[1][1] ~^ image[5][7] + kernel[1][2] ~^ image[5][8] + kernel[1][3] ~^ image[5][9] + kernel[1][4] ~^ image[5][10] + kernel[2][0] ~^ image[6][6] + kernel[2][1] ~^ image[6][7] + kernel[2][2] ~^ image[6][8] + kernel[2][3] ~^ image[6][9] + kernel[2][4] ~^ image[6][10] + kernel[3][0] ~^ image[7][6] + kernel[3][1] ~^ image[7][7] + kernel[3][2] ~^ image[7][8] + kernel[3][3] ~^ image[7][9] + kernel[3][4] ~^ image[7][10] + kernel[4][0] ~^ image[8][6] + kernel[4][1] ~^ image[8][7] + kernel[4][2] ~^ image[8][8] + kernel[4][3] ~^ image[8][9] + kernel[4][4] ~^ image[8][10];
assign xor_sum[4][7] = kernel[0][0] ~^ image[4][7] + kernel[0][1] ~^ image[4][8] + kernel[0][2] ~^ image[4][9] + kernel[0][3] ~^ image[4][10] + kernel[0][4] ~^ image[4][11] + kernel[1][0] ~^ image[5][7] + kernel[1][1] ~^ image[5][8] + kernel[1][2] ~^ image[5][9] + kernel[1][3] ~^ image[5][10] + kernel[1][4] ~^ image[5][11] + kernel[2][0] ~^ image[6][7] + kernel[2][1] ~^ image[6][8] + kernel[2][2] ~^ image[6][9] + kernel[2][3] ~^ image[6][10] + kernel[2][4] ~^ image[6][11] + kernel[3][0] ~^ image[7][7] + kernel[3][1] ~^ image[7][8] + kernel[3][2] ~^ image[7][9] + kernel[3][3] ~^ image[7][10] + kernel[3][4] ~^ image[7][11] + kernel[4][0] ~^ image[8][7] + kernel[4][1] ~^ image[8][8] + kernel[4][2] ~^ image[8][9] + kernel[4][3] ~^ image[8][10] + kernel[4][4] ~^ image[8][11];
assign xor_sum[4][8] = kernel[0][0] ~^ image[4][8] + kernel[0][1] ~^ image[4][9] + kernel[0][2] ~^ image[4][10] + kernel[0][3] ~^ image[4][11] + kernel[0][4] ~^ image[4][12] + kernel[1][0] ~^ image[5][8] + kernel[1][1] ~^ image[5][9] + kernel[1][2] ~^ image[5][10] + kernel[1][3] ~^ image[5][11] + kernel[1][4] ~^ image[5][12] + kernel[2][0] ~^ image[6][8] + kernel[2][1] ~^ image[6][9] + kernel[2][2] ~^ image[6][10] + kernel[2][3] ~^ image[6][11] + kernel[2][4] ~^ image[6][12] + kernel[3][0] ~^ image[7][8] + kernel[3][1] ~^ image[7][9] + kernel[3][2] ~^ image[7][10] + kernel[3][3] ~^ image[7][11] + kernel[3][4] ~^ image[7][12] + kernel[4][0] ~^ image[8][8] + kernel[4][1] ~^ image[8][9] + kernel[4][2] ~^ image[8][10] + kernel[4][3] ~^ image[8][11] + kernel[4][4] ~^ image[8][12];
assign xor_sum[4][9] = kernel[0][0] ~^ image[4][9] + kernel[0][1] ~^ image[4][10] + kernel[0][2] ~^ image[4][11] + kernel[0][3] ~^ image[4][12] + kernel[0][4] ~^ image[4][13] + kernel[1][0] ~^ image[5][9] + kernel[1][1] ~^ image[5][10] + kernel[1][2] ~^ image[5][11] + kernel[1][3] ~^ image[5][12] + kernel[1][4] ~^ image[5][13] + kernel[2][0] ~^ image[6][9] + kernel[2][1] ~^ image[6][10] + kernel[2][2] ~^ image[6][11] + kernel[2][3] ~^ image[6][12] + kernel[2][4] ~^ image[6][13] + kernel[3][0] ~^ image[7][9] + kernel[3][1] ~^ image[7][10] + kernel[3][2] ~^ image[7][11] + kernel[3][3] ~^ image[7][12] + kernel[3][4] ~^ image[7][13] + kernel[4][0] ~^ image[8][9] + kernel[4][1] ~^ image[8][10] + kernel[4][2] ~^ image[8][11] + kernel[4][3] ~^ image[8][12] + kernel[4][4] ~^ image[8][13];
assign xor_sum[4][10] = kernel[0][0] ~^ image[4][10] + kernel[0][1] ~^ image[4][11] + kernel[0][2] ~^ image[4][12] + kernel[0][3] ~^ image[4][13] + kernel[0][4] ~^ image[4][14] + kernel[1][0] ~^ image[5][10] + kernel[1][1] ~^ image[5][11] + kernel[1][2] ~^ image[5][12] + kernel[1][3] ~^ image[5][13] + kernel[1][4] ~^ image[5][14] + kernel[2][0] ~^ image[6][10] + kernel[2][1] ~^ image[6][11] + kernel[2][2] ~^ image[6][12] + kernel[2][3] ~^ image[6][13] + kernel[2][4] ~^ image[6][14] + kernel[3][0] ~^ image[7][10] + kernel[3][1] ~^ image[7][11] + kernel[3][2] ~^ image[7][12] + kernel[3][3] ~^ image[7][13] + kernel[3][4] ~^ image[7][14] + kernel[4][0] ~^ image[8][10] + kernel[4][1] ~^ image[8][11] + kernel[4][2] ~^ image[8][12] + kernel[4][3] ~^ image[8][13] + kernel[4][4] ~^ image[8][14];
assign xor_sum[4][11] = kernel[0][0] ~^ image[4][11] + kernel[0][1] ~^ image[4][12] + kernel[0][2] ~^ image[4][13] + kernel[0][3] ~^ image[4][14] + kernel[0][4] ~^ image[4][15] + kernel[1][0] ~^ image[5][11] + kernel[1][1] ~^ image[5][12] + kernel[1][2] ~^ image[5][13] + kernel[1][3] ~^ image[5][14] + kernel[1][4] ~^ image[5][15] + kernel[2][0] ~^ image[6][11] + kernel[2][1] ~^ image[6][12] + kernel[2][2] ~^ image[6][13] + kernel[2][3] ~^ image[6][14] + kernel[2][4] ~^ image[6][15] + kernel[3][0] ~^ image[7][11] + kernel[3][1] ~^ image[7][12] + kernel[3][2] ~^ image[7][13] + kernel[3][3] ~^ image[7][14] + kernel[3][4] ~^ image[7][15] + kernel[4][0] ~^ image[8][11] + kernel[4][1] ~^ image[8][12] + kernel[4][2] ~^ image[8][13] + kernel[4][3] ~^ image[8][14] + kernel[4][4] ~^ image[8][15];
assign xor_sum[4][12] = kernel[0][0] ~^ image[4][12] + kernel[0][1] ~^ image[4][13] + kernel[0][2] ~^ image[4][14] + kernel[0][3] ~^ image[4][15] + kernel[0][4] ~^ image[4][16] + kernel[1][0] ~^ image[5][12] + kernel[1][1] ~^ image[5][13] + kernel[1][2] ~^ image[5][14] + kernel[1][3] ~^ image[5][15] + kernel[1][4] ~^ image[5][16] + kernel[2][0] ~^ image[6][12] + kernel[2][1] ~^ image[6][13] + kernel[2][2] ~^ image[6][14] + kernel[2][3] ~^ image[6][15] + kernel[2][4] ~^ image[6][16] + kernel[3][0] ~^ image[7][12] + kernel[3][1] ~^ image[7][13] + kernel[3][2] ~^ image[7][14] + kernel[3][3] ~^ image[7][15] + kernel[3][4] ~^ image[7][16] + kernel[4][0] ~^ image[8][12] + kernel[4][1] ~^ image[8][13] + kernel[4][2] ~^ image[8][14] + kernel[4][3] ~^ image[8][15] + kernel[4][4] ~^ image[8][16];
assign xor_sum[4][13] = kernel[0][0] ~^ image[4][13] + kernel[0][1] ~^ image[4][14] + kernel[0][2] ~^ image[4][15] + kernel[0][3] ~^ image[4][16] + kernel[0][4] ~^ image[4][17] + kernel[1][0] ~^ image[5][13] + kernel[1][1] ~^ image[5][14] + kernel[1][2] ~^ image[5][15] + kernel[1][3] ~^ image[5][16] + kernel[1][4] ~^ image[5][17] + kernel[2][0] ~^ image[6][13] + kernel[2][1] ~^ image[6][14] + kernel[2][2] ~^ image[6][15] + kernel[2][3] ~^ image[6][16] + kernel[2][4] ~^ image[6][17] + kernel[3][0] ~^ image[7][13] + kernel[3][1] ~^ image[7][14] + kernel[3][2] ~^ image[7][15] + kernel[3][3] ~^ image[7][16] + kernel[3][4] ~^ image[7][17] + kernel[4][0] ~^ image[8][13] + kernel[4][1] ~^ image[8][14] + kernel[4][2] ~^ image[8][15] + kernel[4][3] ~^ image[8][16] + kernel[4][4] ~^ image[8][17];
assign xor_sum[4][14] = kernel[0][0] ~^ image[4][14] + kernel[0][1] ~^ image[4][15] + kernel[0][2] ~^ image[4][16] + kernel[0][3] ~^ image[4][17] + kernel[0][4] ~^ image[4][18] + kernel[1][0] ~^ image[5][14] + kernel[1][1] ~^ image[5][15] + kernel[1][2] ~^ image[5][16] + kernel[1][3] ~^ image[5][17] + kernel[1][4] ~^ image[5][18] + kernel[2][0] ~^ image[6][14] + kernel[2][1] ~^ image[6][15] + kernel[2][2] ~^ image[6][16] + kernel[2][3] ~^ image[6][17] + kernel[2][4] ~^ image[6][18] + kernel[3][0] ~^ image[7][14] + kernel[3][1] ~^ image[7][15] + kernel[3][2] ~^ image[7][16] + kernel[3][3] ~^ image[7][17] + kernel[3][4] ~^ image[7][18] + kernel[4][0] ~^ image[8][14] + kernel[4][1] ~^ image[8][15] + kernel[4][2] ~^ image[8][16] + kernel[4][3] ~^ image[8][17] + kernel[4][4] ~^ image[8][18];
assign xor_sum[4][15] = kernel[0][0] ~^ image[4][15] + kernel[0][1] ~^ image[4][16] + kernel[0][2] ~^ image[4][17] + kernel[0][3] ~^ image[4][18] + kernel[0][4] ~^ image[4][19] + kernel[1][0] ~^ image[5][15] + kernel[1][1] ~^ image[5][16] + kernel[1][2] ~^ image[5][17] + kernel[1][3] ~^ image[5][18] + kernel[1][4] ~^ image[5][19] + kernel[2][0] ~^ image[6][15] + kernel[2][1] ~^ image[6][16] + kernel[2][2] ~^ image[6][17] + kernel[2][3] ~^ image[6][18] + kernel[2][4] ~^ image[6][19] + kernel[3][0] ~^ image[7][15] + kernel[3][1] ~^ image[7][16] + kernel[3][2] ~^ image[7][17] + kernel[3][3] ~^ image[7][18] + kernel[3][4] ~^ image[7][19] + kernel[4][0] ~^ image[8][15] + kernel[4][1] ~^ image[8][16] + kernel[4][2] ~^ image[8][17] + kernel[4][3] ~^ image[8][18] + kernel[4][4] ~^ image[8][19];
assign xor_sum[4][16] = kernel[0][0] ~^ image[4][16] + kernel[0][1] ~^ image[4][17] + kernel[0][2] ~^ image[4][18] + kernel[0][3] ~^ image[4][19] + kernel[0][4] ~^ image[4][20] + kernel[1][0] ~^ image[5][16] + kernel[1][1] ~^ image[5][17] + kernel[1][2] ~^ image[5][18] + kernel[1][3] ~^ image[5][19] + kernel[1][4] ~^ image[5][20] + kernel[2][0] ~^ image[6][16] + kernel[2][1] ~^ image[6][17] + kernel[2][2] ~^ image[6][18] + kernel[2][3] ~^ image[6][19] + kernel[2][4] ~^ image[6][20] + kernel[3][0] ~^ image[7][16] + kernel[3][1] ~^ image[7][17] + kernel[3][2] ~^ image[7][18] + kernel[3][3] ~^ image[7][19] + kernel[3][4] ~^ image[7][20] + kernel[4][0] ~^ image[8][16] + kernel[4][1] ~^ image[8][17] + kernel[4][2] ~^ image[8][18] + kernel[4][3] ~^ image[8][19] + kernel[4][4] ~^ image[8][20];
assign xor_sum[4][17] = kernel[0][0] ~^ image[4][17] + kernel[0][1] ~^ image[4][18] + kernel[0][2] ~^ image[4][19] + kernel[0][3] ~^ image[4][20] + kernel[0][4] ~^ image[4][21] + kernel[1][0] ~^ image[5][17] + kernel[1][1] ~^ image[5][18] + kernel[1][2] ~^ image[5][19] + kernel[1][3] ~^ image[5][20] + kernel[1][4] ~^ image[5][21] + kernel[2][0] ~^ image[6][17] + kernel[2][1] ~^ image[6][18] + kernel[2][2] ~^ image[6][19] + kernel[2][3] ~^ image[6][20] + kernel[2][4] ~^ image[6][21] + kernel[3][0] ~^ image[7][17] + kernel[3][1] ~^ image[7][18] + kernel[3][2] ~^ image[7][19] + kernel[3][3] ~^ image[7][20] + kernel[3][4] ~^ image[7][21] + kernel[4][0] ~^ image[8][17] + kernel[4][1] ~^ image[8][18] + kernel[4][2] ~^ image[8][19] + kernel[4][3] ~^ image[8][20] + kernel[4][4] ~^ image[8][21];
assign xor_sum[4][18] = kernel[0][0] ~^ image[4][18] + kernel[0][1] ~^ image[4][19] + kernel[0][2] ~^ image[4][20] + kernel[0][3] ~^ image[4][21] + kernel[0][4] ~^ image[4][22] + kernel[1][0] ~^ image[5][18] + kernel[1][1] ~^ image[5][19] + kernel[1][2] ~^ image[5][20] + kernel[1][3] ~^ image[5][21] + kernel[1][4] ~^ image[5][22] + kernel[2][0] ~^ image[6][18] + kernel[2][1] ~^ image[6][19] + kernel[2][2] ~^ image[6][20] + kernel[2][3] ~^ image[6][21] + kernel[2][4] ~^ image[6][22] + kernel[3][0] ~^ image[7][18] + kernel[3][1] ~^ image[7][19] + kernel[3][2] ~^ image[7][20] + kernel[3][3] ~^ image[7][21] + kernel[3][4] ~^ image[7][22] + kernel[4][0] ~^ image[8][18] + kernel[4][1] ~^ image[8][19] + kernel[4][2] ~^ image[8][20] + kernel[4][3] ~^ image[8][21] + kernel[4][4] ~^ image[8][22];
assign xor_sum[4][19] = kernel[0][0] ~^ image[4][19] + kernel[0][1] ~^ image[4][20] + kernel[0][2] ~^ image[4][21] + kernel[0][3] ~^ image[4][22] + kernel[0][4] ~^ image[4][23] + kernel[1][0] ~^ image[5][19] + kernel[1][1] ~^ image[5][20] + kernel[1][2] ~^ image[5][21] + kernel[1][3] ~^ image[5][22] + kernel[1][4] ~^ image[5][23] + kernel[2][0] ~^ image[6][19] + kernel[2][1] ~^ image[6][20] + kernel[2][2] ~^ image[6][21] + kernel[2][3] ~^ image[6][22] + kernel[2][4] ~^ image[6][23] + kernel[3][0] ~^ image[7][19] + kernel[3][1] ~^ image[7][20] + kernel[3][2] ~^ image[7][21] + kernel[3][3] ~^ image[7][22] + kernel[3][4] ~^ image[7][23] + kernel[4][0] ~^ image[8][19] + kernel[4][1] ~^ image[8][20] + kernel[4][2] ~^ image[8][21] + kernel[4][3] ~^ image[8][22] + kernel[4][4] ~^ image[8][23];
assign xor_sum[4][20] = kernel[0][0] ~^ image[4][20] + kernel[0][1] ~^ image[4][21] + kernel[0][2] ~^ image[4][22] + kernel[0][3] ~^ image[4][23] + kernel[0][4] ~^ image[4][24] + kernel[1][0] ~^ image[5][20] + kernel[1][1] ~^ image[5][21] + kernel[1][2] ~^ image[5][22] + kernel[1][3] ~^ image[5][23] + kernel[1][4] ~^ image[5][24] + kernel[2][0] ~^ image[6][20] + kernel[2][1] ~^ image[6][21] + kernel[2][2] ~^ image[6][22] + kernel[2][3] ~^ image[6][23] + kernel[2][4] ~^ image[6][24] + kernel[3][0] ~^ image[7][20] + kernel[3][1] ~^ image[7][21] + kernel[3][2] ~^ image[7][22] + kernel[3][3] ~^ image[7][23] + kernel[3][4] ~^ image[7][24] + kernel[4][0] ~^ image[8][20] + kernel[4][1] ~^ image[8][21] + kernel[4][2] ~^ image[8][22] + kernel[4][3] ~^ image[8][23] + kernel[4][4] ~^ image[8][24];
assign xor_sum[4][21] = kernel[0][0] ~^ image[4][21] + kernel[0][1] ~^ image[4][22] + kernel[0][2] ~^ image[4][23] + kernel[0][3] ~^ image[4][24] + kernel[0][4] ~^ image[4][25] + kernel[1][0] ~^ image[5][21] + kernel[1][1] ~^ image[5][22] + kernel[1][2] ~^ image[5][23] + kernel[1][3] ~^ image[5][24] + kernel[1][4] ~^ image[5][25] + kernel[2][0] ~^ image[6][21] + kernel[2][1] ~^ image[6][22] + kernel[2][2] ~^ image[6][23] + kernel[2][3] ~^ image[6][24] + kernel[2][4] ~^ image[6][25] + kernel[3][0] ~^ image[7][21] + kernel[3][1] ~^ image[7][22] + kernel[3][2] ~^ image[7][23] + kernel[3][3] ~^ image[7][24] + kernel[3][4] ~^ image[7][25] + kernel[4][0] ~^ image[8][21] + kernel[4][1] ~^ image[8][22] + kernel[4][2] ~^ image[8][23] + kernel[4][3] ~^ image[8][24] + kernel[4][4] ~^ image[8][25];
assign xor_sum[4][22] = kernel[0][0] ~^ image[4][22] + kernel[0][1] ~^ image[4][23] + kernel[0][2] ~^ image[4][24] + kernel[0][3] ~^ image[4][25] + kernel[0][4] ~^ image[4][26] + kernel[1][0] ~^ image[5][22] + kernel[1][1] ~^ image[5][23] + kernel[1][2] ~^ image[5][24] + kernel[1][3] ~^ image[5][25] + kernel[1][4] ~^ image[5][26] + kernel[2][0] ~^ image[6][22] + kernel[2][1] ~^ image[6][23] + kernel[2][2] ~^ image[6][24] + kernel[2][3] ~^ image[6][25] + kernel[2][4] ~^ image[6][26] + kernel[3][0] ~^ image[7][22] + kernel[3][1] ~^ image[7][23] + kernel[3][2] ~^ image[7][24] + kernel[3][3] ~^ image[7][25] + kernel[3][4] ~^ image[7][26] + kernel[4][0] ~^ image[8][22] + kernel[4][1] ~^ image[8][23] + kernel[4][2] ~^ image[8][24] + kernel[4][3] ~^ image[8][25] + kernel[4][4] ~^ image[8][26];
assign xor_sum[4][23] = kernel[0][0] ~^ image[4][23] + kernel[0][1] ~^ image[4][24] + kernel[0][2] ~^ image[4][25] + kernel[0][3] ~^ image[4][26] + kernel[0][4] ~^ image[4][27] + kernel[1][0] ~^ image[5][23] + kernel[1][1] ~^ image[5][24] + kernel[1][2] ~^ image[5][25] + kernel[1][3] ~^ image[5][26] + kernel[1][4] ~^ image[5][27] + kernel[2][0] ~^ image[6][23] + kernel[2][1] ~^ image[6][24] + kernel[2][2] ~^ image[6][25] + kernel[2][3] ~^ image[6][26] + kernel[2][4] ~^ image[6][27] + kernel[3][0] ~^ image[7][23] + kernel[3][1] ~^ image[7][24] + kernel[3][2] ~^ image[7][25] + kernel[3][3] ~^ image[7][26] + kernel[3][4] ~^ image[7][27] + kernel[4][0] ~^ image[8][23] + kernel[4][1] ~^ image[8][24] + kernel[4][2] ~^ image[8][25] + kernel[4][3] ~^ image[8][26] + kernel[4][4] ~^ image[8][27];
assign xor_sum[5][0] = kernel[0][0] ~^ image[5][0] + kernel[0][1] ~^ image[5][1] + kernel[0][2] ~^ image[5][2] + kernel[0][3] ~^ image[5][3] + kernel[0][4] ~^ image[5][4] + kernel[1][0] ~^ image[6][0] + kernel[1][1] ~^ image[6][1] + kernel[1][2] ~^ image[6][2] + kernel[1][3] ~^ image[6][3] + kernel[1][4] ~^ image[6][4] + kernel[2][0] ~^ image[7][0] + kernel[2][1] ~^ image[7][1] + kernel[2][2] ~^ image[7][2] + kernel[2][3] ~^ image[7][3] + kernel[2][4] ~^ image[7][4] + kernel[3][0] ~^ image[8][0] + kernel[3][1] ~^ image[8][1] + kernel[3][2] ~^ image[8][2] + kernel[3][3] ~^ image[8][3] + kernel[3][4] ~^ image[8][4] + kernel[4][0] ~^ image[9][0] + kernel[4][1] ~^ image[9][1] + kernel[4][2] ~^ image[9][2] + kernel[4][3] ~^ image[9][3] + kernel[4][4] ~^ image[9][4];
assign xor_sum[5][1] = kernel[0][0] ~^ image[5][1] + kernel[0][1] ~^ image[5][2] + kernel[0][2] ~^ image[5][3] + kernel[0][3] ~^ image[5][4] + kernel[0][4] ~^ image[5][5] + kernel[1][0] ~^ image[6][1] + kernel[1][1] ~^ image[6][2] + kernel[1][2] ~^ image[6][3] + kernel[1][3] ~^ image[6][4] + kernel[1][4] ~^ image[6][5] + kernel[2][0] ~^ image[7][1] + kernel[2][1] ~^ image[7][2] + kernel[2][2] ~^ image[7][3] + kernel[2][3] ~^ image[7][4] + kernel[2][4] ~^ image[7][5] + kernel[3][0] ~^ image[8][1] + kernel[3][1] ~^ image[8][2] + kernel[3][2] ~^ image[8][3] + kernel[3][3] ~^ image[8][4] + kernel[3][4] ~^ image[8][5] + kernel[4][0] ~^ image[9][1] + kernel[4][1] ~^ image[9][2] + kernel[4][2] ~^ image[9][3] + kernel[4][3] ~^ image[9][4] + kernel[4][4] ~^ image[9][5];
assign xor_sum[5][2] = kernel[0][0] ~^ image[5][2] + kernel[0][1] ~^ image[5][3] + kernel[0][2] ~^ image[5][4] + kernel[0][3] ~^ image[5][5] + kernel[0][4] ~^ image[5][6] + kernel[1][0] ~^ image[6][2] + kernel[1][1] ~^ image[6][3] + kernel[1][2] ~^ image[6][4] + kernel[1][3] ~^ image[6][5] + kernel[1][4] ~^ image[6][6] + kernel[2][0] ~^ image[7][2] + kernel[2][1] ~^ image[7][3] + kernel[2][2] ~^ image[7][4] + kernel[2][3] ~^ image[7][5] + kernel[2][4] ~^ image[7][6] + kernel[3][0] ~^ image[8][2] + kernel[3][1] ~^ image[8][3] + kernel[3][2] ~^ image[8][4] + kernel[3][3] ~^ image[8][5] + kernel[3][4] ~^ image[8][6] + kernel[4][0] ~^ image[9][2] + kernel[4][1] ~^ image[9][3] + kernel[4][2] ~^ image[9][4] + kernel[4][3] ~^ image[9][5] + kernel[4][4] ~^ image[9][6];
assign xor_sum[5][3] = kernel[0][0] ~^ image[5][3] + kernel[0][1] ~^ image[5][4] + kernel[0][2] ~^ image[5][5] + kernel[0][3] ~^ image[5][6] + kernel[0][4] ~^ image[5][7] + kernel[1][0] ~^ image[6][3] + kernel[1][1] ~^ image[6][4] + kernel[1][2] ~^ image[6][5] + kernel[1][3] ~^ image[6][6] + kernel[1][4] ~^ image[6][7] + kernel[2][0] ~^ image[7][3] + kernel[2][1] ~^ image[7][4] + kernel[2][2] ~^ image[7][5] + kernel[2][3] ~^ image[7][6] + kernel[2][4] ~^ image[7][7] + kernel[3][0] ~^ image[8][3] + kernel[3][1] ~^ image[8][4] + kernel[3][2] ~^ image[8][5] + kernel[3][3] ~^ image[8][6] + kernel[3][4] ~^ image[8][7] + kernel[4][0] ~^ image[9][3] + kernel[4][1] ~^ image[9][4] + kernel[4][2] ~^ image[9][5] + kernel[4][3] ~^ image[9][6] + kernel[4][4] ~^ image[9][7];
assign xor_sum[5][4] = kernel[0][0] ~^ image[5][4] + kernel[0][1] ~^ image[5][5] + kernel[0][2] ~^ image[5][6] + kernel[0][3] ~^ image[5][7] + kernel[0][4] ~^ image[5][8] + kernel[1][0] ~^ image[6][4] + kernel[1][1] ~^ image[6][5] + kernel[1][2] ~^ image[6][6] + kernel[1][3] ~^ image[6][7] + kernel[1][4] ~^ image[6][8] + kernel[2][0] ~^ image[7][4] + kernel[2][1] ~^ image[7][5] + kernel[2][2] ~^ image[7][6] + kernel[2][3] ~^ image[7][7] + kernel[2][4] ~^ image[7][8] + kernel[3][0] ~^ image[8][4] + kernel[3][1] ~^ image[8][5] + kernel[3][2] ~^ image[8][6] + kernel[3][3] ~^ image[8][7] + kernel[3][4] ~^ image[8][8] + kernel[4][0] ~^ image[9][4] + kernel[4][1] ~^ image[9][5] + kernel[4][2] ~^ image[9][6] + kernel[4][3] ~^ image[9][7] + kernel[4][4] ~^ image[9][8];
assign xor_sum[5][5] = kernel[0][0] ~^ image[5][5] + kernel[0][1] ~^ image[5][6] + kernel[0][2] ~^ image[5][7] + kernel[0][3] ~^ image[5][8] + kernel[0][4] ~^ image[5][9] + kernel[1][0] ~^ image[6][5] + kernel[1][1] ~^ image[6][6] + kernel[1][2] ~^ image[6][7] + kernel[1][3] ~^ image[6][8] + kernel[1][4] ~^ image[6][9] + kernel[2][0] ~^ image[7][5] + kernel[2][1] ~^ image[7][6] + kernel[2][2] ~^ image[7][7] + kernel[2][3] ~^ image[7][8] + kernel[2][4] ~^ image[7][9] + kernel[3][0] ~^ image[8][5] + kernel[3][1] ~^ image[8][6] + kernel[3][2] ~^ image[8][7] + kernel[3][3] ~^ image[8][8] + kernel[3][4] ~^ image[8][9] + kernel[4][0] ~^ image[9][5] + kernel[4][1] ~^ image[9][6] + kernel[4][2] ~^ image[9][7] + kernel[4][3] ~^ image[9][8] + kernel[4][4] ~^ image[9][9];
assign xor_sum[5][6] = kernel[0][0] ~^ image[5][6] + kernel[0][1] ~^ image[5][7] + kernel[0][2] ~^ image[5][8] + kernel[0][3] ~^ image[5][9] + kernel[0][4] ~^ image[5][10] + kernel[1][0] ~^ image[6][6] + kernel[1][1] ~^ image[6][7] + kernel[1][2] ~^ image[6][8] + kernel[1][3] ~^ image[6][9] + kernel[1][4] ~^ image[6][10] + kernel[2][0] ~^ image[7][6] + kernel[2][1] ~^ image[7][7] + kernel[2][2] ~^ image[7][8] + kernel[2][3] ~^ image[7][9] + kernel[2][4] ~^ image[7][10] + kernel[3][0] ~^ image[8][6] + kernel[3][1] ~^ image[8][7] + kernel[3][2] ~^ image[8][8] + kernel[3][3] ~^ image[8][9] + kernel[3][4] ~^ image[8][10] + kernel[4][0] ~^ image[9][6] + kernel[4][1] ~^ image[9][7] + kernel[4][2] ~^ image[9][8] + kernel[4][3] ~^ image[9][9] + kernel[4][4] ~^ image[9][10];
assign xor_sum[5][7] = kernel[0][0] ~^ image[5][7] + kernel[0][1] ~^ image[5][8] + kernel[0][2] ~^ image[5][9] + kernel[0][3] ~^ image[5][10] + kernel[0][4] ~^ image[5][11] + kernel[1][0] ~^ image[6][7] + kernel[1][1] ~^ image[6][8] + kernel[1][2] ~^ image[6][9] + kernel[1][3] ~^ image[6][10] + kernel[1][4] ~^ image[6][11] + kernel[2][0] ~^ image[7][7] + kernel[2][1] ~^ image[7][8] + kernel[2][2] ~^ image[7][9] + kernel[2][3] ~^ image[7][10] + kernel[2][4] ~^ image[7][11] + kernel[3][0] ~^ image[8][7] + kernel[3][1] ~^ image[8][8] + kernel[3][2] ~^ image[8][9] + kernel[3][3] ~^ image[8][10] + kernel[3][4] ~^ image[8][11] + kernel[4][0] ~^ image[9][7] + kernel[4][1] ~^ image[9][8] + kernel[4][2] ~^ image[9][9] + kernel[4][3] ~^ image[9][10] + kernel[4][4] ~^ image[9][11];
assign xor_sum[5][8] = kernel[0][0] ~^ image[5][8] + kernel[0][1] ~^ image[5][9] + kernel[0][2] ~^ image[5][10] + kernel[0][3] ~^ image[5][11] + kernel[0][4] ~^ image[5][12] + kernel[1][0] ~^ image[6][8] + kernel[1][1] ~^ image[6][9] + kernel[1][2] ~^ image[6][10] + kernel[1][3] ~^ image[6][11] + kernel[1][4] ~^ image[6][12] + kernel[2][0] ~^ image[7][8] + kernel[2][1] ~^ image[7][9] + kernel[2][2] ~^ image[7][10] + kernel[2][3] ~^ image[7][11] + kernel[2][4] ~^ image[7][12] + kernel[3][0] ~^ image[8][8] + kernel[3][1] ~^ image[8][9] + kernel[3][2] ~^ image[8][10] + kernel[3][3] ~^ image[8][11] + kernel[3][4] ~^ image[8][12] + kernel[4][0] ~^ image[9][8] + kernel[4][1] ~^ image[9][9] + kernel[4][2] ~^ image[9][10] + kernel[4][3] ~^ image[9][11] + kernel[4][4] ~^ image[9][12];
assign xor_sum[5][9] = kernel[0][0] ~^ image[5][9] + kernel[0][1] ~^ image[5][10] + kernel[0][2] ~^ image[5][11] + kernel[0][3] ~^ image[5][12] + kernel[0][4] ~^ image[5][13] + kernel[1][0] ~^ image[6][9] + kernel[1][1] ~^ image[6][10] + kernel[1][2] ~^ image[6][11] + kernel[1][3] ~^ image[6][12] + kernel[1][4] ~^ image[6][13] + kernel[2][0] ~^ image[7][9] + kernel[2][1] ~^ image[7][10] + kernel[2][2] ~^ image[7][11] + kernel[2][3] ~^ image[7][12] + kernel[2][4] ~^ image[7][13] + kernel[3][0] ~^ image[8][9] + kernel[3][1] ~^ image[8][10] + kernel[3][2] ~^ image[8][11] + kernel[3][3] ~^ image[8][12] + kernel[3][4] ~^ image[8][13] + kernel[4][0] ~^ image[9][9] + kernel[4][1] ~^ image[9][10] + kernel[4][2] ~^ image[9][11] + kernel[4][3] ~^ image[9][12] + kernel[4][4] ~^ image[9][13];
assign xor_sum[5][10] = kernel[0][0] ~^ image[5][10] + kernel[0][1] ~^ image[5][11] + kernel[0][2] ~^ image[5][12] + kernel[0][3] ~^ image[5][13] + kernel[0][4] ~^ image[5][14] + kernel[1][0] ~^ image[6][10] + kernel[1][1] ~^ image[6][11] + kernel[1][2] ~^ image[6][12] + kernel[1][3] ~^ image[6][13] + kernel[1][4] ~^ image[6][14] + kernel[2][0] ~^ image[7][10] + kernel[2][1] ~^ image[7][11] + kernel[2][2] ~^ image[7][12] + kernel[2][3] ~^ image[7][13] + kernel[2][4] ~^ image[7][14] + kernel[3][0] ~^ image[8][10] + kernel[3][1] ~^ image[8][11] + kernel[3][2] ~^ image[8][12] + kernel[3][3] ~^ image[8][13] + kernel[3][4] ~^ image[8][14] + kernel[4][0] ~^ image[9][10] + kernel[4][1] ~^ image[9][11] + kernel[4][2] ~^ image[9][12] + kernel[4][3] ~^ image[9][13] + kernel[4][4] ~^ image[9][14];
assign xor_sum[5][11] = kernel[0][0] ~^ image[5][11] + kernel[0][1] ~^ image[5][12] + kernel[0][2] ~^ image[5][13] + kernel[0][3] ~^ image[5][14] + kernel[0][4] ~^ image[5][15] + kernel[1][0] ~^ image[6][11] + kernel[1][1] ~^ image[6][12] + kernel[1][2] ~^ image[6][13] + kernel[1][3] ~^ image[6][14] + kernel[1][4] ~^ image[6][15] + kernel[2][0] ~^ image[7][11] + kernel[2][1] ~^ image[7][12] + kernel[2][2] ~^ image[7][13] + kernel[2][3] ~^ image[7][14] + kernel[2][4] ~^ image[7][15] + kernel[3][0] ~^ image[8][11] + kernel[3][1] ~^ image[8][12] + kernel[3][2] ~^ image[8][13] + kernel[3][3] ~^ image[8][14] + kernel[3][4] ~^ image[8][15] + kernel[4][0] ~^ image[9][11] + kernel[4][1] ~^ image[9][12] + kernel[4][2] ~^ image[9][13] + kernel[4][3] ~^ image[9][14] + kernel[4][4] ~^ image[9][15];
assign xor_sum[5][12] = kernel[0][0] ~^ image[5][12] + kernel[0][1] ~^ image[5][13] + kernel[0][2] ~^ image[5][14] + kernel[0][3] ~^ image[5][15] + kernel[0][4] ~^ image[5][16] + kernel[1][0] ~^ image[6][12] + kernel[1][1] ~^ image[6][13] + kernel[1][2] ~^ image[6][14] + kernel[1][3] ~^ image[6][15] + kernel[1][4] ~^ image[6][16] + kernel[2][0] ~^ image[7][12] + kernel[2][1] ~^ image[7][13] + kernel[2][2] ~^ image[7][14] + kernel[2][3] ~^ image[7][15] + kernel[2][4] ~^ image[7][16] + kernel[3][0] ~^ image[8][12] + kernel[3][1] ~^ image[8][13] + kernel[3][2] ~^ image[8][14] + kernel[3][3] ~^ image[8][15] + kernel[3][4] ~^ image[8][16] + kernel[4][0] ~^ image[9][12] + kernel[4][1] ~^ image[9][13] + kernel[4][2] ~^ image[9][14] + kernel[4][3] ~^ image[9][15] + kernel[4][4] ~^ image[9][16];
assign xor_sum[5][13] = kernel[0][0] ~^ image[5][13] + kernel[0][1] ~^ image[5][14] + kernel[0][2] ~^ image[5][15] + kernel[0][3] ~^ image[5][16] + kernel[0][4] ~^ image[5][17] + kernel[1][0] ~^ image[6][13] + kernel[1][1] ~^ image[6][14] + kernel[1][2] ~^ image[6][15] + kernel[1][3] ~^ image[6][16] + kernel[1][4] ~^ image[6][17] + kernel[2][0] ~^ image[7][13] + kernel[2][1] ~^ image[7][14] + kernel[2][2] ~^ image[7][15] + kernel[2][3] ~^ image[7][16] + kernel[2][4] ~^ image[7][17] + kernel[3][0] ~^ image[8][13] + kernel[3][1] ~^ image[8][14] + kernel[3][2] ~^ image[8][15] + kernel[3][3] ~^ image[8][16] + kernel[3][4] ~^ image[8][17] + kernel[4][0] ~^ image[9][13] + kernel[4][1] ~^ image[9][14] + kernel[4][2] ~^ image[9][15] + kernel[4][3] ~^ image[9][16] + kernel[4][4] ~^ image[9][17];
assign xor_sum[5][14] = kernel[0][0] ~^ image[5][14] + kernel[0][1] ~^ image[5][15] + kernel[0][2] ~^ image[5][16] + kernel[0][3] ~^ image[5][17] + kernel[0][4] ~^ image[5][18] + kernel[1][0] ~^ image[6][14] + kernel[1][1] ~^ image[6][15] + kernel[1][2] ~^ image[6][16] + kernel[1][3] ~^ image[6][17] + kernel[1][4] ~^ image[6][18] + kernel[2][0] ~^ image[7][14] + kernel[2][1] ~^ image[7][15] + kernel[2][2] ~^ image[7][16] + kernel[2][3] ~^ image[7][17] + kernel[2][4] ~^ image[7][18] + kernel[3][0] ~^ image[8][14] + kernel[3][1] ~^ image[8][15] + kernel[3][2] ~^ image[8][16] + kernel[3][3] ~^ image[8][17] + kernel[3][4] ~^ image[8][18] + kernel[4][0] ~^ image[9][14] + kernel[4][1] ~^ image[9][15] + kernel[4][2] ~^ image[9][16] + kernel[4][3] ~^ image[9][17] + kernel[4][4] ~^ image[9][18];
assign xor_sum[5][15] = kernel[0][0] ~^ image[5][15] + kernel[0][1] ~^ image[5][16] + kernel[0][2] ~^ image[5][17] + kernel[0][3] ~^ image[5][18] + kernel[0][4] ~^ image[5][19] + kernel[1][0] ~^ image[6][15] + kernel[1][1] ~^ image[6][16] + kernel[1][2] ~^ image[6][17] + kernel[1][3] ~^ image[6][18] + kernel[1][4] ~^ image[6][19] + kernel[2][0] ~^ image[7][15] + kernel[2][1] ~^ image[7][16] + kernel[2][2] ~^ image[7][17] + kernel[2][3] ~^ image[7][18] + kernel[2][4] ~^ image[7][19] + kernel[3][0] ~^ image[8][15] + kernel[3][1] ~^ image[8][16] + kernel[3][2] ~^ image[8][17] + kernel[3][3] ~^ image[8][18] + kernel[3][4] ~^ image[8][19] + kernel[4][0] ~^ image[9][15] + kernel[4][1] ~^ image[9][16] + kernel[4][2] ~^ image[9][17] + kernel[4][3] ~^ image[9][18] + kernel[4][4] ~^ image[9][19];
assign xor_sum[5][16] = kernel[0][0] ~^ image[5][16] + kernel[0][1] ~^ image[5][17] + kernel[0][2] ~^ image[5][18] + kernel[0][3] ~^ image[5][19] + kernel[0][4] ~^ image[5][20] + kernel[1][0] ~^ image[6][16] + kernel[1][1] ~^ image[6][17] + kernel[1][2] ~^ image[6][18] + kernel[1][3] ~^ image[6][19] + kernel[1][4] ~^ image[6][20] + kernel[2][0] ~^ image[7][16] + kernel[2][1] ~^ image[7][17] + kernel[2][2] ~^ image[7][18] + kernel[2][3] ~^ image[7][19] + kernel[2][4] ~^ image[7][20] + kernel[3][0] ~^ image[8][16] + kernel[3][1] ~^ image[8][17] + kernel[3][2] ~^ image[8][18] + kernel[3][3] ~^ image[8][19] + kernel[3][4] ~^ image[8][20] + kernel[4][0] ~^ image[9][16] + kernel[4][1] ~^ image[9][17] + kernel[4][2] ~^ image[9][18] + kernel[4][3] ~^ image[9][19] + kernel[4][4] ~^ image[9][20];
assign xor_sum[5][17] = kernel[0][0] ~^ image[5][17] + kernel[0][1] ~^ image[5][18] + kernel[0][2] ~^ image[5][19] + kernel[0][3] ~^ image[5][20] + kernel[0][4] ~^ image[5][21] + kernel[1][0] ~^ image[6][17] + kernel[1][1] ~^ image[6][18] + kernel[1][2] ~^ image[6][19] + kernel[1][3] ~^ image[6][20] + kernel[1][4] ~^ image[6][21] + kernel[2][0] ~^ image[7][17] + kernel[2][1] ~^ image[7][18] + kernel[2][2] ~^ image[7][19] + kernel[2][3] ~^ image[7][20] + kernel[2][4] ~^ image[7][21] + kernel[3][0] ~^ image[8][17] + kernel[3][1] ~^ image[8][18] + kernel[3][2] ~^ image[8][19] + kernel[3][3] ~^ image[8][20] + kernel[3][4] ~^ image[8][21] + kernel[4][0] ~^ image[9][17] + kernel[4][1] ~^ image[9][18] + kernel[4][2] ~^ image[9][19] + kernel[4][3] ~^ image[9][20] + kernel[4][4] ~^ image[9][21];
assign xor_sum[5][18] = kernel[0][0] ~^ image[5][18] + kernel[0][1] ~^ image[5][19] + kernel[0][2] ~^ image[5][20] + kernel[0][3] ~^ image[5][21] + kernel[0][4] ~^ image[5][22] + kernel[1][0] ~^ image[6][18] + kernel[1][1] ~^ image[6][19] + kernel[1][2] ~^ image[6][20] + kernel[1][3] ~^ image[6][21] + kernel[1][4] ~^ image[6][22] + kernel[2][0] ~^ image[7][18] + kernel[2][1] ~^ image[7][19] + kernel[2][2] ~^ image[7][20] + kernel[2][3] ~^ image[7][21] + kernel[2][4] ~^ image[7][22] + kernel[3][0] ~^ image[8][18] + kernel[3][1] ~^ image[8][19] + kernel[3][2] ~^ image[8][20] + kernel[3][3] ~^ image[8][21] + kernel[3][4] ~^ image[8][22] + kernel[4][0] ~^ image[9][18] + kernel[4][1] ~^ image[9][19] + kernel[4][2] ~^ image[9][20] + kernel[4][3] ~^ image[9][21] + kernel[4][4] ~^ image[9][22];
assign xor_sum[5][19] = kernel[0][0] ~^ image[5][19] + kernel[0][1] ~^ image[5][20] + kernel[0][2] ~^ image[5][21] + kernel[0][3] ~^ image[5][22] + kernel[0][4] ~^ image[5][23] + kernel[1][0] ~^ image[6][19] + kernel[1][1] ~^ image[6][20] + kernel[1][2] ~^ image[6][21] + kernel[1][3] ~^ image[6][22] + kernel[1][4] ~^ image[6][23] + kernel[2][0] ~^ image[7][19] + kernel[2][1] ~^ image[7][20] + kernel[2][2] ~^ image[7][21] + kernel[2][3] ~^ image[7][22] + kernel[2][4] ~^ image[7][23] + kernel[3][0] ~^ image[8][19] + kernel[3][1] ~^ image[8][20] + kernel[3][2] ~^ image[8][21] + kernel[3][3] ~^ image[8][22] + kernel[3][4] ~^ image[8][23] + kernel[4][0] ~^ image[9][19] + kernel[4][1] ~^ image[9][20] + kernel[4][2] ~^ image[9][21] + kernel[4][3] ~^ image[9][22] + kernel[4][4] ~^ image[9][23];
assign xor_sum[5][20] = kernel[0][0] ~^ image[5][20] + kernel[0][1] ~^ image[5][21] + kernel[0][2] ~^ image[5][22] + kernel[0][3] ~^ image[5][23] + kernel[0][4] ~^ image[5][24] + kernel[1][0] ~^ image[6][20] + kernel[1][1] ~^ image[6][21] + kernel[1][2] ~^ image[6][22] + kernel[1][3] ~^ image[6][23] + kernel[1][4] ~^ image[6][24] + kernel[2][0] ~^ image[7][20] + kernel[2][1] ~^ image[7][21] + kernel[2][2] ~^ image[7][22] + kernel[2][3] ~^ image[7][23] + kernel[2][4] ~^ image[7][24] + kernel[3][0] ~^ image[8][20] + kernel[3][1] ~^ image[8][21] + kernel[3][2] ~^ image[8][22] + kernel[3][3] ~^ image[8][23] + kernel[3][4] ~^ image[8][24] + kernel[4][0] ~^ image[9][20] + kernel[4][1] ~^ image[9][21] + kernel[4][2] ~^ image[9][22] + kernel[4][3] ~^ image[9][23] + kernel[4][4] ~^ image[9][24];
assign xor_sum[5][21] = kernel[0][0] ~^ image[5][21] + kernel[0][1] ~^ image[5][22] + kernel[0][2] ~^ image[5][23] + kernel[0][3] ~^ image[5][24] + kernel[0][4] ~^ image[5][25] + kernel[1][0] ~^ image[6][21] + kernel[1][1] ~^ image[6][22] + kernel[1][2] ~^ image[6][23] + kernel[1][3] ~^ image[6][24] + kernel[1][4] ~^ image[6][25] + kernel[2][0] ~^ image[7][21] + kernel[2][1] ~^ image[7][22] + kernel[2][2] ~^ image[7][23] + kernel[2][3] ~^ image[7][24] + kernel[2][4] ~^ image[7][25] + kernel[3][0] ~^ image[8][21] + kernel[3][1] ~^ image[8][22] + kernel[3][2] ~^ image[8][23] + kernel[3][3] ~^ image[8][24] + kernel[3][4] ~^ image[8][25] + kernel[4][0] ~^ image[9][21] + kernel[4][1] ~^ image[9][22] + kernel[4][2] ~^ image[9][23] + kernel[4][3] ~^ image[9][24] + kernel[4][4] ~^ image[9][25];
assign xor_sum[5][22] = kernel[0][0] ~^ image[5][22] + kernel[0][1] ~^ image[5][23] + kernel[0][2] ~^ image[5][24] + kernel[0][3] ~^ image[5][25] + kernel[0][4] ~^ image[5][26] + kernel[1][0] ~^ image[6][22] + kernel[1][1] ~^ image[6][23] + kernel[1][2] ~^ image[6][24] + kernel[1][3] ~^ image[6][25] + kernel[1][4] ~^ image[6][26] + kernel[2][0] ~^ image[7][22] + kernel[2][1] ~^ image[7][23] + kernel[2][2] ~^ image[7][24] + kernel[2][3] ~^ image[7][25] + kernel[2][4] ~^ image[7][26] + kernel[3][0] ~^ image[8][22] + kernel[3][1] ~^ image[8][23] + kernel[3][2] ~^ image[8][24] + kernel[3][3] ~^ image[8][25] + kernel[3][4] ~^ image[8][26] + kernel[4][0] ~^ image[9][22] + kernel[4][1] ~^ image[9][23] + kernel[4][2] ~^ image[9][24] + kernel[4][3] ~^ image[9][25] + kernel[4][4] ~^ image[9][26];
assign xor_sum[5][23] = kernel[0][0] ~^ image[5][23] + kernel[0][1] ~^ image[5][24] + kernel[0][2] ~^ image[5][25] + kernel[0][3] ~^ image[5][26] + kernel[0][4] ~^ image[5][27] + kernel[1][0] ~^ image[6][23] + kernel[1][1] ~^ image[6][24] + kernel[1][2] ~^ image[6][25] + kernel[1][3] ~^ image[6][26] + kernel[1][4] ~^ image[6][27] + kernel[2][0] ~^ image[7][23] + kernel[2][1] ~^ image[7][24] + kernel[2][2] ~^ image[7][25] + kernel[2][3] ~^ image[7][26] + kernel[2][4] ~^ image[7][27] + kernel[3][0] ~^ image[8][23] + kernel[3][1] ~^ image[8][24] + kernel[3][2] ~^ image[8][25] + kernel[3][3] ~^ image[8][26] + kernel[3][4] ~^ image[8][27] + kernel[4][0] ~^ image[9][23] + kernel[4][1] ~^ image[9][24] + kernel[4][2] ~^ image[9][25] + kernel[4][3] ~^ image[9][26] + kernel[4][4] ~^ image[9][27];
assign xor_sum[6][0] = kernel[0][0] ~^ image[6][0] + kernel[0][1] ~^ image[6][1] + kernel[0][2] ~^ image[6][2] + kernel[0][3] ~^ image[6][3] + kernel[0][4] ~^ image[6][4] + kernel[1][0] ~^ image[7][0] + kernel[1][1] ~^ image[7][1] + kernel[1][2] ~^ image[7][2] + kernel[1][3] ~^ image[7][3] + kernel[1][4] ~^ image[7][4] + kernel[2][0] ~^ image[8][0] + kernel[2][1] ~^ image[8][1] + kernel[2][2] ~^ image[8][2] + kernel[2][3] ~^ image[8][3] + kernel[2][4] ~^ image[8][4] + kernel[3][0] ~^ image[9][0] + kernel[3][1] ~^ image[9][1] + kernel[3][2] ~^ image[9][2] + kernel[3][3] ~^ image[9][3] + kernel[3][4] ~^ image[9][4] + kernel[4][0] ~^ image[10][0] + kernel[4][1] ~^ image[10][1] + kernel[4][2] ~^ image[10][2] + kernel[4][3] ~^ image[10][3] + kernel[4][4] ~^ image[10][4];
assign xor_sum[6][1] = kernel[0][0] ~^ image[6][1] + kernel[0][1] ~^ image[6][2] + kernel[0][2] ~^ image[6][3] + kernel[0][3] ~^ image[6][4] + kernel[0][4] ~^ image[6][5] + kernel[1][0] ~^ image[7][1] + kernel[1][1] ~^ image[7][2] + kernel[1][2] ~^ image[7][3] + kernel[1][3] ~^ image[7][4] + kernel[1][4] ~^ image[7][5] + kernel[2][0] ~^ image[8][1] + kernel[2][1] ~^ image[8][2] + kernel[2][2] ~^ image[8][3] + kernel[2][3] ~^ image[8][4] + kernel[2][4] ~^ image[8][5] + kernel[3][0] ~^ image[9][1] + kernel[3][1] ~^ image[9][2] + kernel[3][2] ~^ image[9][3] + kernel[3][3] ~^ image[9][4] + kernel[3][4] ~^ image[9][5] + kernel[4][0] ~^ image[10][1] + kernel[4][1] ~^ image[10][2] + kernel[4][2] ~^ image[10][3] + kernel[4][3] ~^ image[10][4] + kernel[4][4] ~^ image[10][5];
assign xor_sum[6][2] = kernel[0][0] ~^ image[6][2] + kernel[0][1] ~^ image[6][3] + kernel[0][2] ~^ image[6][4] + kernel[0][3] ~^ image[6][5] + kernel[0][4] ~^ image[6][6] + kernel[1][0] ~^ image[7][2] + kernel[1][1] ~^ image[7][3] + kernel[1][2] ~^ image[7][4] + kernel[1][3] ~^ image[7][5] + kernel[1][4] ~^ image[7][6] + kernel[2][0] ~^ image[8][2] + kernel[2][1] ~^ image[8][3] + kernel[2][2] ~^ image[8][4] + kernel[2][3] ~^ image[8][5] + kernel[2][4] ~^ image[8][6] + kernel[3][0] ~^ image[9][2] + kernel[3][1] ~^ image[9][3] + kernel[3][2] ~^ image[9][4] + kernel[3][3] ~^ image[9][5] + kernel[3][4] ~^ image[9][6] + kernel[4][0] ~^ image[10][2] + kernel[4][1] ~^ image[10][3] + kernel[4][2] ~^ image[10][4] + kernel[4][3] ~^ image[10][5] + kernel[4][4] ~^ image[10][6];
assign xor_sum[6][3] = kernel[0][0] ~^ image[6][3] + kernel[0][1] ~^ image[6][4] + kernel[0][2] ~^ image[6][5] + kernel[0][3] ~^ image[6][6] + kernel[0][4] ~^ image[6][7] + kernel[1][0] ~^ image[7][3] + kernel[1][1] ~^ image[7][4] + kernel[1][2] ~^ image[7][5] + kernel[1][3] ~^ image[7][6] + kernel[1][4] ~^ image[7][7] + kernel[2][0] ~^ image[8][3] + kernel[2][1] ~^ image[8][4] + kernel[2][2] ~^ image[8][5] + kernel[2][3] ~^ image[8][6] + kernel[2][4] ~^ image[8][7] + kernel[3][0] ~^ image[9][3] + kernel[3][1] ~^ image[9][4] + kernel[3][2] ~^ image[9][5] + kernel[3][3] ~^ image[9][6] + kernel[3][4] ~^ image[9][7] + kernel[4][0] ~^ image[10][3] + kernel[4][1] ~^ image[10][4] + kernel[4][2] ~^ image[10][5] + kernel[4][3] ~^ image[10][6] + kernel[4][4] ~^ image[10][7];
assign xor_sum[6][4] = kernel[0][0] ~^ image[6][4] + kernel[0][1] ~^ image[6][5] + kernel[0][2] ~^ image[6][6] + kernel[0][3] ~^ image[6][7] + kernel[0][4] ~^ image[6][8] + kernel[1][0] ~^ image[7][4] + kernel[1][1] ~^ image[7][5] + kernel[1][2] ~^ image[7][6] + kernel[1][3] ~^ image[7][7] + kernel[1][4] ~^ image[7][8] + kernel[2][0] ~^ image[8][4] + kernel[2][1] ~^ image[8][5] + kernel[2][2] ~^ image[8][6] + kernel[2][3] ~^ image[8][7] + kernel[2][4] ~^ image[8][8] + kernel[3][0] ~^ image[9][4] + kernel[3][1] ~^ image[9][5] + kernel[3][2] ~^ image[9][6] + kernel[3][3] ~^ image[9][7] + kernel[3][4] ~^ image[9][8] + kernel[4][0] ~^ image[10][4] + kernel[4][1] ~^ image[10][5] + kernel[4][2] ~^ image[10][6] + kernel[4][3] ~^ image[10][7] + kernel[4][4] ~^ image[10][8];
assign xor_sum[6][5] = kernel[0][0] ~^ image[6][5] + kernel[0][1] ~^ image[6][6] + kernel[0][2] ~^ image[6][7] + kernel[0][3] ~^ image[6][8] + kernel[0][4] ~^ image[6][9] + kernel[1][0] ~^ image[7][5] + kernel[1][1] ~^ image[7][6] + kernel[1][2] ~^ image[7][7] + kernel[1][3] ~^ image[7][8] + kernel[1][4] ~^ image[7][9] + kernel[2][0] ~^ image[8][5] + kernel[2][1] ~^ image[8][6] + kernel[2][2] ~^ image[8][7] + kernel[2][3] ~^ image[8][8] + kernel[2][4] ~^ image[8][9] + kernel[3][0] ~^ image[9][5] + kernel[3][1] ~^ image[9][6] + kernel[3][2] ~^ image[9][7] + kernel[3][3] ~^ image[9][8] + kernel[3][4] ~^ image[9][9] + kernel[4][0] ~^ image[10][5] + kernel[4][1] ~^ image[10][6] + kernel[4][2] ~^ image[10][7] + kernel[4][3] ~^ image[10][8] + kernel[4][4] ~^ image[10][9];
assign xor_sum[6][6] = kernel[0][0] ~^ image[6][6] + kernel[0][1] ~^ image[6][7] + kernel[0][2] ~^ image[6][8] + kernel[0][3] ~^ image[6][9] + kernel[0][4] ~^ image[6][10] + kernel[1][0] ~^ image[7][6] + kernel[1][1] ~^ image[7][7] + kernel[1][2] ~^ image[7][8] + kernel[1][3] ~^ image[7][9] + kernel[1][4] ~^ image[7][10] + kernel[2][0] ~^ image[8][6] + kernel[2][1] ~^ image[8][7] + kernel[2][2] ~^ image[8][8] + kernel[2][3] ~^ image[8][9] + kernel[2][4] ~^ image[8][10] + kernel[3][0] ~^ image[9][6] + kernel[3][1] ~^ image[9][7] + kernel[3][2] ~^ image[9][8] + kernel[3][3] ~^ image[9][9] + kernel[3][4] ~^ image[9][10] + kernel[4][0] ~^ image[10][6] + kernel[4][1] ~^ image[10][7] + kernel[4][2] ~^ image[10][8] + kernel[4][3] ~^ image[10][9] + kernel[4][4] ~^ image[10][10];
assign xor_sum[6][7] = kernel[0][0] ~^ image[6][7] + kernel[0][1] ~^ image[6][8] + kernel[0][2] ~^ image[6][9] + kernel[0][3] ~^ image[6][10] + kernel[0][4] ~^ image[6][11] + kernel[1][0] ~^ image[7][7] + kernel[1][1] ~^ image[7][8] + kernel[1][2] ~^ image[7][9] + kernel[1][3] ~^ image[7][10] + kernel[1][4] ~^ image[7][11] + kernel[2][0] ~^ image[8][7] + kernel[2][1] ~^ image[8][8] + kernel[2][2] ~^ image[8][9] + kernel[2][3] ~^ image[8][10] + kernel[2][4] ~^ image[8][11] + kernel[3][0] ~^ image[9][7] + kernel[3][1] ~^ image[9][8] + kernel[3][2] ~^ image[9][9] + kernel[3][3] ~^ image[9][10] + kernel[3][4] ~^ image[9][11] + kernel[4][0] ~^ image[10][7] + kernel[4][1] ~^ image[10][8] + kernel[4][2] ~^ image[10][9] + kernel[4][3] ~^ image[10][10] + kernel[4][4] ~^ image[10][11];
assign xor_sum[6][8] = kernel[0][0] ~^ image[6][8] + kernel[0][1] ~^ image[6][9] + kernel[0][2] ~^ image[6][10] + kernel[0][3] ~^ image[6][11] + kernel[0][4] ~^ image[6][12] + kernel[1][0] ~^ image[7][8] + kernel[1][1] ~^ image[7][9] + kernel[1][2] ~^ image[7][10] + kernel[1][3] ~^ image[7][11] + kernel[1][4] ~^ image[7][12] + kernel[2][0] ~^ image[8][8] + kernel[2][1] ~^ image[8][9] + kernel[2][2] ~^ image[8][10] + kernel[2][3] ~^ image[8][11] + kernel[2][4] ~^ image[8][12] + kernel[3][0] ~^ image[9][8] + kernel[3][1] ~^ image[9][9] + kernel[3][2] ~^ image[9][10] + kernel[3][3] ~^ image[9][11] + kernel[3][4] ~^ image[9][12] + kernel[4][0] ~^ image[10][8] + kernel[4][1] ~^ image[10][9] + kernel[4][2] ~^ image[10][10] + kernel[4][3] ~^ image[10][11] + kernel[4][4] ~^ image[10][12];
assign xor_sum[6][9] = kernel[0][0] ~^ image[6][9] + kernel[0][1] ~^ image[6][10] + kernel[0][2] ~^ image[6][11] + kernel[0][3] ~^ image[6][12] + kernel[0][4] ~^ image[6][13] + kernel[1][0] ~^ image[7][9] + kernel[1][1] ~^ image[7][10] + kernel[1][2] ~^ image[7][11] + kernel[1][3] ~^ image[7][12] + kernel[1][4] ~^ image[7][13] + kernel[2][0] ~^ image[8][9] + kernel[2][1] ~^ image[8][10] + kernel[2][2] ~^ image[8][11] + kernel[2][3] ~^ image[8][12] + kernel[2][4] ~^ image[8][13] + kernel[3][0] ~^ image[9][9] + kernel[3][1] ~^ image[9][10] + kernel[3][2] ~^ image[9][11] + kernel[3][3] ~^ image[9][12] + kernel[3][4] ~^ image[9][13] + kernel[4][0] ~^ image[10][9] + kernel[4][1] ~^ image[10][10] + kernel[4][2] ~^ image[10][11] + kernel[4][3] ~^ image[10][12] + kernel[4][4] ~^ image[10][13];
assign xor_sum[6][10] = kernel[0][0] ~^ image[6][10] + kernel[0][1] ~^ image[6][11] + kernel[0][2] ~^ image[6][12] + kernel[0][3] ~^ image[6][13] + kernel[0][4] ~^ image[6][14] + kernel[1][0] ~^ image[7][10] + kernel[1][1] ~^ image[7][11] + kernel[1][2] ~^ image[7][12] + kernel[1][3] ~^ image[7][13] + kernel[1][4] ~^ image[7][14] + kernel[2][0] ~^ image[8][10] + kernel[2][1] ~^ image[8][11] + kernel[2][2] ~^ image[8][12] + kernel[2][3] ~^ image[8][13] + kernel[2][4] ~^ image[8][14] + kernel[3][0] ~^ image[9][10] + kernel[3][1] ~^ image[9][11] + kernel[3][2] ~^ image[9][12] + kernel[3][3] ~^ image[9][13] + kernel[3][4] ~^ image[9][14] + kernel[4][0] ~^ image[10][10] + kernel[4][1] ~^ image[10][11] + kernel[4][2] ~^ image[10][12] + kernel[4][3] ~^ image[10][13] + kernel[4][4] ~^ image[10][14];
assign xor_sum[6][11] = kernel[0][0] ~^ image[6][11] + kernel[0][1] ~^ image[6][12] + kernel[0][2] ~^ image[6][13] + kernel[0][3] ~^ image[6][14] + kernel[0][4] ~^ image[6][15] + kernel[1][0] ~^ image[7][11] + kernel[1][1] ~^ image[7][12] + kernel[1][2] ~^ image[7][13] + kernel[1][3] ~^ image[7][14] + kernel[1][4] ~^ image[7][15] + kernel[2][0] ~^ image[8][11] + kernel[2][1] ~^ image[8][12] + kernel[2][2] ~^ image[8][13] + kernel[2][3] ~^ image[8][14] + kernel[2][4] ~^ image[8][15] + kernel[3][0] ~^ image[9][11] + kernel[3][1] ~^ image[9][12] + kernel[3][2] ~^ image[9][13] + kernel[3][3] ~^ image[9][14] + kernel[3][4] ~^ image[9][15] + kernel[4][0] ~^ image[10][11] + kernel[4][1] ~^ image[10][12] + kernel[4][2] ~^ image[10][13] + kernel[4][3] ~^ image[10][14] + kernel[4][4] ~^ image[10][15];
assign xor_sum[6][12] = kernel[0][0] ~^ image[6][12] + kernel[0][1] ~^ image[6][13] + kernel[0][2] ~^ image[6][14] + kernel[0][3] ~^ image[6][15] + kernel[0][4] ~^ image[6][16] + kernel[1][0] ~^ image[7][12] + kernel[1][1] ~^ image[7][13] + kernel[1][2] ~^ image[7][14] + kernel[1][3] ~^ image[7][15] + kernel[1][4] ~^ image[7][16] + kernel[2][0] ~^ image[8][12] + kernel[2][1] ~^ image[8][13] + kernel[2][2] ~^ image[8][14] + kernel[2][3] ~^ image[8][15] + kernel[2][4] ~^ image[8][16] + kernel[3][0] ~^ image[9][12] + kernel[3][1] ~^ image[9][13] + kernel[3][2] ~^ image[9][14] + kernel[3][3] ~^ image[9][15] + kernel[3][4] ~^ image[9][16] + kernel[4][0] ~^ image[10][12] + kernel[4][1] ~^ image[10][13] + kernel[4][2] ~^ image[10][14] + kernel[4][3] ~^ image[10][15] + kernel[4][4] ~^ image[10][16];
assign xor_sum[6][13] = kernel[0][0] ~^ image[6][13] + kernel[0][1] ~^ image[6][14] + kernel[0][2] ~^ image[6][15] + kernel[0][3] ~^ image[6][16] + kernel[0][4] ~^ image[6][17] + kernel[1][0] ~^ image[7][13] + kernel[1][1] ~^ image[7][14] + kernel[1][2] ~^ image[7][15] + kernel[1][3] ~^ image[7][16] + kernel[1][4] ~^ image[7][17] + kernel[2][0] ~^ image[8][13] + kernel[2][1] ~^ image[8][14] + kernel[2][2] ~^ image[8][15] + kernel[2][3] ~^ image[8][16] + kernel[2][4] ~^ image[8][17] + kernel[3][0] ~^ image[9][13] + kernel[3][1] ~^ image[9][14] + kernel[3][2] ~^ image[9][15] + kernel[3][3] ~^ image[9][16] + kernel[3][4] ~^ image[9][17] + kernel[4][0] ~^ image[10][13] + kernel[4][1] ~^ image[10][14] + kernel[4][2] ~^ image[10][15] + kernel[4][3] ~^ image[10][16] + kernel[4][4] ~^ image[10][17];
assign xor_sum[6][14] = kernel[0][0] ~^ image[6][14] + kernel[0][1] ~^ image[6][15] + kernel[0][2] ~^ image[6][16] + kernel[0][3] ~^ image[6][17] + kernel[0][4] ~^ image[6][18] + kernel[1][0] ~^ image[7][14] + kernel[1][1] ~^ image[7][15] + kernel[1][2] ~^ image[7][16] + kernel[1][3] ~^ image[7][17] + kernel[1][4] ~^ image[7][18] + kernel[2][0] ~^ image[8][14] + kernel[2][1] ~^ image[8][15] + kernel[2][2] ~^ image[8][16] + kernel[2][3] ~^ image[8][17] + kernel[2][4] ~^ image[8][18] + kernel[3][0] ~^ image[9][14] + kernel[3][1] ~^ image[9][15] + kernel[3][2] ~^ image[9][16] + kernel[3][3] ~^ image[9][17] + kernel[3][4] ~^ image[9][18] + kernel[4][0] ~^ image[10][14] + kernel[4][1] ~^ image[10][15] + kernel[4][2] ~^ image[10][16] + kernel[4][3] ~^ image[10][17] + kernel[4][4] ~^ image[10][18];
assign xor_sum[6][15] = kernel[0][0] ~^ image[6][15] + kernel[0][1] ~^ image[6][16] + kernel[0][2] ~^ image[6][17] + kernel[0][3] ~^ image[6][18] + kernel[0][4] ~^ image[6][19] + kernel[1][0] ~^ image[7][15] + kernel[1][1] ~^ image[7][16] + kernel[1][2] ~^ image[7][17] + kernel[1][3] ~^ image[7][18] + kernel[1][4] ~^ image[7][19] + kernel[2][0] ~^ image[8][15] + kernel[2][1] ~^ image[8][16] + kernel[2][2] ~^ image[8][17] + kernel[2][3] ~^ image[8][18] + kernel[2][4] ~^ image[8][19] + kernel[3][0] ~^ image[9][15] + kernel[3][1] ~^ image[9][16] + kernel[3][2] ~^ image[9][17] + kernel[3][3] ~^ image[9][18] + kernel[3][4] ~^ image[9][19] + kernel[4][0] ~^ image[10][15] + kernel[4][1] ~^ image[10][16] + kernel[4][2] ~^ image[10][17] + kernel[4][3] ~^ image[10][18] + kernel[4][4] ~^ image[10][19];
assign xor_sum[6][16] = kernel[0][0] ~^ image[6][16] + kernel[0][1] ~^ image[6][17] + kernel[0][2] ~^ image[6][18] + kernel[0][3] ~^ image[6][19] + kernel[0][4] ~^ image[6][20] + kernel[1][0] ~^ image[7][16] + kernel[1][1] ~^ image[7][17] + kernel[1][2] ~^ image[7][18] + kernel[1][3] ~^ image[7][19] + kernel[1][4] ~^ image[7][20] + kernel[2][0] ~^ image[8][16] + kernel[2][1] ~^ image[8][17] + kernel[2][2] ~^ image[8][18] + kernel[2][3] ~^ image[8][19] + kernel[2][4] ~^ image[8][20] + kernel[3][0] ~^ image[9][16] + kernel[3][1] ~^ image[9][17] + kernel[3][2] ~^ image[9][18] + kernel[3][3] ~^ image[9][19] + kernel[3][4] ~^ image[9][20] + kernel[4][0] ~^ image[10][16] + kernel[4][1] ~^ image[10][17] + kernel[4][2] ~^ image[10][18] + kernel[4][3] ~^ image[10][19] + kernel[4][4] ~^ image[10][20];
assign xor_sum[6][17] = kernel[0][0] ~^ image[6][17] + kernel[0][1] ~^ image[6][18] + kernel[0][2] ~^ image[6][19] + kernel[0][3] ~^ image[6][20] + kernel[0][4] ~^ image[6][21] + kernel[1][0] ~^ image[7][17] + kernel[1][1] ~^ image[7][18] + kernel[1][2] ~^ image[7][19] + kernel[1][3] ~^ image[7][20] + kernel[1][4] ~^ image[7][21] + kernel[2][0] ~^ image[8][17] + kernel[2][1] ~^ image[8][18] + kernel[2][2] ~^ image[8][19] + kernel[2][3] ~^ image[8][20] + kernel[2][4] ~^ image[8][21] + kernel[3][0] ~^ image[9][17] + kernel[3][1] ~^ image[9][18] + kernel[3][2] ~^ image[9][19] + kernel[3][3] ~^ image[9][20] + kernel[3][4] ~^ image[9][21] + kernel[4][0] ~^ image[10][17] + kernel[4][1] ~^ image[10][18] + kernel[4][2] ~^ image[10][19] + kernel[4][3] ~^ image[10][20] + kernel[4][4] ~^ image[10][21];
assign xor_sum[6][18] = kernel[0][0] ~^ image[6][18] + kernel[0][1] ~^ image[6][19] + kernel[0][2] ~^ image[6][20] + kernel[0][3] ~^ image[6][21] + kernel[0][4] ~^ image[6][22] + kernel[1][0] ~^ image[7][18] + kernel[1][1] ~^ image[7][19] + kernel[1][2] ~^ image[7][20] + kernel[1][3] ~^ image[7][21] + kernel[1][4] ~^ image[7][22] + kernel[2][0] ~^ image[8][18] + kernel[2][1] ~^ image[8][19] + kernel[2][2] ~^ image[8][20] + kernel[2][3] ~^ image[8][21] + kernel[2][4] ~^ image[8][22] + kernel[3][0] ~^ image[9][18] + kernel[3][1] ~^ image[9][19] + kernel[3][2] ~^ image[9][20] + kernel[3][3] ~^ image[9][21] + kernel[3][4] ~^ image[9][22] + kernel[4][0] ~^ image[10][18] + kernel[4][1] ~^ image[10][19] + kernel[4][2] ~^ image[10][20] + kernel[4][3] ~^ image[10][21] + kernel[4][4] ~^ image[10][22];
assign xor_sum[6][19] = kernel[0][0] ~^ image[6][19] + kernel[0][1] ~^ image[6][20] + kernel[0][2] ~^ image[6][21] + kernel[0][3] ~^ image[6][22] + kernel[0][4] ~^ image[6][23] + kernel[1][0] ~^ image[7][19] + kernel[1][1] ~^ image[7][20] + kernel[1][2] ~^ image[7][21] + kernel[1][3] ~^ image[7][22] + kernel[1][4] ~^ image[7][23] + kernel[2][0] ~^ image[8][19] + kernel[2][1] ~^ image[8][20] + kernel[2][2] ~^ image[8][21] + kernel[2][3] ~^ image[8][22] + kernel[2][4] ~^ image[8][23] + kernel[3][0] ~^ image[9][19] + kernel[3][1] ~^ image[9][20] + kernel[3][2] ~^ image[9][21] + kernel[3][3] ~^ image[9][22] + kernel[3][4] ~^ image[9][23] + kernel[4][0] ~^ image[10][19] + kernel[4][1] ~^ image[10][20] + kernel[4][2] ~^ image[10][21] + kernel[4][3] ~^ image[10][22] + kernel[4][4] ~^ image[10][23];
assign xor_sum[6][20] = kernel[0][0] ~^ image[6][20] + kernel[0][1] ~^ image[6][21] + kernel[0][2] ~^ image[6][22] + kernel[0][3] ~^ image[6][23] + kernel[0][4] ~^ image[6][24] + kernel[1][0] ~^ image[7][20] + kernel[1][1] ~^ image[7][21] + kernel[1][2] ~^ image[7][22] + kernel[1][3] ~^ image[7][23] + kernel[1][4] ~^ image[7][24] + kernel[2][0] ~^ image[8][20] + kernel[2][1] ~^ image[8][21] + kernel[2][2] ~^ image[8][22] + kernel[2][3] ~^ image[8][23] + kernel[2][4] ~^ image[8][24] + kernel[3][0] ~^ image[9][20] + kernel[3][1] ~^ image[9][21] + kernel[3][2] ~^ image[9][22] + kernel[3][3] ~^ image[9][23] + kernel[3][4] ~^ image[9][24] + kernel[4][0] ~^ image[10][20] + kernel[4][1] ~^ image[10][21] + kernel[4][2] ~^ image[10][22] + kernel[4][3] ~^ image[10][23] + kernel[4][4] ~^ image[10][24];
assign xor_sum[6][21] = kernel[0][0] ~^ image[6][21] + kernel[0][1] ~^ image[6][22] + kernel[0][2] ~^ image[6][23] + kernel[0][3] ~^ image[6][24] + kernel[0][4] ~^ image[6][25] + kernel[1][0] ~^ image[7][21] + kernel[1][1] ~^ image[7][22] + kernel[1][2] ~^ image[7][23] + kernel[1][3] ~^ image[7][24] + kernel[1][4] ~^ image[7][25] + kernel[2][0] ~^ image[8][21] + kernel[2][1] ~^ image[8][22] + kernel[2][2] ~^ image[8][23] + kernel[2][3] ~^ image[8][24] + kernel[2][4] ~^ image[8][25] + kernel[3][0] ~^ image[9][21] + kernel[3][1] ~^ image[9][22] + kernel[3][2] ~^ image[9][23] + kernel[3][3] ~^ image[9][24] + kernel[3][4] ~^ image[9][25] + kernel[4][0] ~^ image[10][21] + kernel[4][1] ~^ image[10][22] + kernel[4][2] ~^ image[10][23] + kernel[4][3] ~^ image[10][24] + kernel[4][4] ~^ image[10][25];
assign xor_sum[6][22] = kernel[0][0] ~^ image[6][22] + kernel[0][1] ~^ image[6][23] + kernel[0][2] ~^ image[6][24] + kernel[0][3] ~^ image[6][25] + kernel[0][4] ~^ image[6][26] + kernel[1][0] ~^ image[7][22] + kernel[1][1] ~^ image[7][23] + kernel[1][2] ~^ image[7][24] + kernel[1][3] ~^ image[7][25] + kernel[1][4] ~^ image[7][26] + kernel[2][0] ~^ image[8][22] + kernel[2][1] ~^ image[8][23] + kernel[2][2] ~^ image[8][24] + kernel[2][3] ~^ image[8][25] + kernel[2][4] ~^ image[8][26] + kernel[3][0] ~^ image[9][22] + kernel[3][1] ~^ image[9][23] + kernel[3][2] ~^ image[9][24] + kernel[3][3] ~^ image[9][25] + kernel[3][4] ~^ image[9][26] + kernel[4][0] ~^ image[10][22] + kernel[4][1] ~^ image[10][23] + kernel[4][2] ~^ image[10][24] + kernel[4][3] ~^ image[10][25] + kernel[4][4] ~^ image[10][26];
assign xor_sum[6][23] = kernel[0][0] ~^ image[6][23] + kernel[0][1] ~^ image[6][24] + kernel[0][2] ~^ image[6][25] + kernel[0][3] ~^ image[6][26] + kernel[0][4] ~^ image[6][27] + kernel[1][0] ~^ image[7][23] + kernel[1][1] ~^ image[7][24] + kernel[1][2] ~^ image[7][25] + kernel[1][3] ~^ image[7][26] + kernel[1][4] ~^ image[7][27] + kernel[2][0] ~^ image[8][23] + kernel[2][1] ~^ image[8][24] + kernel[2][2] ~^ image[8][25] + kernel[2][3] ~^ image[8][26] + kernel[2][4] ~^ image[8][27] + kernel[3][0] ~^ image[9][23] + kernel[3][1] ~^ image[9][24] + kernel[3][2] ~^ image[9][25] + kernel[3][3] ~^ image[9][26] + kernel[3][4] ~^ image[9][27] + kernel[4][0] ~^ image[10][23] + kernel[4][1] ~^ image[10][24] + kernel[4][2] ~^ image[10][25] + kernel[4][3] ~^ image[10][26] + kernel[4][4] ~^ image[10][27];
assign xor_sum[7][0] = kernel[0][0] ~^ image[7][0] + kernel[0][1] ~^ image[7][1] + kernel[0][2] ~^ image[7][2] + kernel[0][3] ~^ image[7][3] + kernel[0][4] ~^ image[7][4] + kernel[1][0] ~^ image[8][0] + kernel[1][1] ~^ image[8][1] + kernel[1][2] ~^ image[8][2] + kernel[1][3] ~^ image[8][3] + kernel[1][4] ~^ image[8][4] + kernel[2][0] ~^ image[9][0] + kernel[2][1] ~^ image[9][1] + kernel[2][2] ~^ image[9][2] + kernel[2][3] ~^ image[9][3] + kernel[2][4] ~^ image[9][4] + kernel[3][0] ~^ image[10][0] + kernel[3][1] ~^ image[10][1] + kernel[3][2] ~^ image[10][2] + kernel[3][3] ~^ image[10][3] + kernel[3][4] ~^ image[10][4] + kernel[4][0] ~^ image[11][0] + kernel[4][1] ~^ image[11][1] + kernel[4][2] ~^ image[11][2] + kernel[4][3] ~^ image[11][3] + kernel[4][4] ~^ image[11][4];
assign xor_sum[7][1] = kernel[0][0] ~^ image[7][1] + kernel[0][1] ~^ image[7][2] + kernel[0][2] ~^ image[7][3] + kernel[0][3] ~^ image[7][4] + kernel[0][4] ~^ image[7][5] + kernel[1][0] ~^ image[8][1] + kernel[1][1] ~^ image[8][2] + kernel[1][2] ~^ image[8][3] + kernel[1][3] ~^ image[8][4] + kernel[1][4] ~^ image[8][5] + kernel[2][0] ~^ image[9][1] + kernel[2][1] ~^ image[9][2] + kernel[2][2] ~^ image[9][3] + kernel[2][3] ~^ image[9][4] + kernel[2][4] ~^ image[9][5] + kernel[3][0] ~^ image[10][1] + kernel[3][1] ~^ image[10][2] + kernel[3][2] ~^ image[10][3] + kernel[3][3] ~^ image[10][4] + kernel[3][4] ~^ image[10][5] + kernel[4][0] ~^ image[11][1] + kernel[4][1] ~^ image[11][2] + kernel[4][2] ~^ image[11][3] + kernel[4][3] ~^ image[11][4] + kernel[4][4] ~^ image[11][5];
assign xor_sum[7][2] = kernel[0][0] ~^ image[7][2] + kernel[0][1] ~^ image[7][3] + kernel[0][2] ~^ image[7][4] + kernel[0][3] ~^ image[7][5] + kernel[0][4] ~^ image[7][6] + kernel[1][0] ~^ image[8][2] + kernel[1][1] ~^ image[8][3] + kernel[1][2] ~^ image[8][4] + kernel[1][3] ~^ image[8][5] + kernel[1][4] ~^ image[8][6] + kernel[2][0] ~^ image[9][2] + kernel[2][1] ~^ image[9][3] + kernel[2][2] ~^ image[9][4] + kernel[2][3] ~^ image[9][5] + kernel[2][4] ~^ image[9][6] + kernel[3][0] ~^ image[10][2] + kernel[3][1] ~^ image[10][3] + kernel[3][2] ~^ image[10][4] + kernel[3][3] ~^ image[10][5] + kernel[3][4] ~^ image[10][6] + kernel[4][0] ~^ image[11][2] + kernel[4][1] ~^ image[11][3] + kernel[4][2] ~^ image[11][4] + kernel[4][3] ~^ image[11][5] + kernel[4][4] ~^ image[11][6];
assign xor_sum[7][3] = kernel[0][0] ~^ image[7][3] + kernel[0][1] ~^ image[7][4] + kernel[0][2] ~^ image[7][5] + kernel[0][3] ~^ image[7][6] + kernel[0][4] ~^ image[7][7] + kernel[1][0] ~^ image[8][3] + kernel[1][1] ~^ image[8][4] + kernel[1][2] ~^ image[8][5] + kernel[1][3] ~^ image[8][6] + kernel[1][4] ~^ image[8][7] + kernel[2][0] ~^ image[9][3] + kernel[2][1] ~^ image[9][4] + kernel[2][2] ~^ image[9][5] + kernel[2][3] ~^ image[9][6] + kernel[2][4] ~^ image[9][7] + kernel[3][0] ~^ image[10][3] + kernel[3][1] ~^ image[10][4] + kernel[3][2] ~^ image[10][5] + kernel[3][3] ~^ image[10][6] + kernel[3][4] ~^ image[10][7] + kernel[4][0] ~^ image[11][3] + kernel[4][1] ~^ image[11][4] + kernel[4][2] ~^ image[11][5] + kernel[4][3] ~^ image[11][6] + kernel[4][4] ~^ image[11][7];
assign xor_sum[7][4] = kernel[0][0] ~^ image[7][4] + kernel[0][1] ~^ image[7][5] + kernel[0][2] ~^ image[7][6] + kernel[0][3] ~^ image[7][7] + kernel[0][4] ~^ image[7][8] + kernel[1][0] ~^ image[8][4] + kernel[1][1] ~^ image[8][5] + kernel[1][2] ~^ image[8][6] + kernel[1][3] ~^ image[8][7] + kernel[1][4] ~^ image[8][8] + kernel[2][0] ~^ image[9][4] + kernel[2][1] ~^ image[9][5] + kernel[2][2] ~^ image[9][6] + kernel[2][3] ~^ image[9][7] + kernel[2][4] ~^ image[9][8] + kernel[3][0] ~^ image[10][4] + kernel[3][1] ~^ image[10][5] + kernel[3][2] ~^ image[10][6] + kernel[3][3] ~^ image[10][7] + kernel[3][4] ~^ image[10][8] + kernel[4][0] ~^ image[11][4] + kernel[4][1] ~^ image[11][5] + kernel[4][2] ~^ image[11][6] + kernel[4][3] ~^ image[11][7] + kernel[4][4] ~^ image[11][8];
assign xor_sum[7][5] = kernel[0][0] ~^ image[7][5] + kernel[0][1] ~^ image[7][6] + kernel[0][2] ~^ image[7][7] + kernel[0][3] ~^ image[7][8] + kernel[0][4] ~^ image[7][9] + kernel[1][0] ~^ image[8][5] + kernel[1][1] ~^ image[8][6] + kernel[1][2] ~^ image[8][7] + kernel[1][3] ~^ image[8][8] + kernel[1][4] ~^ image[8][9] + kernel[2][0] ~^ image[9][5] + kernel[2][1] ~^ image[9][6] + kernel[2][2] ~^ image[9][7] + kernel[2][3] ~^ image[9][8] + kernel[2][4] ~^ image[9][9] + kernel[3][0] ~^ image[10][5] + kernel[3][1] ~^ image[10][6] + kernel[3][2] ~^ image[10][7] + kernel[3][3] ~^ image[10][8] + kernel[3][4] ~^ image[10][9] + kernel[4][0] ~^ image[11][5] + kernel[4][1] ~^ image[11][6] + kernel[4][2] ~^ image[11][7] + kernel[4][3] ~^ image[11][8] + kernel[4][4] ~^ image[11][9];
assign xor_sum[7][6] = kernel[0][0] ~^ image[7][6] + kernel[0][1] ~^ image[7][7] + kernel[0][2] ~^ image[7][8] + kernel[0][3] ~^ image[7][9] + kernel[0][4] ~^ image[7][10] + kernel[1][0] ~^ image[8][6] + kernel[1][1] ~^ image[8][7] + kernel[1][2] ~^ image[8][8] + kernel[1][3] ~^ image[8][9] + kernel[1][4] ~^ image[8][10] + kernel[2][0] ~^ image[9][6] + kernel[2][1] ~^ image[9][7] + kernel[2][2] ~^ image[9][8] + kernel[2][3] ~^ image[9][9] + kernel[2][4] ~^ image[9][10] + kernel[3][0] ~^ image[10][6] + kernel[3][1] ~^ image[10][7] + kernel[3][2] ~^ image[10][8] + kernel[3][3] ~^ image[10][9] + kernel[3][4] ~^ image[10][10] + kernel[4][0] ~^ image[11][6] + kernel[4][1] ~^ image[11][7] + kernel[4][2] ~^ image[11][8] + kernel[4][3] ~^ image[11][9] + kernel[4][4] ~^ image[11][10];
assign xor_sum[7][7] = kernel[0][0] ~^ image[7][7] + kernel[0][1] ~^ image[7][8] + kernel[0][2] ~^ image[7][9] + kernel[0][3] ~^ image[7][10] + kernel[0][4] ~^ image[7][11] + kernel[1][0] ~^ image[8][7] + kernel[1][1] ~^ image[8][8] + kernel[1][2] ~^ image[8][9] + kernel[1][3] ~^ image[8][10] + kernel[1][4] ~^ image[8][11] + kernel[2][0] ~^ image[9][7] + kernel[2][1] ~^ image[9][8] + kernel[2][2] ~^ image[9][9] + kernel[2][3] ~^ image[9][10] + kernel[2][4] ~^ image[9][11] + kernel[3][0] ~^ image[10][7] + kernel[3][1] ~^ image[10][8] + kernel[3][2] ~^ image[10][9] + kernel[3][3] ~^ image[10][10] + kernel[3][4] ~^ image[10][11] + kernel[4][0] ~^ image[11][7] + kernel[4][1] ~^ image[11][8] + kernel[4][2] ~^ image[11][9] + kernel[4][3] ~^ image[11][10] + kernel[4][4] ~^ image[11][11];
assign xor_sum[7][8] = kernel[0][0] ~^ image[7][8] + kernel[0][1] ~^ image[7][9] + kernel[0][2] ~^ image[7][10] + kernel[0][3] ~^ image[7][11] + kernel[0][4] ~^ image[7][12] + kernel[1][0] ~^ image[8][8] + kernel[1][1] ~^ image[8][9] + kernel[1][2] ~^ image[8][10] + kernel[1][3] ~^ image[8][11] + kernel[1][4] ~^ image[8][12] + kernel[2][0] ~^ image[9][8] + kernel[2][1] ~^ image[9][9] + kernel[2][2] ~^ image[9][10] + kernel[2][3] ~^ image[9][11] + kernel[2][4] ~^ image[9][12] + kernel[3][0] ~^ image[10][8] + kernel[3][1] ~^ image[10][9] + kernel[3][2] ~^ image[10][10] + kernel[3][3] ~^ image[10][11] + kernel[3][4] ~^ image[10][12] + kernel[4][0] ~^ image[11][8] + kernel[4][1] ~^ image[11][9] + kernel[4][2] ~^ image[11][10] + kernel[4][3] ~^ image[11][11] + kernel[4][4] ~^ image[11][12];
assign xor_sum[7][9] = kernel[0][0] ~^ image[7][9] + kernel[0][1] ~^ image[7][10] + kernel[0][2] ~^ image[7][11] + kernel[0][3] ~^ image[7][12] + kernel[0][4] ~^ image[7][13] + kernel[1][0] ~^ image[8][9] + kernel[1][1] ~^ image[8][10] + kernel[1][2] ~^ image[8][11] + kernel[1][3] ~^ image[8][12] + kernel[1][4] ~^ image[8][13] + kernel[2][0] ~^ image[9][9] + kernel[2][1] ~^ image[9][10] + kernel[2][2] ~^ image[9][11] + kernel[2][3] ~^ image[9][12] + kernel[2][4] ~^ image[9][13] + kernel[3][0] ~^ image[10][9] + kernel[3][1] ~^ image[10][10] + kernel[3][2] ~^ image[10][11] + kernel[3][3] ~^ image[10][12] + kernel[3][4] ~^ image[10][13] + kernel[4][0] ~^ image[11][9] + kernel[4][1] ~^ image[11][10] + kernel[4][2] ~^ image[11][11] + kernel[4][3] ~^ image[11][12] + kernel[4][4] ~^ image[11][13];
assign xor_sum[7][10] = kernel[0][0] ~^ image[7][10] + kernel[0][1] ~^ image[7][11] + kernel[0][2] ~^ image[7][12] + kernel[0][3] ~^ image[7][13] + kernel[0][4] ~^ image[7][14] + kernel[1][0] ~^ image[8][10] + kernel[1][1] ~^ image[8][11] + kernel[1][2] ~^ image[8][12] + kernel[1][3] ~^ image[8][13] + kernel[1][4] ~^ image[8][14] + kernel[2][0] ~^ image[9][10] + kernel[2][1] ~^ image[9][11] + kernel[2][2] ~^ image[9][12] + kernel[2][3] ~^ image[9][13] + kernel[2][4] ~^ image[9][14] + kernel[3][0] ~^ image[10][10] + kernel[3][1] ~^ image[10][11] + kernel[3][2] ~^ image[10][12] + kernel[3][3] ~^ image[10][13] + kernel[3][4] ~^ image[10][14] + kernel[4][0] ~^ image[11][10] + kernel[4][1] ~^ image[11][11] + kernel[4][2] ~^ image[11][12] + kernel[4][3] ~^ image[11][13] + kernel[4][4] ~^ image[11][14];
assign xor_sum[7][11] = kernel[0][0] ~^ image[7][11] + kernel[0][1] ~^ image[7][12] + kernel[0][2] ~^ image[7][13] + kernel[0][3] ~^ image[7][14] + kernel[0][4] ~^ image[7][15] + kernel[1][0] ~^ image[8][11] + kernel[1][1] ~^ image[8][12] + kernel[1][2] ~^ image[8][13] + kernel[1][3] ~^ image[8][14] + kernel[1][4] ~^ image[8][15] + kernel[2][0] ~^ image[9][11] + kernel[2][1] ~^ image[9][12] + kernel[2][2] ~^ image[9][13] + kernel[2][3] ~^ image[9][14] + kernel[2][4] ~^ image[9][15] + kernel[3][0] ~^ image[10][11] + kernel[3][1] ~^ image[10][12] + kernel[3][2] ~^ image[10][13] + kernel[3][3] ~^ image[10][14] + kernel[3][4] ~^ image[10][15] + kernel[4][0] ~^ image[11][11] + kernel[4][1] ~^ image[11][12] + kernel[4][2] ~^ image[11][13] + kernel[4][3] ~^ image[11][14] + kernel[4][4] ~^ image[11][15];
assign xor_sum[7][12] = kernel[0][0] ~^ image[7][12] + kernel[0][1] ~^ image[7][13] + kernel[0][2] ~^ image[7][14] + kernel[0][3] ~^ image[7][15] + kernel[0][4] ~^ image[7][16] + kernel[1][0] ~^ image[8][12] + kernel[1][1] ~^ image[8][13] + kernel[1][2] ~^ image[8][14] + kernel[1][3] ~^ image[8][15] + kernel[1][4] ~^ image[8][16] + kernel[2][0] ~^ image[9][12] + kernel[2][1] ~^ image[9][13] + kernel[2][2] ~^ image[9][14] + kernel[2][3] ~^ image[9][15] + kernel[2][4] ~^ image[9][16] + kernel[3][0] ~^ image[10][12] + kernel[3][1] ~^ image[10][13] + kernel[3][2] ~^ image[10][14] + kernel[3][3] ~^ image[10][15] + kernel[3][4] ~^ image[10][16] + kernel[4][0] ~^ image[11][12] + kernel[4][1] ~^ image[11][13] + kernel[4][2] ~^ image[11][14] + kernel[4][3] ~^ image[11][15] + kernel[4][4] ~^ image[11][16];
assign xor_sum[7][13] = kernel[0][0] ~^ image[7][13] + kernel[0][1] ~^ image[7][14] + kernel[0][2] ~^ image[7][15] + kernel[0][3] ~^ image[7][16] + kernel[0][4] ~^ image[7][17] + kernel[1][0] ~^ image[8][13] + kernel[1][1] ~^ image[8][14] + kernel[1][2] ~^ image[8][15] + kernel[1][3] ~^ image[8][16] + kernel[1][4] ~^ image[8][17] + kernel[2][0] ~^ image[9][13] + kernel[2][1] ~^ image[9][14] + kernel[2][2] ~^ image[9][15] + kernel[2][3] ~^ image[9][16] + kernel[2][4] ~^ image[9][17] + kernel[3][0] ~^ image[10][13] + kernel[3][1] ~^ image[10][14] + kernel[3][2] ~^ image[10][15] + kernel[3][3] ~^ image[10][16] + kernel[3][4] ~^ image[10][17] + kernel[4][0] ~^ image[11][13] + kernel[4][1] ~^ image[11][14] + kernel[4][2] ~^ image[11][15] + kernel[4][3] ~^ image[11][16] + kernel[4][4] ~^ image[11][17];
assign xor_sum[7][14] = kernel[0][0] ~^ image[7][14] + kernel[0][1] ~^ image[7][15] + kernel[0][2] ~^ image[7][16] + kernel[0][3] ~^ image[7][17] + kernel[0][4] ~^ image[7][18] + kernel[1][0] ~^ image[8][14] + kernel[1][1] ~^ image[8][15] + kernel[1][2] ~^ image[8][16] + kernel[1][3] ~^ image[8][17] + kernel[1][4] ~^ image[8][18] + kernel[2][0] ~^ image[9][14] + kernel[2][1] ~^ image[9][15] + kernel[2][2] ~^ image[9][16] + kernel[2][3] ~^ image[9][17] + kernel[2][4] ~^ image[9][18] + kernel[3][0] ~^ image[10][14] + kernel[3][1] ~^ image[10][15] + kernel[3][2] ~^ image[10][16] + kernel[3][3] ~^ image[10][17] + kernel[3][4] ~^ image[10][18] + kernel[4][0] ~^ image[11][14] + kernel[4][1] ~^ image[11][15] + kernel[4][2] ~^ image[11][16] + kernel[4][3] ~^ image[11][17] + kernel[4][4] ~^ image[11][18];
assign xor_sum[7][15] = kernel[0][0] ~^ image[7][15] + kernel[0][1] ~^ image[7][16] + kernel[0][2] ~^ image[7][17] + kernel[0][3] ~^ image[7][18] + kernel[0][4] ~^ image[7][19] + kernel[1][0] ~^ image[8][15] + kernel[1][1] ~^ image[8][16] + kernel[1][2] ~^ image[8][17] + kernel[1][3] ~^ image[8][18] + kernel[1][4] ~^ image[8][19] + kernel[2][0] ~^ image[9][15] + kernel[2][1] ~^ image[9][16] + kernel[2][2] ~^ image[9][17] + kernel[2][3] ~^ image[9][18] + kernel[2][4] ~^ image[9][19] + kernel[3][0] ~^ image[10][15] + kernel[3][1] ~^ image[10][16] + kernel[3][2] ~^ image[10][17] + kernel[3][3] ~^ image[10][18] + kernel[3][4] ~^ image[10][19] + kernel[4][0] ~^ image[11][15] + kernel[4][1] ~^ image[11][16] + kernel[4][2] ~^ image[11][17] + kernel[4][3] ~^ image[11][18] + kernel[4][4] ~^ image[11][19];
assign xor_sum[7][16] = kernel[0][0] ~^ image[7][16] + kernel[0][1] ~^ image[7][17] + kernel[0][2] ~^ image[7][18] + kernel[0][3] ~^ image[7][19] + kernel[0][4] ~^ image[7][20] + kernel[1][0] ~^ image[8][16] + kernel[1][1] ~^ image[8][17] + kernel[1][2] ~^ image[8][18] + kernel[1][3] ~^ image[8][19] + kernel[1][4] ~^ image[8][20] + kernel[2][0] ~^ image[9][16] + kernel[2][1] ~^ image[9][17] + kernel[2][2] ~^ image[9][18] + kernel[2][3] ~^ image[9][19] + kernel[2][4] ~^ image[9][20] + kernel[3][0] ~^ image[10][16] + kernel[3][1] ~^ image[10][17] + kernel[3][2] ~^ image[10][18] + kernel[3][3] ~^ image[10][19] + kernel[3][4] ~^ image[10][20] + kernel[4][0] ~^ image[11][16] + kernel[4][1] ~^ image[11][17] + kernel[4][2] ~^ image[11][18] + kernel[4][3] ~^ image[11][19] + kernel[4][4] ~^ image[11][20];
assign xor_sum[7][17] = kernel[0][0] ~^ image[7][17] + kernel[0][1] ~^ image[7][18] + kernel[0][2] ~^ image[7][19] + kernel[0][3] ~^ image[7][20] + kernel[0][4] ~^ image[7][21] + kernel[1][0] ~^ image[8][17] + kernel[1][1] ~^ image[8][18] + kernel[1][2] ~^ image[8][19] + kernel[1][3] ~^ image[8][20] + kernel[1][4] ~^ image[8][21] + kernel[2][0] ~^ image[9][17] + kernel[2][1] ~^ image[9][18] + kernel[2][2] ~^ image[9][19] + kernel[2][3] ~^ image[9][20] + kernel[2][4] ~^ image[9][21] + kernel[3][0] ~^ image[10][17] + kernel[3][1] ~^ image[10][18] + kernel[3][2] ~^ image[10][19] + kernel[3][3] ~^ image[10][20] + kernel[3][4] ~^ image[10][21] + kernel[4][0] ~^ image[11][17] + kernel[4][1] ~^ image[11][18] + kernel[4][2] ~^ image[11][19] + kernel[4][3] ~^ image[11][20] + kernel[4][4] ~^ image[11][21];
assign xor_sum[7][18] = kernel[0][0] ~^ image[7][18] + kernel[0][1] ~^ image[7][19] + kernel[0][2] ~^ image[7][20] + kernel[0][3] ~^ image[7][21] + kernel[0][4] ~^ image[7][22] + kernel[1][0] ~^ image[8][18] + kernel[1][1] ~^ image[8][19] + kernel[1][2] ~^ image[8][20] + kernel[1][3] ~^ image[8][21] + kernel[1][4] ~^ image[8][22] + kernel[2][0] ~^ image[9][18] + kernel[2][1] ~^ image[9][19] + kernel[2][2] ~^ image[9][20] + kernel[2][3] ~^ image[9][21] + kernel[2][4] ~^ image[9][22] + kernel[3][0] ~^ image[10][18] + kernel[3][1] ~^ image[10][19] + kernel[3][2] ~^ image[10][20] + kernel[3][3] ~^ image[10][21] + kernel[3][4] ~^ image[10][22] + kernel[4][0] ~^ image[11][18] + kernel[4][1] ~^ image[11][19] + kernel[4][2] ~^ image[11][20] + kernel[4][3] ~^ image[11][21] + kernel[4][4] ~^ image[11][22];
assign xor_sum[7][19] = kernel[0][0] ~^ image[7][19] + kernel[0][1] ~^ image[7][20] + kernel[0][2] ~^ image[7][21] + kernel[0][3] ~^ image[7][22] + kernel[0][4] ~^ image[7][23] + kernel[1][0] ~^ image[8][19] + kernel[1][1] ~^ image[8][20] + kernel[1][2] ~^ image[8][21] + kernel[1][3] ~^ image[8][22] + kernel[1][4] ~^ image[8][23] + kernel[2][0] ~^ image[9][19] + kernel[2][1] ~^ image[9][20] + kernel[2][2] ~^ image[9][21] + kernel[2][3] ~^ image[9][22] + kernel[2][4] ~^ image[9][23] + kernel[3][0] ~^ image[10][19] + kernel[3][1] ~^ image[10][20] + kernel[3][2] ~^ image[10][21] + kernel[3][3] ~^ image[10][22] + kernel[3][4] ~^ image[10][23] + kernel[4][0] ~^ image[11][19] + kernel[4][1] ~^ image[11][20] + kernel[4][2] ~^ image[11][21] + kernel[4][3] ~^ image[11][22] + kernel[4][4] ~^ image[11][23];
assign xor_sum[7][20] = kernel[0][0] ~^ image[7][20] + kernel[0][1] ~^ image[7][21] + kernel[0][2] ~^ image[7][22] + kernel[0][3] ~^ image[7][23] + kernel[0][4] ~^ image[7][24] + kernel[1][0] ~^ image[8][20] + kernel[1][1] ~^ image[8][21] + kernel[1][2] ~^ image[8][22] + kernel[1][3] ~^ image[8][23] + kernel[1][4] ~^ image[8][24] + kernel[2][0] ~^ image[9][20] + kernel[2][1] ~^ image[9][21] + kernel[2][2] ~^ image[9][22] + kernel[2][3] ~^ image[9][23] + kernel[2][4] ~^ image[9][24] + kernel[3][0] ~^ image[10][20] + kernel[3][1] ~^ image[10][21] + kernel[3][2] ~^ image[10][22] + kernel[3][3] ~^ image[10][23] + kernel[3][4] ~^ image[10][24] + kernel[4][0] ~^ image[11][20] + kernel[4][1] ~^ image[11][21] + kernel[4][2] ~^ image[11][22] + kernel[4][3] ~^ image[11][23] + kernel[4][4] ~^ image[11][24];
assign xor_sum[7][21] = kernel[0][0] ~^ image[7][21] + kernel[0][1] ~^ image[7][22] + kernel[0][2] ~^ image[7][23] + kernel[0][3] ~^ image[7][24] + kernel[0][4] ~^ image[7][25] + kernel[1][0] ~^ image[8][21] + kernel[1][1] ~^ image[8][22] + kernel[1][2] ~^ image[8][23] + kernel[1][3] ~^ image[8][24] + kernel[1][4] ~^ image[8][25] + kernel[2][0] ~^ image[9][21] + kernel[2][1] ~^ image[9][22] + kernel[2][2] ~^ image[9][23] + kernel[2][3] ~^ image[9][24] + kernel[2][4] ~^ image[9][25] + kernel[3][0] ~^ image[10][21] + kernel[3][1] ~^ image[10][22] + kernel[3][2] ~^ image[10][23] + kernel[3][3] ~^ image[10][24] + kernel[3][4] ~^ image[10][25] + kernel[4][0] ~^ image[11][21] + kernel[4][1] ~^ image[11][22] + kernel[4][2] ~^ image[11][23] + kernel[4][3] ~^ image[11][24] + kernel[4][4] ~^ image[11][25];
assign xor_sum[7][22] = kernel[0][0] ~^ image[7][22] + kernel[0][1] ~^ image[7][23] + kernel[0][2] ~^ image[7][24] + kernel[0][3] ~^ image[7][25] + kernel[0][4] ~^ image[7][26] + kernel[1][0] ~^ image[8][22] + kernel[1][1] ~^ image[8][23] + kernel[1][2] ~^ image[8][24] + kernel[1][3] ~^ image[8][25] + kernel[1][4] ~^ image[8][26] + kernel[2][0] ~^ image[9][22] + kernel[2][1] ~^ image[9][23] + kernel[2][2] ~^ image[9][24] + kernel[2][3] ~^ image[9][25] + kernel[2][4] ~^ image[9][26] + kernel[3][0] ~^ image[10][22] + kernel[3][1] ~^ image[10][23] + kernel[3][2] ~^ image[10][24] + kernel[3][3] ~^ image[10][25] + kernel[3][4] ~^ image[10][26] + kernel[4][0] ~^ image[11][22] + kernel[4][1] ~^ image[11][23] + kernel[4][2] ~^ image[11][24] + kernel[4][3] ~^ image[11][25] + kernel[4][4] ~^ image[11][26];
assign xor_sum[7][23] = kernel[0][0] ~^ image[7][23] + kernel[0][1] ~^ image[7][24] + kernel[0][2] ~^ image[7][25] + kernel[0][3] ~^ image[7][26] + kernel[0][4] ~^ image[7][27] + kernel[1][0] ~^ image[8][23] + kernel[1][1] ~^ image[8][24] + kernel[1][2] ~^ image[8][25] + kernel[1][3] ~^ image[8][26] + kernel[1][4] ~^ image[8][27] + kernel[2][0] ~^ image[9][23] + kernel[2][1] ~^ image[9][24] + kernel[2][2] ~^ image[9][25] + kernel[2][3] ~^ image[9][26] + kernel[2][4] ~^ image[9][27] + kernel[3][0] ~^ image[10][23] + kernel[3][1] ~^ image[10][24] + kernel[3][2] ~^ image[10][25] + kernel[3][3] ~^ image[10][26] + kernel[3][4] ~^ image[10][27] + kernel[4][0] ~^ image[11][23] + kernel[4][1] ~^ image[11][24] + kernel[4][2] ~^ image[11][25] + kernel[4][3] ~^ image[11][26] + kernel[4][4] ~^ image[11][27];
assign xor_sum[8][0] = kernel[0][0] ~^ image[8][0] + kernel[0][1] ~^ image[8][1] + kernel[0][2] ~^ image[8][2] + kernel[0][3] ~^ image[8][3] + kernel[0][4] ~^ image[8][4] + kernel[1][0] ~^ image[9][0] + kernel[1][1] ~^ image[9][1] + kernel[1][2] ~^ image[9][2] + kernel[1][3] ~^ image[9][3] + kernel[1][4] ~^ image[9][4] + kernel[2][0] ~^ image[10][0] + kernel[2][1] ~^ image[10][1] + kernel[2][2] ~^ image[10][2] + kernel[2][3] ~^ image[10][3] + kernel[2][4] ~^ image[10][4] + kernel[3][0] ~^ image[11][0] + kernel[3][1] ~^ image[11][1] + kernel[3][2] ~^ image[11][2] + kernel[3][3] ~^ image[11][3] + kernel[3][4] ~^ image[11][4] + kernel[4][0] ~^ image[12][0] + kernel[4][1] ~^ image[12][1] + kernel[4][2] ~^ image[12][2] + kernel[4][3] ~^ image[12][3] + kernel[4][4] ~^ image[12][4];
assign xor_sum[8][1] = kernel[0][0] ~^ image[8][1] + kernel[0][1] ~^ image[8][2] + kernel[0][2] ~^ image[8][3] + kernel[0][3] ~^ image[8][4] + kernel[0][4] ~^ image[8][5] + kernel[1][0] ~^ image[9][1] + kernel[1][1] ~^ image[9][2] + kernel[1][2] ~^ image[9][3] + kernel[1][3] ~^ image[9][4] + kernel[1][4] ~^ image[9][5] + kernel[2][0] ~^ image[10][1] + kernel[2][1] ~^ image[10][2] + kernel[2][2] ~^ image[10][3] + kernel[2][3] ~^ image[10][4] + kernel[2][4] ~^ image[10][5] + kernel[3][0] ~^ image[11][1] + kernel[3][1] ~^ image[11][2] + kernel[3][2] ~^ image[11][3] + kernel[3][3] ~^ image[11][4] + kernel[3][4] ~^ image[11][5] + kernel[4][0] ~^ image[12][1] + kernel[4][1] ~^ image[12][2] + kernel[4][2] ~^ image[12][3] + kernel[4][3] ~^ image[12][4] + kernel[4][4] ~^ image[12][5];
assign xor_sum[8][2] = kernel[0][0] ~^ image[8][2] + kernel[0][1] ~^ image[8][3] + kernel[0][2] ~^ image[8][4] + kernel[0][3] ~^ image[8][5] + kernel[0][4] ~^ image[8][6] + kernel[1][0] ~^ image[9][2] + kernel[1][1] ~^ image[9][3] + kernel[1][2] ~^ image[9][4] + kernel[1][3] ~^ image[9][5] + kernel[1][4] ~^ image[9][6] + kernel[2][0] ~^ image[10][2] + kernel[2][1] ~^ image[10][3] + kernel[2][2] ~^ image[10][4] + kernel[2][3] ~^ image[10][5] + kernel[2][4] ~^ image[10][6] + kernel[3][0] ~^ image[11][2] + kernel[3][1] ~^ image[11][3] + kernel[3][2] ~^ image[11][4] + kernel[3][3] ~^ image[11][5] + kernel[3][4] ~^ image[11][6] + kernel[4][0] ~^ image[12][2] + kernel[4][1] ~^ image[12][3] + kernel[4][2] ~^ image[12][4] + kernel[4][3] ~^ image[12][5] + kernel[4][4] ~^ image[12][6];
assign xor_sum[8][3] = kernel[0][0] ~^ image[8][3] + kernel[0][1] ~^ image[8][4] + kernel[0][2] ~^ image[8][5] + kernel[0][3] ~^ image[8][6] + kernel[0][4] ~^ image[8][7] + kernel[1][0] ~^ image[9][3] + kernel[1][1] ~^ image[9][4] + kernel[1][2] ~^ image[9][5] + kernel[1][3] ~^ image[9][6] + kernel[1][4] ~^ image[9][7] + kernel[2][0] ~^ image[10][3] + kernel[2][1] ~^ image[10][4] + kernel[2][2] ~^ image[10][5] + kernel[2][3] ~^ image[10][6] + kernel[2][4] ~^ image[10][7] + kernel[3][0] ~^ image[11][3] + kernel[3][1] ~^ image[11][4] + kernel[3][2] ~^ image[11][5] + kernel[3][3] ~^ image[11][6] + kernel[3][4] ~^ image[11][7] + kernel[4][0] ~^ image[12][3] + kernel[4][1] ~^ image[12][4] + kernel[4][2] ~^ image[12][5] + kernel[4][3] ~^ image[12][6] + kernel[4][4] ~^ image[12][7];
assign xor_sum[8][4] = kernel[0][0] ~^ image[8][4] + kernel[0][1] ~^ image[8][5] + kernel[0][2] ~^ image[8][6] + kernel[0][3] ~^ image[8][7] + kernel[0][4] ~^ image[8][8] + kernel[1][0] ~^ image[9][4] + kernel[1][1] ~^ image[9][5] + kernel[1][2] ~^ image[9][6] + kernel[1][3] ~^ image[9][7] + kernel[1][4] ~^ image[9][8] + kernel[2][0] ~^ image[10][4] + kernel[2][1] ~^ image[10][5] + kernel[2][2] ~^ image[10][6] + kernel[2][3] ~^ image[10][7] + kernel[2][4] ~^ image[10][8] + kernel[3][0] ~^ image[11][4] + kernel[3][1] ~^ image[11][5] + kernel[3][2] ~^ image[11][6] + kernel[3][3] ~^ image[11][7] + kernel[3][4] ~^ image[11][8] + kernel[4][0] ~^ image[12][4] + kernel[4][1] ~^ image[12][5] + kernel[4][2] ~^ image[12][6] + kernel[4][3] ~^ image[12][7] + kernel[4][4] ~^ image[12][8];
assign xor_sum[8][5] = kernel[0][0] ~^ image[8][5] + kernel[0][1] ~^ image[8][6] + kernel[0][2] ~^ image[8][7] + kernel[0][3] ~^ image[8][8] + kernel[0][4] ~^ image[8][9] + kernel[1][0] ~^ image[9][5] + kernel[1][1] ~^ image[9][6] + kernel[1][2] ~^ image[9][7] + kernel[1][3] ~^ image[9][8] + kernel[1][4] ~^ image[9][9] + kernel[2][0] ~^ image[10][5] + kernel[2][1] ~^ image[10][6] + kernel[2][2] ~^ image[10][7] + kernel[2][3] ~^ image[10][8] + kernel[2][4] ~^ image[10][9] + kernel[3][0] ~^ image[11][5] + kernel[3][1] ~^ image[11][6] + kernel[3][2] ~^ image[11][7] + kernel[3][3] ~^ image[11][8] + kernel[3][4] ~^ image[11][9] + kernel[4][0] ~^ image[12][5] + kernel[4][1] ~^ image[12][6] + kernel[4][2] ~^ image[12][7] + kernel[4][3] ~^ image[12][8] + kernel[4][4] ~^ image[12][9];
assign xor_sum[8][6] = kernel[0][0] ~^ image[8][6] + kernel[0][1] ~^ image[8][7] + kernel[0][2] ~^ image[8][8] + kernel[0][3] ~^ image[8][9] + kernel[0][4] ~^ image[8][10] + kernel[1][0] ~^ image[9][6] + kernel[1][1] ~^ image[9][7] + kernel[1][2] ~^ image[9][8] + kernel[1][3] ~^ image[9][9] + kernel[1][4] ~^ image[9][10] + kernel[2][0] ~^ image[10][6] + kernel[2][1] ~^ image[10][7] + kernel[2][2] ~^ image[10][8] + kernel[2][3] ~^ image[10][9] + kernel[2][4] ~^ image[10][10] + kernel[3][0] ~^ image[11][6] + kernel[3][1] ~^ image[11][7] + kernel[3][2] ~^ image[11][8] + kernel[3][3] ~^ image[11][9] + kernel[3][4] ~^ image[11][10] + kernel[4][0] ~^ image[12][6] + kernel[4][1] ~^ image[12][7] + kernel[4][2] ~^ image[12][8] + kernel[4][3] ~^ image[12][9] + kernel[4][4] ~^ image[12][10];
assign xor_sum[8][7] = kernel[0][0] ~^ image[8][7] + kernel[0][1] ~^ image[8][8] + kernel[0][2] ~^ image[8][9] + kernel[0][3] ~^ image[8][10] + kernel[0][4] ~^ image[8][11] + kernel[1][0] ~^ image[9][7] + kernel[1][1] ~^ image[9][8] + kernel[1][2] ~^ image[9][9] + kernel[1][3] ~^ image[9][10] + kernel[1][4] ~^ image[9][11] + kernel[2][0] ~^ image[10][7] + kernel[2][1] ~^ image[10][8] + kernel[2][2] ~^ image[10][9] + kernel[2][3] ~^ image[10][10] + kernel[2][4] ~^ image[10][11] + kernel[3][0] ~^ image[11][7] + kernel[3][1] ~^ image[11][8] + kernel[3][2] ~^ image[11][9] + kernel[3][3] ~^ image[11][10] + kernel[3][4] ~^ image[11][11] + kernel[4][0] ~^ image[12][7] + kernel[4][1] ~^ image[12][8] + kernel[4][2] ~^ image[12][9] + kernel[4][3] ~^ image[12][10] + kernel[4][4] ~^ image[12][11];
assign xor_sum[8][8] = kernel[0][0] ~^ image[8][8] + kernel[0][1] ~^ image[8][9] + kernel[0][2] ~^ image[8][10] + kernel[0][3] ~^ image[8][11] + kernel[0][4] ~^ image[8][12] + kernel[1][0] ~^ image[9][8] + kernel[1][1] ~^ image[9][9] + kernel[1][2] ~^ image[9][10] + kernel[1][3] ~^ image[9][11] + kernel[1][4] ~^ image[9][12] + kernel[2][0] ~^ image[10][8] + kernel[2][1] ~^ image[10][9] + kernel[2][2] ~^ image[10][10] + kernel[2][3] ~^ image[10][11] + kernel[2][4] ~^ image[10][12] + kernel[3][0] ~^ image[11][8] + kernel[3][1] ~^ image[11][9] + kernel[3][2] ~^ image[11][10] + kernel[3][3] ~^ image[11][11] + kernel[3][4] ~^ image[11][12] + kernel[4][0] ~^ image[12][8] + kernel[4][1] ~^ image[12][9] + kernel[4][2] ~^ image[12][10] + kernel[4][3] ~^ image[12][11] + kernel[4][4] ~^ image[12][12];
assign xor_sum[8][9] = kernel[0][0] ~^ image[8][9] + kernel[0][1] ~^ image[8][10] + kernel[0][2] ~^ image[8][11] + kernel[0][3] ~^ image[8][12] + kernel[0][4] ~^ image[8][13] + kernel[1][0] ~^ image[9][9] + kernel[1][1] ~^ image[9][10] + kernel[1][2] ~^ image[9][11] + kernel[1][3] ~^ image[9][12] + kernel[1][4] ~^ image[9][13] + kernel[2][0] ~^ image[10][9] + kernel[2][1] ~^ image[10][10] + kernel[2][2] ~^ image[10][11] + kernel[2][3] ~^ image[10][12] + kernel[2][4] ~^ image[10][13] + kernel[3][0] ~^ image[11][9] + kernel[3][1] ~^ image[11][10] + kernel[3][2] ~^ image[11][11] + kernel[3][3] ~^ image[11][12] + kernel[3][4] ~^ image[11][13] + kernel[4][0] ~^ image[12][9] + kernel[4][1] ~^ image[12][10] + kernel[4][2] ~^ image[12][11] + kernel[4][3] ~^ image[12][12] + kernel[4][4] ~^ image[12][13];
assign xor_sum[8][10] = kernel[0][0] ~^ image[8][10] + kernel[0][1] ~^ image[8][11] + kernel[0][2] ~^ image[8][12] + kernel[0][3] ~^ image[8][13] + kernel[0][4] ~^ image[8][14] + kernel[1][0] ~^ image[9][10] + kernel[1][1] ~^ image[9][11] + kernel[1][2] ~^ image[9][12] + kernel[1][3] ~^ image[9][13] + kernel[1][4] ~^ image[9][14] + kernel[2][0] ~^ image[10][10] + kernel[2][1] ~^ image[10][11] + kernel[2][2] ~^ image[10][12] + kernel[2][3] ~^ image[10][13] + kernel[2][4] ~^ image[10][14] + kernel[3][0] ~^ image[11][10] + kernel[3][1] ~^ image[11][11] + kernel[3][2] ~^ image[11][12] + kernel[3][3] ~^ image[11][13] + kernel[3][4] ~^ image[11][14] + kernel[4][0] ~^ image[12][10] + kernel[4][1] ~^ image[12][11] + kernel[4][2] ~^ image[12][12] + kernel[4][3] ~^ image[12][13] + kernel[4][4] ~^ image[12][14];
assign xor_sum[8][11] = kernel[0][0] ~^ image[8][11] + kernel[0][1] ~^ image[8][12] + kernel[0][2] ~^ image[8][13] + kernel[0][3] ~^ image[8][14] + kernel[0][4] ~^ image[8][15] + kernel[1][0] ~^ image[9][11] + kernel[1][1] ~^ image[9][12] + kernel[1][2] ~^ image[9][13] + kernel[1][3] ~^ image[9][14] + kernel[1][4] ~^ image[9][15] + kernel[2][0] ~^ image[10][11] + kernel[2][1] ~^ image[10][12] + kernel[2][2] ~^ image[10][13] + kernel[2][3] ~^ image[10][14] + kernel[2][4] ~^ image[10][15] + kernel[3][0] ~^ image[11][11] + kernel[3][1] ~^ image[11][12] + kernel[3][2] ~^ image[11][13] + kernel[3][3] ~^ image[11][14] + kernel[3][4] ~^ image[11][15] + kernel[4][0] ~^ image[12][11] + kernel[4][1] ~^ image[12][12] + kernel[4][2] ~^ image[12][13] + kernel[4][3] ~^ image[12][14] + kernel[4][4] ~^ image[12][15];
assign xor_sum[8][12] = kernel[0][0] ~^ image[8][12] + kernel[0][1] ~^ image[8][13] + kernel[0][2] ~^ image[8][14] + kernel[0][3] ~^ image[8][15] + kernel[0][4] ~^ image[8][16] + kernel[1][0] ~^ image[9][12] + kernel[1][1] ~^ image[9][13] + kernel[1][2] ~^ image[9][14] + kernel[1][3] ~^ image[9][15] + kernel[1][4] ~^ image[9][16] + kernel[2][0] ~^ image[10][12] + kernel[2][1] ~^ image[10][13] + kernel[2][2] ~^ image[10][14] + kernel[2][3] ~^ image[10][15] + kernel[2][4] ~^ image[10][16] + kernel[3][0] ~^ image[11][12] + kernel[3][1] ~^ image[11][13] + kernel[3][2] ~^ image[11][14] + kernel[3][3] ~^ image[11][15] + kernel[3][4] ~^ image[11][16] + kernel[4][0] ~^ image[12][12] + kernel[4][1] ~^ image[12][13] + kernel[4][2] ~^ image[12][14] + kernel[4][3] ~^ image[12][15] + kernel[4][4] ~^ image[12][16];
assign xor_sum[8][13] = kernel[0][0] ~^ image[8][13] + kernel[0][1] ~^ image[8][14] + kernel[0][2] ~^ image[8][15] + kernel[0][3] ~^ image[8][16] + kernel[0][4] ~^ image[8][17] + kernel[1][0] ~^ image[9][13] + kernel[1][1] ~^ image[9][14] + kernel[1][2] ~^ image[9][15] + kernel[1][3] ~^ image[9][16] + kernel[1][4] ~^ image[9][17] + kernel[2][0] ~^ image[10][13] + kernel[2][1] ~^ image[10][14] + kernel[2][2] ~^ image[10][15] + kernel[2][3] ~^ image[10][16] + kernel[2][4] ~^ image[10][17] + kernel[3][0] ~^ image[11][13] + kernel[3][1] ~^ image[11][14] + kernel[3][2] ~^ image[11][15] + kernel[3][3] ~^ image[11][16] + kernel[3][4] ~^ image[11][17] + kernel[4][0] ~^ image[12][13] + kernel[4][1] ~^ image[12][14] + kernel[4][2] ~^ image[12][15] + kernel[4][3] ~^ image[12][16] + kernel[4][4] ~^ image[12][17];
assign xor_sum[8][14] = kernel[0][0] ~^ image[8][14] + kernel[0][1] ~^ image[8][15] + kernel[0][2] ~^ image[8][16] + kernel[0][3] ~^ image[8][17] + kernel[0][4] ~^ image[8][18] + kernel[1][0] ~^ image[9][14] + kernel[1][1] ~^ image[9][15] + kernel[1][2] ~^ image[9][16] + kernel[1][3] ~^ image[9][17] + kernel[1][4] ~^ image[9][18] + kernel[2][0] ~^ image[10][14] + kernel[2][1] ~^ image[10][15] + kernel[2][2] ~^ image[10][16] + kernel[2][3] ~^ image[10][17] + kernel[2][4] ~^ image[10][18] + kernel[3][0] ~^ image[11][14] + kernel[3][1] ~^ image[11][15] + kernel[3][2] ~^ image[11][16] + kernel[3][3] ~^ image[11][17] + kernel[3][4] ~^ image[11][18] + kernel[4][0] ~^ image[12][14] + kernel[4][1] ~^ image[12][15] + kernel[4][2] ~^ image[12][16] + kernel[4][3] ~^ image[12][17] + kernel[4][4] ~^ image[12][18];
assign xor_sum[8][15] = kernel[0][0] ~^ image[8][15] + kernel[0][1] ~^ image[8][16] + kernel[0][2] ~^ image[8][17] + kernel[0][3] ~^ image[8][18] + kernel[0][4] ~^ image[8][19] + kernel[1][0] ~^ image[9][15] + kernel[1][1] ~^ image[9][16] + kernel[1][2] ~^ image[9][17] + kernel[1][3] ~^ image[9][18] + kernel[1][4] ~^ image[9][19] + kernel[2][0] ~^ image[10][15] + kernel[2][1] ~^ image[10][16] + kernel[2][2] ~^ image[10][17] + kernel[2][3] ~^ image[10][18] + kernel[2][4] ~^ image[10][19] + kernel[3][0] ~^ image[11][15] + kernel[3][1] ~^ image[11][16] + kernel[3][2] ~^ image[11][17] + kernel[3][3] ~^ image[11][18] + kernel[3][4] ~^ image[11][19] + kernel[4][0] ~^ image[12][15] + kernel[4][1] ~^ image[12][16] + kernel[4][2] ~^ image[12][17] + kernel[4][3] ~^ image[12][18] + kernel[4][4] ~^ image[12][19];
assign xor_sum[8][16] = kernel[0][0] ~^ image[8][16] + kernel[0][1] ~^ image[8][17] + kernel[0][2] ~^ image[8][18] + kernel[0][3] ~^ image[8][19] + kernel[0][4] ~^ image[8][20] + kernel[1][0] ~^ image[9][16] + kernel[1][1] ~^ image[9][17] + kernel[1][2] ~^ image[9][18] + kernel[1][3] ~^ image[9][19] + kernel[1][4] ~^ image[9][20] + kernel[2][0] ~^ image[10][16] + kernel[2][1] ~^ image[10][17] + kernel[2][2] ~^ image[10][18] + kernel[2][3] ~^ image[10][19] + kernel[2][4] ~^ image[10][20] + kernel[3][0] ~^ image[11][16] + kernel[3][1] ~^ image[11][17] + kernel[3][2] ~^ image[11][18] + kernel[3][3] ~^ image[11][19] + kernel[3][4] ~^ image[11][20] + kernel[4][0] ~^ image[12][16] + kernel[4][1] ~^ image[12][17] + kernel[4][2] ~^ image[12][18] + kernel[4][3] ~^ image[12][19] + kernel[4][4] ~^ image[12][20];
assign xor_sum[8][17] = kernel[0][0] ~^ image[8][17] + kernel[0][1] ~^ image[8][18] + kernel[0][2] ~^ image[8][19] + kernel[0][3] ~^ image[8][20] + kernel[0][4] ~^ image[8][21] + kernel[1][0] ~^ image[9][17] + kernel[1][1] ~^ image[9][18] + kernel[1][2] ~^ image[9][19] + kernel[1][3] ~^ image[9][20] + kernel[1][4] ~^ image[9][21] + kernel[2][0] ~^ image[10][17] + kernel[2][1] ~^ image[10][18] + kernel[2][2] ~^ image[10][19] + kernel[2][3] ~^ image[10][20] + kernel[2][4] ~^ image[10][21] + kernel[3][0] ~^ image[11][17] + kernel[3][1] ~^ image[11][18] + kernel[3][2] ~^ image[11][19] + kernel[3][3] ~^ image[11][20] + kernel[3][4] ~^ image[11][21] + kernel[4][0] ~^ image[12][17] + kernel[4][1] ~^ image[12][18] + kernel[4][2] ~^ image[12][19] + kernel[4][3] ~^ image[12][20] + kernel[4][4] ~^ image[12][21];
assign xor_sum[8][18] = kernel[0][0] ~^ image[8][18] + kernel[0][1] ~^ image[8][19] + kernel[0][2] ~^ image[8][20] + kernel[0][3] ~^ image[8][21] + kernel[0][4] ~^ image[8][22] + kernel[1][0] ~^ image[9][18] + kernel[1][1] ~^ image[9][19] + kernel[1][2] ~^ image[9][20] + kernel[1][3] ~^ image[9][21] + kernel[1][4] ~^ image[9][22] + kernel[2][0] ~^ image[10][18] + kernel[2][1] ~^ image[10][19] + kernel[2][2] ~^ image[10][20] + kernel[2][3] ~^ image[10][21] + kernel[2][4] ~^ image[10][22] + kernel[3][0] ~^ image[11][18] + kernel[3][1] ~^ image[11][19] + kernel[3][2] ~^ image[11][20] + kernel[3][3] ~^ image[11][21] + kernel[3][4] ~^ image[11][22] + kernel[4][0] ~^ image[12][18] + kernel[4][1] ~^ image[12][19] + kernel[4][2] ~^ image[12][20] + kernel[4][3] ~^ image[12][21] + kernel[4][4] ~^ image[12][22];
assign xor_sum[8][19] = kernel[0][0] ~^ image[8][19] + kernel[0][1] ~^ image[8][20] + kernel[0][2] ~^ image[8][21] + kernel[0][3] ~^ image[8][22] + kernel[0][4] ~^ image[8][23] + kernel[1][0] ~^ image[9][19] + kernel[1][1] ~^ image[9][20] + kernel[1][2] ~^ image[9][21] + kernel[1][3] ~^ image[9][22] + kernel[1][4] ~^ image[9][23] + kernel[2][0] ~^ image[10][19] + kernel[2][1] ~^ image[10][20] + kernel[2][2] ~^ image[10][21] + kernel[2][3] ~^ image[10][22] + kernel[2][4] ~^ image[10][23] + kernel[3][0] ~^ image[11][19] + kernel[3][1] ~^ image[11][20] + kernel[3][2] ~^ image[11][21] + kernel[3][3] ~^ image[11][22] + kernel[3][4] ~^ image[11][23] + kernel[4][0] ~^ image[12][19] + kernel[4][1] ~^ image[12][20] + kernel[4][2] ~^ image[12][21] + kernel[4][3] ~^ image[12][22] + kernel[4][4] ~^ image[12][23];
assign xor_sum[8][20] = kernel[0][0] ~^ image[8][20] + kernel[0][1] ~^ image[8][21] + kernel[0][2] ~^ image[8][22] + kernel[0][3] ~^ image[8][23] + kernel[0][4] ~^ image[8][24] + kernel[1][0] ~^ image[9][20] + kernel[1][1] ~^ image[9][21] + kernel[1][2] ~^ image[9][22] + kernel[1][3] ~^ image[9][23] + kernel[1][4] ~^ image[9][24] + kernel[2][0] ~^ image[10][20] + kernel[2][1] ~^ image[10][21] + kernel[2][2] ~^ image[10][22] + kernel[2][3] ~^ image[10][23] + kernel[2][4] ~^ image[10][24] + kernel[3][0] ~^ image[11][20] + kernel[3][1] ~^ image[11][21] + kernel[3][2] ~^ image[11][22] + kernel[3][3] ~^ image[11][23] + kernel[3][4] ~^ image[11][24] + kernel[4][0] ~^ image[12][20] + kernel[4][1] ~^ image[12][21] + kernel[4][2] ~^ image[12][22] + kernel[4][3] ~^ image[12][23] + kernel[4][4] ~^ image[12][24];
assign xor_sum[8][21] = kernel[0][0] ~^ image[8][21] + kernel[0][1] ~^ image[8][22] + kernel[0][2] ~^ image[8][23] + kernel[0][3] ~^ image[8][24] + kernel[0][4] ~^ image[8][25] + kernel[1][0] ~^ image[9][21] + kernel[1][1] ~^ image[9][22] + kernel[1][2] ~^ image[9][23] + kernel[1][3] ~^ image[9][24] + kernel[1][4] ~^ image[9][25] + kernel[2][0] ~^ image[10][21] + kernel[2][1] ~^ image[10][22] + kernel[2][2] ~^ image[10][23] + kernel[2][3] ~^ image[10][24] + kernel[2][4] ~^ image[10][25] + kernel[3][0] ~^ image[11][21] + kernel[3][1] ~^ image[11][22] + kernel[3][2] ~^ image[11][23] + kernel[3][3] ~^ image[11][24] + kernel[3][4] ~^ image[11][25] + kernel[4][0] ~^ image[12][21] + kernel[4][1] ~^ image[12][22] + kernel[4][2] ~^ image[12][23] + kernel[4][3] ~^ image[12][24] + kernel[4][4] ~^ image[12][25];
assign xor_sum[8][22] = kernel[0][0] ~^ image[8][22] + kernel[0][1] ~^ image[8][23] + kernel[0][2] ~^ image[8][24] + kernel[0][3] ~^ image[8][25] + kernel[0][4] ~^ image[8][26] + kernel[1][0] ~^ image[9][22] + kernel[1][1] ~^ image[9][23] + kernel[1][2] ~^ image[9][24] + kernel[1][3] ~^ image[9][25] + kernel[1][4] ~^ image[9][26] + kernel[2][0] ~^ image[10][22] + kernel[2][1] ~^ image[10][23] + kernel[2][2] ~^ image[10][24] + kernel[2][3] ~^ image[10][25] + kernel[2][4] ~^ image[10][26] + kernel[3][0] ~^ image[11][22] + kernel[3][1] ~^ image[11][23] + kernel[3][2] ~^ image[11][24] + kernel[3][3] ~^ image[11][25] + kernel[3][4] ~^ image[11][26] + kernel[4][0] ~^ image[12][22] + kernel[4][1] ~^ image[12][23] + kernel[4][2] ~^ image[12][24] + kernel[4][3] ~^ image[12][25] + kernel[4][4] ~^ image[12][26];
assign xor_sum[8][23] = kernel[0][0] ~^ image[8][23] + kernel[0][1] ~^ image[8][24] + kernel[0][2] ~^ image[8][25] + kernel[0][3] ~^ image[8][26] + kernel[0][4] ~^ image[8][27] + kernel[1][0] ~^ image[9][23] + kernel[1][1] ~^ image[9][24] + kernel[1][2] ~^ image[9][25] + kernel[1][3] ~^ image[9][26] + kernel[1][4] ~^ image[9][27] + kernel[2][0] ~^ image[10][23] + kernel[2][1] ~^ image[10][24] + kernel[2][2] ~^ image[10][25] + kernel[2][3] ~^ image[10][26] + kernel[2][4] ~^ image[10][27] + kernel[3][0] ~^ image[11][23] + kernel[3][1] ~^ image[11][24] + kernel[3][2] ~^ image[11][25] + kernel[3][3] ~^ image[11][26] + kernel[3][4] ~^ image[11][27] + kernel[4][0] ~^ image[12][23] + kernel[4][1] ~^ image[12][24] + kernel[4][2] ~^ image[12][25] + kernel[4][3] ~^ image[12][26] + kernel[4][4] ~^ image[12][27];
assign xor_sum[9][0] = kernel[0][0] ~^ image[9][0] + kernel[0][1] ~^ image[9][1] + kernel[0][2] ~^ image[9][2] + kernel[0][3] ~^ image[9][3] + kernel[0][4] ~^ image[9][4] + kernel[1][0] ~^ image[10][0] + kernel[1][1] ~^ image[10][1] + kernel[1][2] ~^ image[10][2] + kernel[1][3] ~^ image[10][3] + kernel[1][4] ~^ image[10][4] + kernel[2][0] ~^ image[11][0] + kernel[2][1] ~^ image[11][1] + kernel[2][2] ~^ image[11][2] + kernel[2][3] ~^ image[11][3] + kernel[2][4] ~^ image[11][4] + kernel[3][0] ~^ image[12][0] + kernel[3][1] ~^ image[12][1] + kernel[3][2] ~^ image[12][2] + kernel[3][3] ~^ image[12][3] + kernel[3][4] ~^ image[12][4] + kernel[4][0] ~^ image[13][0] + kernel[4][1] ~^ image[13][1] + kernel[4][2] ~^ image[13][2] + kernel[4][3] ~^ image[13][3] + kernel[4][4] ~^ image[13][4];
assign xor_sum[9][1] = kernel[0][0] ~^ image[9][1] + kernel[0][1] ~^ image[9][2] + kernel[0][2] ~^ image[9][3] + kernel[0][3] ~^ image[9][4] + kernel[0][4] ~^ image[9][5] + kernel[1][0] ~^ image[10][1] + kernel[1][1] ~^ image[10][2] + kernel[1][2] ~^ image[10][3] + kernel[1][3] ~^ image[10][4] + kernel[1][4] ~^ image[10][5] + kernel[2][0] ~^ image[11][1] + kernel[2][1] ~^ image[11][2] + kernel[2][2] ~^ image[11][3] + kernel[2][3] ~^ image[11][4] + kernel[2][4] ~^ image[11][5] + kernel[3][0] ~^ image[12][1] + kernel[3][1] ~^ image[12][2] + kernel[3][2] ~^ image[12][3] + kernel[3][3] ~^ image[12][4] + kernel[3][4] ~^ image[12][5] + kernel[4][0] ~^ image[13][1] + kernel[4][1] ~^ image[13][2] + kernel[4][2] ~^ image[13][3] + kernel[4][3] ~^ image[13][4] + kernel[4][4] ~^ image[13][5];
assign xor_sum[9][2] = kernel[0][0] ~^ image[9][2] + kernel[0][1] ~^ image[9][3] + kernel[0][2] ~^ image[9][4] + kernel[0][3] ~^ image[9][5] + kernel[0][4] ~^ image[9][6] + kernel[1][0] ~^ image[10][2] + kernel[1][1] ~^ image[10][3] + kernel[1][2] ~^ image[10][4] + kernel[1][3] ~^ image[10][5] + kernel[1][4] ~^ image[10][6] + kernel[2][0] ~^ image[11][2] + kernel[2][1] ~^ image[11][3] + kernel[2][2] ~^ image[11][4] + kernel[2][3] ~^ image[11][5] + kernel[2][4] ~^ image[11][6] + kernel[3][0] ~^ image[12][2] + kernel[3][1] ~^ image[12][3] + kernel[3][2] ~^ image[12][4] + kernel[3][3] ~^ image[12][5] + kernel[3][4] ~^ image[12][6] + kernel[4][0] ~^ image[13][2] + kernel[4][1] ~^ image[13][3] + kernel[4][2] ~^ image[13][4] + kernel[4][3] ~^ image[13][5] + kernel[4][4] ~^ image[13][6];
assign xor_sum[9][3] = kernel[0][0] ~^ image[9][3] + kernel[0][1] ~^ image[9][4] + kernel[0][2] ~^ image[9][5] + kernel[0][3] ~^ image[9][6] + kernel[0][4] ~^ image[9][7] + kernel[1][0] ~^ image[10][3] + kernel[1][1] ~^ image[10][4] + kernel[1][2] ~^ image[10][5] + kernel[1][3] ~^ image[10][6] + kernel[1][4] ~^ image[10][7] + kernel[2][0] ~^ image[11][3] + kernel[2][1] ~^ image[11][4] + kernel[2][2] ~^ image[11][5] + kernel[2][3] ~^ image[11][6] + kernel[2][4] ~^ image[11][7] + kernel[3][0] ~^ image[12][3] + kernel[3][1] ~^ image[12][4] + kernel[3][2] ~^ image[12][5] + kernel[3][3] ~^ image[12][6] + kernel[3][4] ~^ image[12][7] + kernel[4][0] ~^ image[13][3] + kernel[4][1] ~^ image[13][4] + kernel[4][2] ~^ image[13][5] + kernel[4][3] ~^ image[13][6] + kernel[4][4] ~^ image[13][7];
assign xor_sum[9][4] = kernel[0][0] ~^ image[9][4] + kernel[0][1] ~^ image[9][5] + kernel[0][2] ~^ image[9][6] + kernel[0][3] ~^ image[9][7] + kernel[0][4] ~^ image[9][8] + kernel[1][0] ~^ image[10][4] + kernel[1][1] ~^ image[10][5] + kernel[1][2] ~^ image[10][6] + kernel[1][3] ~^ image[10][7] + kernel[1][4] ~^ image[10][8] + kernel[2][0] ~^ image[11][4] + kernel[2][1] ~^ image[11][5] + kernel[2][2] ~^ image[11][6] + kernel[2][3] ~^ image[11][7] + kernel[2][4] ~^ image[11][8] + kernel[3][0] ~^ image[12][4] + kernel[3][1] ~^ image[12][5] + kernel[3][2] ~^ image[12][6] + kernel[3][3] ~^ image[12][7] + kernel[3][4] ~^ image[12][8] + kernel[4][0] ~^ image[13][4] + kernel[4][1] ~^ image[13][5] + kernel[4][2] ~^ image[13][6] + kernel[4][3] ~^ image[13][7] + kernel[4][4] ~^ image[13][8];
assign xor_sum[9][5] = kernel[0][0] ~^ image[9][5] + kernel[0][1] ~^ image[9][6] + kernel[0][2] ~^ image[9][7] + kernel[0][3] ~^ image[9][8] + kernel[0][4] ~^ image[9][9] + kernel[1][0] ~^ image[10][5] + kernel[1][1] ~^ image[10][6] + kernel[1][2] ~^ image[10][7] + kernel[1][3] ~^ image[10][8] + kernel[1][4] ~^ image[10][9] + kernel[2][0] ~^ image[11][5] + kernel[2][1] ~^ image[11][6] + kernel[2][2] ~^ image[11][7] + kernel[2][3] ~^ image[11][8] + kernel[2][4] ~^ image[11][9] + kernel[3][0] ~^ image[12][5] + kernel[3][1] ~^ image[12][6] + kernel[3][2] ~^ image[12][7] + kernel[3][3] ~^ image[12][8] + kernel[3][4] ~^ image[12][9] + kernel[4][0] ~^ image[13][5] + kernel[4][1] ~^ image[13][6] + kernel[4][2] ~^ image[13][7] + kernel[4][3] ~^ image[13][8] + kernel[4][4] ~^ image[13][9];
assign xor_sum[9][6] = kernel[0][0] ~^ image[9][6] + kernel[0][1] ~^ image[9][7] + kernel[0][2] ~^ image[9][8] + kernel[0][3] ~^ image[9][9] + kernel[0][4] ~^ image[9][10] + kernel[1][0] ~^ image[10][6] + kernel[1][1] ~^ image[10][7] + kernel[1][2] ~^ image[10][8] + kernel[1][3] ~^ image[10][9] + kernel[1][4] ~^ image[10][10] + kernel[2][0] ~^ image[11][6] + kernel[2][1] ~^ image[11][7] + kernel[2][2] ~^ image[11][8] + kernel[2][3] ~^ image[11][9] + kernel[2][4] ~^ image[11][10] + kernel[3][0] ~^ image[12][6] + kernel[3][1] ~^ image[12][7] + kernel[3][2] ~^ image[12][8] + kernel[3][3] ~^ image[12][9] + kernel[3][4] ~^ image[12][10] + kernel[4][0] ~^ image[13][6] + kernel[4][1] ~^ image[13][7] + kernel[4][2] ~^ image[13][8] + kernel[4][3] ~^ image[13][9] + kernel[4][4] ~^ image[13][10];
assign xor_sum[9][7] = kernel[0][0] ~^ image[9][7] + kernel[0][1] ~^ image[9][8] + kernel[0][2] ~^ image[9][9] + kernel[0][3] ~^ image[9][10] + kernel[0][4] ~^ image[9][11] + kernel[1][0] ~^ image[10][7] + kernel[1][1] ~^ image[10][8] + kernel[1][2] ~^ image[10][9] + kernel[1][3] ~^ image[10][10] + kernel[1][4] ~^ image[10][11] + kernel[2][0] ~^ image[11][7] + kernel[2][1] ~^ image[11][8] + kernel[2][2] ~^ image[11][9] + kernel[2][3] ~^ image[11][10] + kernel[2][4] ~^ image[11][11] + kernel[3][0] ~^ image[12][7] + kernel[3][1] ~^ image[12][8] + kernel[3][2] ~^ image[12][9] + kernel[3][3] ~^ image[12][10] + kernel[3][4] ~^ image[12][11] + kernel[4][0] ~^ image[13][7] + kernel[4][1] ~^ image[13][8] + kernel[4][2] ~^ image[13][9] + kernel[4][3] ~^ image[13][10] + kernel[4][4] ~^ image[13][11];
assign xor_sum[9][8] = kernel[0][0] ~^ image[9][8] + kernel[0][1] ~^ image[9][9] + kernel[0][2] ~^ image[9][10] + kernel[0][3] ~^ image[9][11] + kernel[0][4] ~^ image[9][12] + kernel[1][0] ~^ image[10][8] + kernel[1][1] ~^ image[10][9] + kernel[1][2] ~^ image[10][10] + kernel[1][3] ~^ image[10][11] + kernel[1][4] ~^ image[10][12] + kernel[2][0] ~^ image[11][8] + kernel[2][1] ~^ image[11][9] + kernel[2][2] ~^ image[11][10] + kernel[2][3] ~^ image[11][11] + kernel[2][4] ~^ image[11][12] + kernel[3][0] ~^ image[12][8] + kernel[3][1] ~^ image[12][9] + kernel[3][2] ~^ image[12][10] + kernel[3][3] ~^ image[12][11] + kernel[3][4] ~^ image[12][12] + kernel[4][0] ~^ image[13][8] + kernel[4][1] ~^ image[13][9] + kernel[4][2] ~^ image[13][10] + kernel[4][3] ~^ image[13][11] + kernel[4][4] ~^ image[13][12];
assign xor_sum[9][9] = kernel[0][0] ~^ image[9][9] + kernel[0][1] ~^ image[9][10] + kernel[0][2] ~^ image[9][11] + kernel[0][3] ~^ image[9][12] + kernel[0][4] ~^ image[9][13] + kernel[1][0] ~^ image[10][9] + kernel[1][1] ~^ image[10][10] + kernel[1][2] ~^ image[10][11] + kernel[1][3] ~^ image[10][12] + kernel[1][4] ~^ image[10][13] + kernel[2][0] ~^ image[11][9] + kernel[2][1] ~^ image[11][10] + kernel[2][2] ~^ image[11][11] + kernel[2][3] ~^ image[11][12] + kernel[2][4] ~^ image[11][13] + kernel[3][0] ~^ image[12][9] + kernel[3][1] ~^ image[12][10] + kernel[3][2] ~^ image[12][11] + kernel[3][3] ~^ image[12][12] + kernel[3][4] ~^ image[12][13] + kernel[4][0] ~^ image[13][9] + kernel[4][1] ~^ image[13][10] + kernel[4][2] ~^ image[13][11] + kernel[4][3] ~^ image[13][12] + kernel[4][4] ~^ image[13][13];
assign xor_sum[9][10] = kernel[0][0] ~^ image[9][10] + kernel[0][1] ~^ image[9][11] + kernel[0][2] ~^ image[9][12] + kernel[0][3] ~^ image[9][13] + kernel[0][4] ~^ image[9][14] + kernel[1][0] ~^ image[10][10] + kernel[1][1] ~^ image[10][11] + kernel[1][2] ~^ image[10][12] + kernel[1][3] ~^ image[10][13] + kernel[1][4] ~^ image[10][14] + kernel[2][0] ~^ image[11][10] + kernel[2][1] ~^ image[11][11] + kernel[2][2] ~^ image[11][12] + kernel[2][3] ~^ image[11][13] + kernel[2][4] ~^ image[11][14] + kernel[3][0] ~^ image[12][10] + kernel[3][1] ~^ image[12][11] + kernel[3][2] ~^ image[12][12] + kernel[3][3] ~^ image[12][13] + kernel[3][4] ~^ image[12][14] + kernel[4][0] ~^ image[13][10] + kernel[4][1] ~^ image[13][11] + kernel[4][2] ~^ image[13][12] + kernel[4][3] ~^ image[13][13] + kernel[4][4] ~^ image[13][14];
assign xor_sum[9][11] = kernel[0][0] ~^ image[9][11] + kernel[0][1] ~^ image[9][12] + kernel[0][2] ~^ image[9][13] + kernel[0][3] ~^ image[9][14] + kernel[0][4] ~^ image[9][15] + kernel[1][0] ~^ image[10][11] + kernel[1][1] ~^ image[10][12] + kernel[1][2] ~^ image[10][13] + kernel[1][3] ~^ image[10][14] + kernel[1][4] ~^ image[10][15] + kernel[2][0] ~^ image[11][11] + kernel[2][1] ~^ image[11][12] + kernel[2][2] ~^ image[11][13] + kernel[2][3] ~^ image[11][14] + kernel[2][4] ~^ image[11][15] + kernel[3][0] ~^ image[12][11] + kernel[3][1] ~^ image[12][12] + kernel[3][2] ~^ image[12][13] + kernel[3][3] ~^ image[12][14] + kernel[3][4] ~^ image[12][15] + kernel[4][0] ~^ image[13][11] + kernel[4][1] ~^ image[13][12] + kernel[4][2] ~^ image[13][13] + kernel[4][3] ~^ image[13][14] + kernel[4][4] ~^ image[13][15];
assign xor_sum[9][12] = kernel[0][0] ~^ image[9][12] + kernel[0][1] ~^ image[9][13] + kernel[0][2] ~^ image[9][14] + kernel[0][3] ~^ image[9][15] + kernel[0][4] ~^ image[9][16] + kernel[1][0] ~^ image[10][12] + kernel[1][1] ~^ image[10][13] + kernel[1][2] ~^ image[10][14] + kernel[1][3] ~^ image[10][15] + kernel[1][4] ~^ image[10][16] + kernel[2][0] ~^ image[11][12] + kernel[2][1] ~^ image[11][13] + kernel[2][2] ~^ image[11][14] + kernel[2][3] ~^ image[11][15] + kernel[2][4] ~^ image[11][16] + kernel[3][0] ~^ image[12][12] + kernel[3][1] ~^ image[12][13] + kernel[3][2] ~^ image[12][14] + kernel[3][3] ~^ image[12][15] + kernel[3][4] ~^ image[12][16] + kernel[4][0] ~^ image[13][12] + kernel[4][1] ~^ image[13][13] + kernel[4][2] ~^ image[13][14] + kernel[4][3] ~^ image[13][15] + kernel[4][4] ~^ image[13][16];
assign xor_sum[9][13] = kernel[0][0] ~^ image[9][13] + kernel[0][1] ~^ image[9][14] + kernel[0][2] ~^ image[9][15] + kernel[0][3] ~^ image[9][16] + kernel[0][4] ~^ image[9][17] + kernel[1][0] ~^ image[10][13] + kernel[1][1] ~^ image[10][14] + kernel[1][2] ~^ image[10][15] + kernel[1][3] ~^ image[10][16] + kernel[1][4] ~^ image[10][17] + kernel[2][0] ~^ image[11][13] + kernel[2][1] ~^ image[11][14] + kernel[2][2] ~^ image[11][15] + kernel[2][3] ~^ image[11][16] + kernel[2][4] ~^ image[11][17] + kernel[3][0] ~^ image[12][13] + kernel[3][1] ~^ image[12][14] + kernel[3][2] ~^ image[12][15] + kernel[3][3] ~^ image[12][16] + kernel[3][4] ~^ image[12][17] + kernel[4][0] ~^ image[13][13] + kernel[4][1] ~^ image[13][14] + kernel[4][2] ~^ image[13][15] + kernel[4][3] ~^ image[13][16] + kernel[4][4] ~^ image[13][17];
assign xor_sum[9][14] = kernel[0][0] ~^ image[9][14] + kernel[0][1] ~^ image[9][15] + kernel[0][2] ~^ image[9][16] + kernel[0][3] ~^ image[9][17] + kernel[0][4] ~^ image[9][18] + kernel[1][0] ~^ image[10][14] + kernel[1][1] ~^ image[10][15] + kernel[1][2] ~^ image[10][16] + kernel[1][3] ~^ image[10][17] + kernel[1][4] ~^ image[10][18] + kernel[2][0] ~^ image[11][14] + kernel[2][1] ~^ image[11][15] + kernel[2][2] ~^ image[11][16] + kernel[2][3] ~^ image[11][17] + kernel[2][4] ~^ image[11][18] + kernel[3][0] ~^ image[12][14] + kernel[3][1] ~^ image[12][15] + kernel[3][2] ~^ image[12][16] + kernel[3][3] ~^ image[12][17] + kernel[3][4] ~^ image[12][18] + kernel[4][0] ~^ image[13][14] + kernel[4][1] ~^ image[13][15] + kernel[4][2] ~^ image[13][16] + kernel[4][3] ~^ image[13][17] + kernel[4][4] ~^ image[13][18];
assign xor_sum[9][15] = kernel[0][0] ~^ image[9][15] + kernel[0][1] ~^ image[9][16] + kernel[0][2] ~^ image[9][17] + kernel[0][3] ~^ image[9][18] + kernel[0][4] ~^ image[9][19] + kernel[1][0] ~^ image[10][15] + kernel[1][1] ~^ image[10][16] + kernel[1][2] ~^ image[10][17] + kernel[1][3] ~^ image[10][18] + kernel[1][4] ~^ image[10][19] + kernel[2][0] ~^ image[11][15] + kernel[2][1] ~^ image[11][16] + kernel[2][2] ~^ image[11][17] + kernel[2][3] ~^ image[11][18] + kernel[2][4] ~^ image[11][19] + kernel[3][0] ~^ image[12][15] + kernel[3][1] ~^ image[12][16] + kernel[3][2] ~^ image[12][17] + kernel[3][3] ~^ image[12][18] + kernel[3][4] ~^ image[12][19] + kernel[4][0] ~^ image[13][15] + kernel[4][1] ~^ image[13][16] + kernel[4][2] ~^ image[13][17] + kernel[4][3] ~^ image[13][18] + kernel[4][4] ~^ image[13][19];
assign xor_sum[9][16] = kernel[0][0] ~^ image[9][16] + kernel[0][1] ~^ image[9][17] + kernel[0][2] ~^ image[9][18] + kernel[0][3] ~^ image[9][19] + kernel[0][4] ~^ image[9][20] + kernel[1][0] ~^ image[10][16] + kernel[1][1] ~^ image[10][17] + kernel[1][2] ~^ image[10][18] + kernel[1][3] ~^ image[10][19] + kernel[1][4] ~^ image[10][20] + kernel[2][0] ~^ image[11][16] + kernel[2][1] ~^ image[11][17] + kernel[2][2] ~^ image[11][18] + kernel[2][3] ~^ image[11][19] + kernel[2][4] ~^ image[11][20] + kernel[3][0] ~^ image[12][16] + kernel[3][1] ~^ image[12][17] + kernel[3][2] ~^ image[12][18] + kernel[3][3] ~^ image[12][19] + kernel[3][4] ~^ image[12][20] + kernel[4][0] ~^ image[13][16] + kernel[4][1] ~^ image[13][17] + kernel[4][2] ~^ image[13][18] + kernel[4][3] ~^ image[13][19] + kernel[4][4] ~^ image[13][20];
assign xor_sum[9][17] = kernel[0][0] ~^ image[9][17] + kernel[0][1] ~^ image[9][18] + kernel[0][2] ~^ image[9][19] + kernel[0][3] ~^ image[9][20] + kernel[0][4] ~^ image[9][21] + kernel[1][0] ~^ image[10][17] + kernel[1][1] ~^ image[10][18] + kernel[1][2] ~^ image[10][19] + kernel[1][3] ~^ image[10][20] + kernel[1][4] ~^ image[10][21] + kernel[2][0] ~^ image[11][17] + kernel[2][1] ~^ image[11][18] + kernel[2][2] ~^ image[11][19] + kernel[2][3] ~^ image[11][20] + kernel[2][4] ~^ image[11][21] + kernel[3][0] ~^ image[12][17] + kernel[3][1] ~^ image[12][18] + kernel[3][2] ~^ image[12][19] + kernel[3][3] ~^ image[12][20] + kernel[3][4] ~^ image[12][21] + kernel[4][0] ~^ image[13][17] + kernel[4][1] ~^ image[13][18] + kernel[4][2] ~^ image[13][19] + kernel[4][3] ~^ image[13][20] + kernel[4][4] ~^ image[13][21];
assign xor_sum[9][18] = kernel[0][0] ~^ image[9][18] + kernel[0][1] ~^ image[9][19] + kernel[0][2] ~^ image[9][20] + kernel[0][3] ~^ image[9][21] + kernel[0][4] ~^ image[9][22] + kernel[1][0] ~^ image[10][18] + kernel[1][1] ~^ image[10][19] + kernel[1][2] ~^ image[10][20] + kernel[1][3] ~^ image[10][21] + kernel[1][4] ~^ image[10][22] + kernel[2][0] ~^ image[11][18] + kernel[2][1] ~^ image[11][19] + kernel[2][2] ~^ image[11][20] + kernel[2][3] ~^ image[11][21] + kernel[2][4] ~^ image[11][22] + kernel[3][0] ~^ image[12][18] + kernel[3][1] ~^ image[12][19] + kernel[3][2] ~^ image[12][20] + kernel[3][3] ~^ image[12][21] + kernel[3][4] ~^ image[12][22] + kernel[4][0] ~^ image[13][18] + kernel[4][1] ~^ image[13][19] + kernel[4][2] ~^ image[13][20] + kernel[4][3] ~^ image[13][21] + kernel[4][4] ~^ image[13][22];
assign xor_sum[9][19] = kernel[0][0] ~^ image[9][19] + kernel[0][1] ~^ image[9][20] + kernel[0][2] ~^ image[9][21] + kernel[0][3] ~^ image[9][22] + kernel[0][4] ~^ image[9][23] + kernel[1][0] ~^ image[10][19] + kernel[1][1] ~^ image[10][20] + kernel[1][2] ~^ image[10][21] + kernel[1][3] ~^ image[10][22] + kernel[1][4] ~^ image[10][23] + kernel[2][0] ~^ image[11][19] + kernel[2][1] ~^ image[11][20] + kernel[2][2] ~^ image[11][21] + kernel[2][3] ~^ image[11][22] + kernel[2][4] ~^ image[11][23] + kernel[3][0] ~^ image[12][19] + kernel[3][1] ~^ image[12][20] + kernel[3][2] ~^ image[12][21] + kernel[3][3] ~^ image[12][22] + kernel[3][4] ~^ image[12][23] + kernel[4][0] ~^ image[13][19] + kernel[4][1] ~^ image[13][20] + kernel[4][2] ~^ image[13][21] + kernel[4][3] ~^ image[13][22] + kernel[4][4] ~^ image[13][23];
assign xor_sum[9][20] = kernel[0][0] ~^ image[9][20] + kernel[0][1] ~^ image[9][21] + kernel[0][2] ~^ image[9][22] + kernel[0][3] ~^ image[9][23] + kernel[0][4] ~^ image[9][24] + kernel[1][0] ~^ image[10][20] + kernel[1][1] ~^ image[10][21] + kernel[1][2] ~^ image[10][22] + kernel[1][3] ~^ image[10][23] + kernel[1][4] ~^ image[10][24] + kernel[2][0] ~^ image[11][20] + kernel[2][1] ~^ image[11][21] + kernel[2][2] ~^ image[11][22] + kernel[2][3] ~^ image[11][23] + kernel[2][4] ~^ image[11][24] + kernel[3][0] ~^ image[12][20] + kernel[3][1] ~^ image[12][21] + kernel[3][2] ~^ image[12][22] + kernel[3][3] ~^ image[12][23] + kernel[3][4] ~^ image[12][24] + kernel[4][0] ~^ image[13][20] + kernel[4][1] ~^ image[13][21] + kernel[4][2] ~^ image[13][22] + kernel[4][3] ~^ image[13][23] + kernel[4][4] ~^ image[13][24];
assign xor_sum[9][21] = kernel[0][0] ~^ image[9][21] + kernel[0][1] ~^ image[9][22] + kernel[0][2] ~^ image[9][23] + kernel[0][3] ~^ image[9][24] + kernel[0][4] ~^ image[9][25] + kernel[1][0] ~^ image[10][21] + kernel[1][1] ~^ image[10][22] + kernel[1][2] ~^ image[10][23] + kernel[1][3] ~^ image[10][24] + kernel[1][4] ~^ image[10][25] + kernel[2][0] ~^ image[11][21] + kernel[2][1] ~^ image[11][22] + kernel[2][2] ~^ image[11][23] + kernel[2][3] ~^ image[11][24] + kernel[2][4] ~^ image[11][25] + kernel[3][0] ~^ image[12][21] + kernel[3][1] ~^ image[12][22] + kernel[3][2] ~^ image[12][23] + kernel[3][3] ~^ image[12][24] + kernel[3][4] ~^ image[12][25] + kernel[4][0] ~^ image[13][21] + kernel[4][1] ~^ image[13][22] + kernel[4][2] ~^ image[13][23] + kernel[4][3] ~^ image[13][24] + kernel[4][4] ~^ image[13][25];
assign xor_sum[9][22] = kernel[0][0] ~^ image[9][22] + kernel[0][1] ~^ image[9][23] + kernel[0][2] ~^ image[9][24] + kernel[0][3] ~^ image[9][25] + kernel[0][4] ~^ image[9][26] + kernel[1][0] ~^ image[10][22] + kernel[1][1] ~^ image[10][23] + kernel[1][2] ~^ image[10][24] + kernel[1][3] ~^ image[10][25] + kernel[1][4] ~^ image[10][26] + kernel[2][0] ~^ image[11][22] + kernel[2][1] ~^ image[11][23] + kernel[2][2] ~^ image[11][24] + kernel[2][3] ~^ image[11][25] + kernel[2][4] ~^ image[11][26] + kernel[3][0] ~^ image[12][22] + kernel[3][1] ~^ image[12][23] + kernel[3][2] ~^ image[12][24] + kernel[3][3] ~^ image[12][25] + kernel[3][4] ~^ image[12][26] + kernel[4][0] ~^ image[13][22] + kernel[4][1] ~^ image[13][23] + kernel[4][2] ~^ image[13][24] + kernel[4][3] ~^ image[13][25] + kernel[4][4] ~^ image[13][26];
assign xor_sum[9][23] = kernel[0][0] ~^ image[9][23] + kernel[0][1] ~^ image[9][24] + kernel[0][2] ~^ image[9][25] + kernel[0][3] ~^ image[9][26] + kernel[0][4] ~^ image[9][27] + kernel[1][0] ~^ image[10][23] + kernel[1][1] ~^ image[10][24] + kernel[1][2] ~^ image[10][25] + kernel[1][3] ~^ image[10][26] + kernel[1][4] ~^ image[10][27] + kernel[2][0] ~^ image[11][23] + kernel[2][1] ~^ image[11][24] + kernel[2][2] ~^ image[11][25] + kernel[2][3] ~^ image[11][26] + kernel[2][4] ~^ image[11][27] + kernel[3][0] ~^ image[12][23] + kernel[3][1] ~^ image[12][24] + kernel[3][2] ~^ image[12][25] + kernel[3][3] ~^ image[12][26] + kernel[3][4] ~^ image[12][27] + kernel[4][0] ~^ image[13][23] + kernel[4][1] ~^ image[13][24] + kernel[4][2] ~^ image[13][25] + kernel[4][3] ~^ image[13][26] + kernel[4][4] ~^ image[13][27];
assign xor_sum[10][0] = kernel[0][0] ~^ image[10][0] + kernel[0][1] ~^ image[10][1] + kernel[0][2] ~^ image[10][2] + kernel[0][3] ~^ image[10][3] + kernel[0][4] ~^ image[10][4] + kernel[1][0] ~^ image[11][0] + kernel[1][1] ~^ image[11][1] + kernel[1][2] ~^ image[11][2] + kernel[1][3] ~^ image[11][3] + kernel[1][4] ~^ image[11][4] + kernel[2][0] ~^ image[12][0] + kernel[2][1] ~^ image[12][1] + kernel[2][2] ~^ image[12][2] + kernel[2][3] ~^ image[12][3] + kernel[2][4] ~^ image[12][4] + kernel[3][0] ~^ image[13][0] + kernel[3][1] ~^ image[13][1] + kernel[3][2] ~^ image[13][2] + kernel[3][3] ~^ image[13][3] + kernel[3][4] ~^ image[13][4] + kernel[4][0] ~^ image[14][0] + kernel[4][1] ~^ image[14][1] + kernel[4][2] ~^ image[14][2] + kernel[4][3] ~^ image[14][3] + kernel[4][4] ~^ image[14][4];
assign xor_sum[10][1] = kernel[0][0] ~^ image[10][1] + kernel[0][1] ~^ image[10][2] + kernel[0][2] ~^ image[10][3] + kernel[0][3] ~^ image[10][4] + kernel[0][4] ~^ image[10][5] + kernel[1][0] ~^ image[11][1] + kernel[1][1] ~^ image[11][2] + kernel[1][2] ~^ image[11][3] + kernel[1][3] ~^ image[11][4] + kernel[1][4] ~^ image[11][5] + kernel[2][0] ~^ image[12][1] + kernel[2][1] ~^ image[12][2] + kernel[2][2] ~^ image[12][3] + kernel[2][3] ~^ image[12][4] + kernel[2][4] ~^ image[12][5] + kernel[3][0] ~^ image[13][1] + kernel[3][1] ~^ image[13][2] + kernel[3][2] ~^ image[13][3] + kernel[3][3] ~^ image[13][4] + kernel[3][4] ~^ image[13][5] + kernel[4][0] ~^ image[14][1] + kernel[4][1] ~^ image[14][2] + kernel[4][2] ~^ image[14][3] + kernel[4][3] ~^ image[14][4] + kernel[4][4] ~^ image[14][5];
assign xor_sum[10][2] = kernel[0][0] ~^ image[10][2] + kernel[0][1] ~^ image[10][3] + kernel[0][2] ~^ image[10][4] + kernel[0][3] ~^ image[10][5] + kernel[0][4] ~^ image[10][6] + kernel[1][0] ~^ image[11][2] + kernel[1][1] ~^ image[11][3] + kernel[1][2] ~^ image[11][4] + kernel[1][3] ~^ image[11][5] + kernel[1][4] ~^ image[11][6] + kernel[2][0] ~^ image[12][2] + kernel[2][1] ~^ image[12][3] + kernel[2][2] ~^ image[12][4] + kernel[2][3] ~^ image[12][5] + kernel[2][4] ~^ image[12][6] + kernel[3][0] ~^ image[13][2] + kernel[3][1] ~^ image[13][3] + kernel[3][2] ~^ image[13][4] + kernel[3][3] ~^ image[13][5] + kernel[3][4] ~^ image[13][6] + kernel[4][0] ~^ image[14][2] + kernel[4][1] ~^ image[14][3] + kernel[4][2] ~^ image[14][4] + kernel[4][3] ~^ image[14][5] + kernel[4][4] ~^ image[14][6];
assign xor_sum[10][3] = kernel[0][0] ~^ image[10][3] + kernel[0][1] ~^ image[10][4] + kernel[0][2] ~^ image[10][5] + kernel[0][3] ~^ image[10][6] + kernel[0][4] ~^ image[10][7] + kernel[1][0] ~^ image[11][3] + kernel[1][1] ~^ image[11][4] + kernel[1][2] ~^ image[11][5] + kernel[1][3] ~^ image[11][6] + kernel[1][4] ~^ image[11][7] + kernel[2][0] ~^ image[12][3] + kernel[2][1] ~^ image[12][4] + kernel[2][2] ~^ image[12][5] + kernel[2][3] ~^ image[12][6] + kernel[2][4] ~^ image[12][7] + kernel[3][0] ~^ image[13][3] + kernel[3][1] ~^ image[13][4] + kernel[3][2] ~^ image[13][5] + kernel[3][3] ~^ image[13][6] + kernel[3][4] ~^ image[13][7] + kernel[4][0] ~^ image[14][3] + kernel[4][1] ~^ image[14][4] + kernel[4][2] ~^ image[14][5] + kernel[4][3] ~^ image[14][6] + kernel[4][4] ~^ image[14][7];
assign xor_sum[10][4] = kernel[0][0] ~^ image[10][4] + kernel[0][1] ~^ image[10][5] + kernel[0][2] ~^ image[10][6] + kernel[0][3] ~^ image[10][7] + kernel[0][4] ~^ image[10][8] + kernel[1][0] ~^ image[11][4] + kernel[1][1] ~^ image[11][5] + kernel[1][2] ~^ image[11][6] + kernel[1][3] ~^ image[11][7] + kernel[1][4] ~^ image[11][8] + kernel[2][0] ~^ image[12][4] + kernel[2][1] ~^ image[12][5] + kernel[2][2] ~^ image[12][6] + kernel[2][3] ~^ image[12][7] + kernel[2][4] ~^ image[12][8] + kernel[3][0] ~^ image[13][4] + kernel[3][1] ~^ image[13][5] + kernel[3][2] ~^ image[13][6] + kernel[3][3] ~^ image[13][7] + kernel[3][4] ~^ image[13][8] + kernel[4][0] ~^ image[14][4] + kernel[4][1] ~^ image[14][5] + kernel[4][2] ~^ image[14][6] + kernel[4][3] ~^ image[14][7] + kernel[4][4] ~^ image[14][8];
assign xor_sum[10][5] = kernel[0][0] ~^ image[10][5] + kernel[0][1] ~^ image[10][6] + kernel[0][2] ~^ image[10][7] + kernel[0][3] ~^ image[10][8] + kernel[0][4] ~^ image[10][9] + kernel[1][0] ~^ image[11][5] + kernel[1][1] ~^ image[11][6] + kernel[1][2] ~^ image[11][7] + kernel[1][3] ~^ image[11][8] + kernel[1][4] ~^ image[11][9] + kernel[2][0] ~^ image[12][5] + kernel[2][1] ~^ image[12][6] + kernel[2][2] ~^ image[12][7] + kernel[2][3] ~^ image[12][8] + kernel[2][4] ~^ image[12][9] + kernel[3][0] ~^ image[13][5] + kernel[3][1] ~^ image[13][6] + kernel[3][2] ~^ image[13][7] + kernel[3][3] ~^ image[13][8] + kernel[3][4] ~^ image[13][9] + kernel[4][0] ~^ image[14][5] + kernel[4][1] ~^ image[14][6] + kernel[4][2] ~^ image[14][7] + kernel[4][3] ~^ image[14][8] + kernel[4][4] ~^ image[14][9];
assign xor_sum[10][6] = kernel[0][0] ~^ image[10][6] + kernel[0][1] ~^ image[10][7] + kernel[0][2] ~^ image[10][8] + kernel[0][3] ~^ image[10][9] + kernel[0][4] ~^ image[10][10] + kernel[1][0] ~^ image[11][6] + kernel[1][1] ~^ image[11][7] + kernel[1][2] ~^ image[11][8] + kernel[1][3] ~^ image[11][9] + kernel[1][4] ~^ image[11][10] + kernel[2][0] ~^ image[12][6] + kernel[2][1] ~^ image[12][7] + kernel[2][2] ~^ image[12][8] + kernel[2][3] ~^ image[12][9] + kernel[2][4] ~^ image[12][10] + kernel[3][0] ~^ image[13][6] + kernel[3][1] ~^ image[13][7] + kernel[3][2] ~^ image[13][8] + kernel[3][3] ~^ image[13][9] + kernel[3][4] ~^ image[13][10] + kernel[4][0] ~^ image[14][6] + kernel[4][1] ~^ image[14][7] + kernel[4][2] ~^ image[14][8] + kernel[4][3] ~^ image[14][9] + kernel[4][4] ~^ image[14][10];
assign xor_sum[10][7] = kernel[0][0] ~^ image[10][7] + kernel[0][1] ~^ image[10][8] + kernel[0][2] ~^ image[10][9] + kernel[0][3] ~^ image[10][10] + kernel[0][4] ~^ image[10][11] + kernel[1][0] ~^ image[11][7] + kernel[1][1] ~^ image[11][8] + kernel[1][2] ~^ image[11][9] + kernel[1][3] ~^ image[11][10] + kernel[1][4] ~^ image[11][11] + kernel[2][0] ~^ image[12][7] + kernel[2][1] ~^ image[12][8] + kernel[2][2] ~^ image[12][9] + kernel[2][3] ~^ image[12][10] + kernel[2][4] ~^ image[12][11] + kernel[3][0] ~^ image[13][7] + kernel[3][1] ~^ image[13][8] + kernel[3][2] ~^ image[13][9] + kernel[3][3] ~^ image[13][10] + kernel[3][4] ~^ image[13][11] + kernel[4][0] ~^ image[14][7] + kernel[4][1] ~^ image[14][8] + kernel[4][2] ~^ image[14][9] + kernel[4][3] ~^ image[14][10] + kernel[4][4] ~^ image[14][11];
assign xor_sum[10][8] = kernel[0][0] ~^ image[10][8] + kernel[0][1] ~^ image[10][9] + kernel[0][2] ~^ image[10][10] + kernel[0][3] ~^ image[10][11] + kernel[0][4] ~^ image[10][12] + kernel[1][0] ~^ image[11][8] + kernel[1][1] ~^ image[11][9] + kernel[1][2] ~^ image[11][10] + kernel[1][3] ~^ image[11][11] + kernel[1][4] ~^ image[11][12] + kernel[2][0] ~^ image[12][8] + kernel[2][1] ~^ image[12][9] + kernel[2][2] ~^ image[12][10] + kernel[2][3] ~^ image[12][11] + kernel[2][4] ~^ image[12][12] + kernel[3][0] ~^ image[13][8] + kernel[3][1] ~^ image[13][9] + kernel[3][2] ~^ image[13][10] + kernel[3][3] ~^ image[13][11] + kernel[3][4] ~^ image[13][12] + kernel[4][0] ~^ image[14][8] + kernel[4][1] ~^ image[14][9] + kernel[4][2] ~^ image[14][10] + kernel[4][3] ~^ image[14][11] + kernel[4][4] ~^ image[14][12];
assign xor_sum[10][9] = kernel[0][0] ~^ image[10][9] + kernel[0][1] ~^ image[10][10] + kernel[0][2] ~^ image[10][11] + kernel[0][3] ~^ image[10][12] + kernel[0][4] ~^ image[10][13] + kernel[1][0] ~^ image[11][9] + kernel[1][1] ~^ image[11][10] + kernel[1][2] ~^ image[11][11] + kernel[1][3] ~^ image[11][12] + kernel[1][4] ~^ image[11][13] + kernel[2][0] ~^ image[12][9] + kernel[2][1] ~^ image[12][10] + kernel[2][2] ~^ image[12][11] + kernel[2][3] ~^ image[12][12] + kernel[2][4] ~^ image[12][13] + kernel[3][0] ~^ image[13][9] + kernel[3][1] ~^ image[13][10] + kernel[3][2] ~^ image[13][11] + kernel[3][3] ~^ image[13][12] + kernel[3][4] ~^ image[13][13] + kernel[4][0] ~^ image[14][9] + kernel[4][1] ~^ image[14][10] + kernel[4][2] ~^ image[14][11] + kernel[4][3] ~^ image[14][12] + kernel[4][4] ~^ image[14][13];
assign xor_sum[10][10] = kernel[0][0] ~^ image[10][10] + kernel[0][1] ~^ image[10][11] + kernel[0][2] ~^ image[10][12] + kernel[0][3] ~^ image[10][13] + kernel[0][4] ~^ image[10][14] + kernel[1][0] ~^ image[11][10] + kernel[1][1] ~^ image[11][11] + kernel[1][2] ~^ image[11][12] + kernel[1][3] ~^ image[11][13] + kernel[1][4] ~^ image[11][14] + kernel[2][0] ~^ image[12][10] + kernel[2][1] ~^ image[12][11] + kernel[2][2] ~^ image[12][12] + kernel[2][3] ~^ image[12][13] + kernel[2][4] ~^ image[12][14] + kernel[3][0] ~^ image[13][10] + kernel[3][1] ~^ image[13][11] + kernel[3][2] ~^ image[13][12] + kernel[3][3] ~^ image[13][13] + kernel[3][4] ~^ image[13][14] + kernel[4][0] ~^ image[14][10] + kernel[4][1] ~^ image[14][11] + kernel[4][2] ~^ image[14][12] + kernel[4][3] ~^ image[14][13] + kernel[4][4] ~^ image[14][14];
assign xor_sum[10][11] = kernel[0][0] ~^ image[10][11] + kernel[0][1] ~^ image[10][12] + kernel[0][2] ~^ image[10][13] + kernel[0][3] ~^ image[10][14] + kernel[0][4] ~^ image[10][15] + kernel[1][0] ~^ image[11][11] + kernel[1][1] ~^ image[11][12] + kernel[1][2] ~^ image[11][13] + kernel[1][3] ~^ image[11][14] + kernel[1][4] ~^ image[11][15] + kernel[2][0] ~^ image[12][11] + kernel[2][1] ~^ image[12][12] + kernel[2][2] ~^ image[12][13] + kernel[2][3] ~^ image[12][14] + kernel[2][4] ~^ image[12][15] + kernel[3][0] ~^ image[13][11] + kernel[3][1] ~^ image[13][12] + kernel[3][2] ~^ image[13][13] + kernel[3][3] ~^ image[13][14] + kernel[3][4] ~^ image[13][15] + kernel[4][0] ~^ image[14][11] + kernel[4][1] ~^ image[14][12] + kernel[4][2] ~^ image[14][13] + kernel[4][3] ~^ image[14][14] + kernel[4][4] ~^ image[14][15];
assign xor_sum[10][12] = kernel[0][0] ~^ image[10][12] + kernel[0][1] ~^ image[10][13] + kernel[0][2] ~^ image[10][14] + kernel[0][3] ~^ image[10][15] + kernel[0][4] ~^ image[10][16] + kernel[1][0] ~^ image[11][12] + kernel[1][1] ~^ image[11][13] + kernel[1][2] ~^ image[11][14] + kernel[1][3] ~^ image[11][15] + kernel[1][4] ~^ image[11][16] + kernel[2][0] ~^ image[12][12] + kernel[2][1] ~^ image[12][13] + kernel[2][2] ~^ image[12][14] + kernel[2][3] ~^ image[12][15] + kernel[2][4] ~^ image[12][16] + kernel[3][0] ~^ image[13][12] + kernel[3][1] ~^ image[13][13] + kernel[3][2] ~^ image[13][14] + kernel[3][3] ~^ image[13][15] + kernel[3][4] ~^ image[13][16] + kernel[4][0] ~^ image[14][12] + kernel[4][1] ~^ image[14][13] + kernel[4][2] ~^ image[14][14] + kernel[4][3] ~^ image[14][15] + kernel[4][4] ~^ image[14][16];
assign xor_sum[10][13] = kernel[0][0] ~^ image[10][13] + kernel[0][1] ~^ image[10][14] + kernel[0][2] ~^ image[10][15] + kernel[0][3] ~^ image[10][16] + kernel[0][4] ~^ image[10][17] + kernel[1][0] ~^ image[11][13] + kernel[1][1] ~^ image[11][14] + kernel[1][2] ~^ image[11][15] + kernel[1][3] ~^ image[11][16] + kernel[1][4] ~^ image[11][17] + kernel[2][0] ~^ image[12][13] + kernel[2][1] ~^ image[12][14] + kernel[2][2] ~^ image[12][15] + kernel[2][3] ~^ image[12][16] + kernel[2][4] ~^ image[12][17] + kernel[3][0] ~^ image[13][13] + kernel[3][1] ~^ image[13][14] + kernel[3][2] ~^ image[13][15] + kernel[3][3] ~^ image[13][16] + kernel[3][4] ~^ image[13][17] + kernel[4][0] ~^ image[14][13] + kernel[4][1] ~^ image[14][14] + kernel[4][2] ~^ image[14][15] + kernel[4][3] ~^ image[14][16] + kernel[4][4] ~^ image[14][17];
assign xor_sum[10][14] = kernel[0][0] ~^ image[10][14] + kernel[0][1] ~^ image[10][15] + kernel[0][2] ~^ image[10][16] + kernel[0][3] ~^ image[10][17] + kernel[0][4] ~^ image[10][18] + kernel[1][0] ~^ image[11][14] + kernel[1][1] ~^ image[11][15] + kernel[1][2] ~^ image[11][16] + kernel[1][3] ~^ image[11][17] + kernel[1][4] ~^ image[11][18] + kernel[2][0] ~^ image[12][14] + kernel[2][1] ~^ image[12][15] + kernel[2][2] ~^ image[12][16] + kernel[2][3] ~^ image[12][17] + kernel[2][4] ~^ image[12][18] + kernel[3][0] ~^ image[13][14] + kernel[3][1] ~^ image[13][15] + kernel[3][2] ~^ image[13][16] + kernel[3][3] ~^ image[13][17] + kernel[3][4] ~^ image[13][18] + kernel[4][0] ~^ image[14][14] + kernel[4][1] ~^ image[14][15] + kernel[4][2] ~^ image[14][16] + kernel[4][3] ~^ image[14][17] + kernel[4][4] ~^ image[14][18];
assign xor_sum[10][15] = kernel[0][0] ~^ image[10][15] + kernel[0][1] ~^ image[10][16] + kernel[0][2] ~^ image[10][17] + kernel[0][3] ~^ image[10][18] + kernel[0][4] ~^ image[10][19] + kernel[1][0] ~^ image[11][15] + kernel[1][1] ~^ image[11][16] + kernel[1][2] ~^ image[11][17] + kernel[1][3] ~^ image[11][18] + kernel[1][4] ~^ image[11][19] + kernel[2][0] ~^ image[12][15] + kernel[2][1] ~^ image[12][16] + kernel[2][2] ~^ image[12][17] + kernel[2][3] ~^ image[12][18] + kernel[2][4] ~^ image[12][19] + kernel[3][0] ~^ image[13][15] + kernel[3][1] ~^ image[13][16] + kernel[3][2] ~^ image[13][17] + kernel[3][3] ~^ image[13][18] + kernel[3][4] ~^ image[13][19] + kernel[4][0] ~^ image[14][15] + kernel[4][1] ~^ image[14][16] + kernel[4][2] ~^ image[14][17] + kernel[4][3] ~^ image[14][18] + kernel[4][4] ~^ image[14][19];
assign xor_sum[10][16] = kernel[0][0] ~^ image[10][16] + kernel[0][1] ~^ image[10][17] + kernel[0][2] ~^ image[10][18] + kernel[0][3] ~^ image[10][19] + kernel[0][4] ~^ image[10][20] + kernel[1][0] ~^ image[11][16] + kernel[1][1] ~^ image[11][17] + kernel[1][2] ~^ image[11][18] + kernel[1][3] ~^ image[11][19] + kernel[1][4] ~^ image[11][20] + kernel[2][0] ~^ image[12][16] + kernel[2][1] ~^ image[12][17] + kernel[2][2] ~^ image[12][18] + kernel[2][3] ~^ image[12][19] + kernel[2][4] ~^ image[12][20] + kernel[3][0] ~^ image[13][16] + kernel[3][1] ~^ image[13][17] + kernel[3][2] ~^ image[13][18] + kernel[3][3] ~^ image[13][19] + kernel[3][4] ~^ image[13][20] + kernel[4][0] ~^ image[14][16] + kernel[4][1] ~^ image[14][17] + kernel[4][2] ~^ image[14][18] + kernel[4][3] ~^ image[14][19] + kernel[4][4] ~^ image[14][20];
assign xor_sum[10][17] = kernel[0][0] ~^ image[10][17] + kernel[0][1] ~^ image[10][18] + kernel[0][2] ~^ image[10][19] + kernel[0][3] ~^ image[10][20] + kernel[0][4] ~^ image[10][21] + kernel[1][0] ~^ image[11][17] + kernel[1][1] ~^ image[11][18] + kernel[1][2] ~^ image[11][19] + kernel[1][3] ~^ image[11][20] + kernel[1][4] ~^ image[11][21] + kernel[2][0] ~^ image[12][17] + kernel[2][1] ~^ image[12][18] + kernel[2][2] ~^ image[12][19] + kernel[2][3] ~^ image[12][20] + kernel[2][4] ~^ image[12][21] + kernel[3][0] ~^ image[13][17] + kernel[3][1] ~^ image[13][18] + kernel[3][2] ~^ image[13][19] + kernel[3][3] ~^ image[13][20] + kernel[3][4] ~^ image[13][21] + kernel[4][0] ~^ image[14][17] + kernel[4][1] ~^ image[14][18] + kernel[4][2] ~^ image[14][19] + kernel[4][3] ~^ image[14][20] + kernel[4][4] ~^ image[14][21];
assign xor_sum[10][18] = kernel[0][0] ~^ image[10][18] + kernel[0][1] ~^ image[10][19] + kernel[0][2] ~^ image[10][20] + kernel[0][3] ~^ image[10][21] + kernel[0][4] ~^ image[10][22] + kernel[1][0] ~^ image[11][18] + kernel[1][1] ~^ image[11][19] + kernel[1][2] ~^ image[11][20] + kernel[1][3] ~^ image[11][21] + kernel[1][4] ~^ image[11][22] + kernel[2][0] ~^ image[12][18] + kernel[2][1] ~^ image[12][19] + kernel[2][2] ~^ image[12][20] + kernel[2][3] ~^ image[12][21] + kernel[2][4] ~^ image[12][22] + kernel[3][0] ~^ image[13][18] + kernel[3][1] ~^ image[13][19] + kernel[3][2] ~^ image[13][20] + kernel[3][3] ~^ image[13][21] + kernel[3][4] ~^ image[13][22] + kernel[4][0] ~^ image[14][18] + kernel[4][1] ~^ image[14][19] + kernel[4][2] ~^ image[14][20] + kernel[4][3] ~^ image[14][21] + kernel[4][4] ~^ image[14][22];
assign xor_sum[10][19] = kernel[0][0] ~^ image[10][19] + kernel[0][1] ~^ image[10][20] + kernel[0][2] ~^ image[10][21] + kernel[0][3] ~^ image[10][22] + kernel[0][4] ~^ image[10][23] + kernel[1][0] ~^ image[11][19] + kernel[1][1] ~^ image[11][20] + kernel[1][2] ~^ image[11][21] + kernel[1][3] ~^ image[11][22] + kernel[1][4] ~^ image[11][23] + kernel[2][0] ~^ image[12][19] + kernel[2][1] ~^ image[12][20] + kernel[2][2] ~^ image[12][21] + kernel[2][3] ~^ image[12][22] + kernel[2][4] ~^ image[12][23] + kernel[3][0] ~^ image[13][19] + kernel[3][1] ~^ image[13][20] + kernel[3][2] ~^ image[13][21] + kernel[3][3] ~^ image[13][22] + kernel[3][4] ~^ image[13][23] + kernel[4][0] ~^ image[14][19] + kernel[4][1] ~^ image[14][20] + kernel[4][2] ~^ image[14][21] + kernel[4][3] ~^ image[14][22] + kernel[4][4] ~^ image[14][23];
assign xor_sum[10][20] = kernel[0][0] ~^ image[10][20] + kernel[0][1] ~^ image[10][21] + kernel[0][2] ~^ image[10][22] + kernel[0][3] ~^ image[10][23] + kernel[0][4] ~^ image[10][24] + kernel[1][0] ~^ image[11][20] + kernel[1][1] ~^ image[11][21] + kernel[1][2] ~^ image[11][22] + kernel[1][3] ~^ image[11][23] + kernel[1][4] ~^ image[11][24] + kernel[2][0] ~^ image[12][20] + kernel[2][1] ~^ image[12][21] + kernel[2][2] ~^ image[12][22] + kernel[2][3] ~^ image[12][23] + kernel[2][4] ~^ image[12][24] + kernel[3][0] ~^ image[13][20] + kernel[3][1] ~^ image[13][21] + kernel[3][2] ~^ image[13][22] + kernel[3][3] ~^ image[13][23] + kernel[3][4] ~^ image[13][24] + kernel[4][0] ~^ image[14][20] + kernel[4][1] ~^ image[14][21] + kernel[4][2] ~^ image[14][22] + kernel[4][3] ~^ image[14][23] + kernel[4][4] ~^ image[14][24];
assign xor_sum[10][21] = kernel[0][0] ~^ image[10][21] + kernel[0][1] ~^ image[10][22] + kernel[0][2] ~^ image[10][23] + kernel[0][3] ~^ image[10][24] + kernel[0][4] ~^ image[10][25] + kernel[1][0] ~^ image[11][21] + kernel[1][1] ~^ image[11][22] + kernel[1][2] ~^ image[11][23] + kernel[1][3] ~^ image[11][24] + kernel[1][4] ~^ image[11][25] + kernel[2][0] ~^ image[12][21] + kernel[2][1] ~^ image[12][22] + kernel[2][2] ~^ image[12][23] + kernel[2][3] ~^ image[12][24] + kernel[2][4] ~^ image[12][25] + kernel[3][0] ~^ image[13][21] + kernel[3][1] ~^ image[13][22] + kernel[3][2] ~^ image[13][23] + kernel[3][3] ~^ image[13][24] + kernel[3][4] ~^ image[13][25] + kernel[4][0] ~^ image[14][21] + kernel[4][1] ~^ image[14][22] + kernel[4][2] ~^ image[14][23] + kernel[4][3] ~^ image[14][24] + kernel[4][4] ~^ image[14][25];
assign xor_sum[10][22] = kernel[0][0] ~^ image[10][22] + kernel[0][1] ~^ image[10][23] + kernel[0][2] ~^ image[10][24] + kernel[0][3] ~^ image[10][25] + kernel[0][4] ~^ image[10][26] + kernel[1][0] ~^ image[11][22] + kernel[1][1] ~^ image[11][23] + kernel[1][2] ~^ image[11][24] + kernel[1][3] ~^ image[11][25] + kernel[1][4] ~^ image[11][26] + kernel[2][0] ~^ image[12][22] + kernel[2][1] ~^ image[12][23] + kernel[2][2] ~^ image[12][24] + kernel[2][3] ~^ image[12][25] + kernel[2][4] ~^ image[12][26] + kernel[3][0] ~^ image[13][22] + kernel[3][1] ~^ image[13][23] + kernel[3][2] ~^ image[13][24] + kernel[3][3] ~^ image[13][25] + kernel[3][4] ~^ image[13][26] + kernel[4][0] ~^ image[14][22] + kernel[4][1] ~^ image[14][23] + kernel[4][2] ~^ image[14][24] + kernel[4][3] ~^ image[14][25] + kernel[4][4] ~^ image[14][26];
assign xor_sum[10][23] = kernel[0][0] ~^ image[10][23] + kernel[0][1] ~^ image[10][24] + kernel[0][2] ~^ image[10][25] + kernel[0][3] ~^ image[10][26] + kernel[0][4] ~^ image[10][27] + kernel[1][0] ~^ image[11][23] + kernel[1][1] ~^ image[11][24] + kernel[1][2] ~^ image[11][25] + kernel[1][3] ~^ image[11][26] + kernel[1][4] ~^ image[11][27] + kernel[2][0] ~^ image[12][23] + kernel[2][1] ~^ image[12][24] + kernel[2][2] ~^ image[12][25] + kernel[2][3] ~^ image[12][26] + kernel[2][4] ~^ image[12][27] + kernel[3][0] ~^ image[13][23] + kernel[3][1] ~^ image[13][24] + kernel[3][2] ~^ image[13][25] + kernel[3][3] ~^ image[13][26] + kernel[3][4] ~^ image[13][27] + kernel[4][0] ~^ image[14][23] + kernel[4][1] ~^ image[14][24] + kernel[4][2] ~^ image[14][25] + kernel[4][3] ~^ image[14][26] + kernel[4][4] ~^ image[14][27];
assign xor_sum[11][0] = kernel[0][0] ~^ image[11][0] + kernel[0][1] ~^ image[11][1] + kernel[0][2] ~^ image[11][2] + kernel[0][3] ~^ image[11][3] + kernel[0][4] ~^ image[11][4] + kernel[1][0] ~^ image[12][0] + kernel[1][1] ~^ image[12][1] + kernel[1][2] ~^ image[12][2] + kernel[1][3] ~^ image[12][3] + kernel[1][4] ~^ image[12][4] + kernel[2][0] ~^ image[13][0] + kernel[2][1] ~^ image[13][1] + kernel[2][2] ~^ image[13][2] + kernel[2][3] ~^ image[13][3] + kernel[2][4] ~^ image[13][4] + kernel[3][0] ~^ image[14][0] + kernel[3][1] ~^ image[14][1] + kernel[3][2] ~^ image[14][2] + kernel[3][3] ~^ image[14][3] + kernel[3][4] ~^ image[14][4] + kernel[4][0] ~^ image[15][0] + kernel[4][1] ~^ image[15][1] + kernel[4][2] ~^ image[15][2] + kernel[4][3] ~^ image[15][3] + kernel[4][4] ~^ image[15][4];
assign xor_sum[11][1] = kernel[0][0] ~^ image[11][1] + kernel[0][1] ~^ image[11][2] + kernel[0][2] ~^ image[11][3] + kernel[0][3] ~^ image[11][4] + kernel[0][4] ~^ image[11][5] + kernel[1][0] ~^ image[12][1] + kernel[1][1] ~^ image[12][2] + kernel[1][2] ~^ image[12][3] + kernel[1][3] ~^ image[12][4] + kernel[1][4] ~^ image[12][5] + kernel[2][0] ~^ image[13][1] + kernel[2][1] ~^ image[13][2] + kernel[2][2] ~^ image[13][3] + kernel[2][3] ~^ image[13][4] + kernel[2][4] ~^ image[13][5] + kernel[3][0] ~^ image[14][1] + kernel[3][1] ~^ image[14][2] + kernel[3][2] ~^ image[14][3] + kernel[3][3] ~^ image[14][4] + kernel[3][4] ~^ image[14][5] + kernel[4][0] ~^ image[15][1] + kernel[4][1] ~^ image[15][2] + kernel[4][2] ~^ image[15][3] + kernel[4][3] ~^ image[15][4] + kernel[4][4] ~^ image[15][5];
assign xor_sum[11][2] = kernel[0][0] ~^ image[11][2] + kernel[0][1] ~^ image[11][3] + kernel[0][2] ~^ image[11][4] + kernel[0][3] ~^ image[11][5] + kernel[0][4] ~^ image[11][6] + kernel[1][0] ~^ image[12][2] + kernel[1][1] ~^ image[12][3] + kernel[1][2] ~^ image[12][4] + kernel[1][3] ~^ image[12][5] + kernel[1][4] ~^ image[12][6] + kernel[2][0] ~^ image[13][2] + kernel[2][1] ~^ image[13][3] + kernel[2][2] ~^ image[13][4] + kernel[2][3] ~^ image[13][5] + kernel[2][4] ~^ image[13][6] + kernel[3][0] ~^ image[14][2] + kernel[3][1] ~^ image[14][3] + kernel[3][2] ~^ image[14][4] + kernel[3][3] ~^ image[14][5] + kernel[3][4] ~^ image[14][6] + kernel[4][0] ~^ image[15][2] + kernel[4][1] ~^ image[15][3] + kernel[4][2] ~^ image[15][4] + kernel[4][3] ~^ image[15][5] + kernel[4][4] ~^ image[15][6];
assign xor_sum[11][3] = kernel[0][0] ~^ image[11][3] + kernel[0][1] ~^ image[11][4] + kernel[0][2] ~^ image[11][5] + kernel[0][3] ~^ image[11][6] + kernel[0][4] ~^ image[11][7] + kernel[1][0] ~^ image[12][3] + kernel[1][1] ~^ image[12][4] + kernel[1][2] ~^ image[12][5] + kernel[1][3] ~^ image[12][6] + kernel[1][4] ~^ image[12][7] + kernel[2][0] ~^ image[13][3] + kernel[2][1] ~^ image[13][4] + kernel[2][2] ~^ image[13][5] + kernel[2][3] ~^ image[13][6] + kernel[2][4] ~^ image[13][7] + kernel[3][0] ~^ image[14][3] + kernel[3][1] ~^ image[14][4] + kernel[3][2] ~^ image[14][5] + kernel[3][3] ~^ image[14][6] + kernel[3][4] ~^ image[14][7] + kernel[4][0] ~^ image[15][3] + kernel[4][1] ~^ image[15][4] + kernel[4][2] ~^ image[15][5] + kernel[4][3] ~^ image[15][6] + kernel[4][4] ~^ image[15][7];
assign xor_sum[11][4] = kernel[0][0] ~^ image[11][4] + kernel[0][1] ~^ image[11][5] + kernel[0][2] ~^ image[11][6] + kernel[0][3] ~^ image[11][7] + kernel[0][4] ~^ image[11][8] + kernel[1][0] ~^ image[12][4] + kernel[1][1] ~^ image[12][5] + kernel[1][2] ~^ image[12][6] + kernel[1][3] ~^ image[12][7] + kernel[1][4] ~^ image[12][8] + kernel[2][0] ~^ image[13][4] + kernel[2][1] ~^ image[13][5] + kernel[2][2] ~^ image[13][6] + kernel[2][3] ~^ image[13][7] + kernel[2][4] ~^ image[13][8] + kernel[3][0] ~^ image[14][4] + kernel[3][1] ~^ image[14][5] + kernel[3][2] ~^ image[14][6] + kernel[3][3] ~^ image[14][7] + kernel[3][4] ~^ image[14][8] + kernel[4][0] ~^ image[15][4] + kernel[4][1] ~^ image[15][5] + kernel[4][2] ~^ image[15][6] + kernel[4][3] ~^ image[15][7] + kernel[4][4] ~^ image[15][8];
assign xor_sum[11][5] = kernel[0][0] ~^ image[11][5] + kernel[0][1] ~^ image[11][6] + kernel[0][2] ~^ image[11][7] + kernel[0][3] ~^ image[11][8] + kernel[0][4] ~^ image[11][9] + kernel[1][0] ~^ image[12][5] + kernel[1][1] ~^ image[12][6] + kernel[1][2] ~^ image[12][7] + kernel[1][3] ~^ image[12][8] + kernel[1][4] ~^ image[12][9] + kernel[2][0] ~^ image[13][5] + kernel[2][1] ~^ image[13][6] + kernel[2][2] ~^ image[13][7] + kernel[2][3] ~^ image[13][8] + kernel[2][4] ~^ image[13][9] + kernel[3][0] ~^ image[14][5] + kernel[3][1] ~^ image[14][6] + kernel[3][2] ~^ image[14][7] + kernel[3][3] ~^ image[14][8] + kernel[3][4] ~^ image[14][9] + kernel[4][0] ~^ image[15][5] + kernel[4][1] ~^ image[15][6] + kernel[4][2] ~^ image[15][7] + kernel[4][3] ~^ image[15][8] + kernel[4][4] ~^ image[15][9];
assign xor_sum[11][6] = kernel[0][0] ~^ image[11][6] + kernel[0][1] ~^ image[11][7] + kernel[0][2] ~^ image[11][8] + kernel[0][3] ~^ image[11][9] + kernel[0][4] ~^ image[11][10] + kernel[1][0] ~^ image[12][6] + kernel[1][1] ~^ image[12][7] + kernel[1][2] ~^ image[12][8] + kernel[1][3] ~^ image[12][9] + kernel[1][4] ~^ image[12][10] + kernel[2][0] ~^ image[13][6] + kernel[2][1] ~^ image[13][7] + kernel[2][2] ~^ image[13][8] + kernel[2][3] ~^ image[13][9] + kernel[2][4] ~^ image[13][10] + kernel[3][0] ~^ image[14][6] + kernel[3][1] ~^ image[14][7] + kernel[3][2] ~^ image[14][8] + kernel[3][3] ~^ image[14][9] + kernel[3][4] ~^ image[14][10] + kernel[4][0] ~^ image[15][6] + kernel[4][1] ~^ image[15][7] + kernel[4][2] ~^ image[15][8] + kernel[4][3] ~^ image[15][9] + kernel[4][4] ~^ image[15][10];
assign xor_sum[11][7] = kernel[0][0] ~^ image[11][7] + kernel[0][1] ~^ image[11][8] + kernel[0][2] ~^ image[11][9] + kernel[0][3] ~^ image[11][10] + kernel[0][4] ~^ image[11][11] + kernel[1][0] ~^ image[12][7] + kernel[1][1] ~^ image[12][8] + kernel[1][2] ~^ image[12][9] + kernel[1][3] ~^ image[12][10] + kernel[1][4] ~^ image[12][11] + kernel[2][0] ~^ image[13][7] + kernel[2][1] ~^ image[13][8] + kernel[2][2] ~^ image[13][9] + kernel[2][3] ~^ image[13][10] + kernel[2][4] ~^ image[13][11] + kernel[3][0] ~^ image[14][7] + kernel[3][1] ~^ image[14][8] + kernel[3][2] ~^ image[14][9] + kernel[3][3] ~^ image[14][10] + kernel[3][4] ~^ image[14][11] + kernel[4][0] ~^ image[15][7] + kernel[4][1] ~^ image[15][8] + kernel[4][2] ~^ image[15][9] + kernel[4][3] ~^ image[15][10] + kernel[4][4] ~^ image[15][11];
assign xor_sum[11][8] = kernel[0][0] ~^ image[11][8] + kernel[0][1] ~^ image[11][9] + kernel[0][2] ~^ image[11][10] + kernel[0][3] ~^ image[11][11] + kernel[0][4] ~^ image[11][12] + kernel[1][0] ~^ image[12][8] + kernel[1][1] ~^ image[12][9] + kernel[1][2] ~^ image[12][10] + kernel[1][3] ~^ image[12][11] + kernel[1][4] ~^ image[12][12] + kernel[2][0] ~^ image[13][8] + kernel[2][1] ~^ image[13][9] + kernel[2][2] ~^ image[13][10] + kernel[2][3] ~^ image[13][11] + kernel[2][4] ~^ image[13][12] + kernel[3][0] ~^ image[14][8] + kernel[3][1] ~^ image[14][9] + kernel[3][2] ~^ image[14][10] + kernel[3][3] ~^ image[14][11] + kernel[3][4] ~^ image[14][12] + kernel[4][0] ~^ image[15][8] + kernel[4][1] ~^ image[15][9] + kernel[4][2] ~^ image[15][10] + kernel[4][3] ~^ image[15][11] + kernel[4][4] ~^ image[15][12];
assign xor_sum[11][9] = kernel[0][0] ~^ image[11][9] + kernel[0][1] ~^ image[11][10] + kernel[0][2] ~^ image[11][11] + kernel[0][3] ~^ image[11][12] + kernel[0][4] ~^ image[11][13] + kernel[1][0] ~^ image[12][9] + kernel[1][1] ~^ image[12][10] + kernel[1][2] ~^ image[12][11] + kernel[1][3] ~^ image[12][12] + kernel[1][4] ~^ image[12][13] + kernel[2][0] ~^ image[13][9] + kernel[2][1] ~^ image[13][10] + kernel[2][2] ~^ image[13][11] + kernel[2][3] ~^ image[13][12] + kernel[2][4] ~^ image[13][13] + kernel[3][0] ~^ image[14][9] + kernel[3][1] ~^ image[14][10] + kernel[3][2] ~^ image[14][11] + kernel[3][3] ~^ image[14][12] + kernel[3][4] ~^ image[14][13] + kernel[4][0] ~^ image[15][9] + kernel[4][1] ~^ image[15][10] + kernel[4][2] ~^ image[15][11] + kernel[4][3] ~^ image[15][12] + kernel[4][4] ~^ image[15][13];
assign xor_sum[11][10] = kernel[0][0] ~^ image[11][10] + kernel[0][1] ~^ image[11][11] + kernel[0][2] ~^ image[11][12] + kernel[0][3] ~^ image[11][13] + kernel[0][4] ~^ image[11][14] + kernel[1][0] ~^ image[12][10] + kernel[1][1] ~^ image[12][11] + kernel[1][2] ~^ image[12][12] + kernel[1][3] ~^ image[12][13] + kernel[1][4] ~^ image[12][14] + kernel[2][0] ~^ image[13][10] + kernel[2][1] ~^ image[13][11] + kernel[2][2] ~^ image[13][12] + kernel[2][3] ~^ image[13][13] + kernel[2][4] ~^ image[13][14] + kernel[3][0] ~^ image[14][10] + kernel[3][1] ~^ image[14][11] + kernel[3][2] ~^ image[14][12] + kernel[3][3] ~^ image[14][13] + kernel[3][4] ~^ image[14][14] + kernel[4][0] ~^ image[15][10] + kernel[4][1] ~^ image[15][11] + kernel[4][2] ~^ image[15][12] + kernel[4][3] ~^ image[15][13] + kernel[4][4] ~^ image[15][14];
assign xor_sum[11][11] = kernel[0][0] ~^ image[11][11] + kernel[0][1] ~^ image[11][12] + kernel[0][2] ~^ image[11][13] + kernel[0][3] ~^ image[11][14] + kernel[0][4] ~^ image[11][15] + kernel[1][0] ~^ image[12][11] + kernel[1][1] ~^ image[12][12] + kernel[1][2] ~^ image[12][13] + kernel[1][3] ~^ image[12][14] + kernel[1][4] ~^ image[12][15] + kernel[2][0] ~^ image[13][11] + kernel[2][1] ~^ image[13][12] + kernel[2][2] ~^ image[13][13] + kernel[2][3] ~^ image[13][14] + kernel[2][4] ~^ image[13][15] + kernel[3][0] ~^ image[14][11] + kernel[3][1] ~^ image[14][12] + kernel[3][2] ~^ image[14][13] + kernel[3][3] ~^ image[14][14] + kernel[3][4] ~^ image[14][15] + kernel[4][0] ~^ image[15][11] + kernel[4][1] ~^ image[15][12] + kernel[4][2] ~^ image[15][13] + kernel[4][3] ~^ image[15][14] + kernel[4][4] ~^ image[15][15];
assign xor_sum[11][12] = kernel[0][0] ~^ image[11][12] + kernel[0][1] ~^ image[11][13] + kernel[0][2] ~^ image[11][14] + kernel[0][3] ~^ image[11][15] + kernel[0][4] ~^ image[11][16] + kernel[1][0] ~^ image[12][12] + kernel[1][1] ~^ image[12][13] + kernel[1][2] ~^ image[12][14] + kernel[1][3] ~^ image[12][15] + kernel[1][4] ~^ image[12][16] + kernel[2][0] ~^ image[13][12] + kernel[2][1] ~^ image[13][13] + kernel[2][2] ~^ image[13][14] + kernel[2][3] ~^ image[13][15] + kernel[2][4] ~^ image[13][16] + kernel[3][0] ~^ image[14][12] + kernel[3][1] ~^ image[14][13] + kernel[3][2] ~^ image[14][14] + kernel[3][3] ~^ image[14][15] + kernel[3][4] ~^ image[14][16] + kernel[4][0] ~^ image[15][12] + kernel[4][1] ~^ image[15][13] + kernel[4][2] ~^ image[15][14] + kernel[4][3] ~^ image[15][15] + kernel[4][4] ~^ image[15][16];
assign xor_sum[11][13] = kernel[0][0] ~^ image[11][13] + kernel[0][1] ~^ image[11][14] + kernel[0][2] ~^ image[11][15] + kernel[0][3] ~^ image[11][16] + kernel[0][4] ~^ image[11][17] + kernel[1][0] ~^ image[12][13] + kernel[1][1] ~^ image[12][14] + kernel[1][2] ~^ image[12][15] + kernel[1][3] ~^ image[12][16] + kernel[1][4] ~^ image[12][17] + kernel[2][0] ~^ image[13][13] + kernel[2][1] ~^ image[13][14] + kernel[2][2] ~^ image[13][15] + kernel[2][3] ~^ image[13][16] + kernel[2][4] ~^ image[13][17] + kernel[3][0] ~^ image[14][13] + kernel[3][1] ~^ image[14][14] + kernel[3][2] ~^ image[14][15] + kernel[3][3] ~^ image[14][16] + kernel[3][4] ~^ image[14][17] + kernel[4][0] ~^ image[15][13] + kernel[4][1] ~^ image[15][14] + kernel[4][2] ~^ image[15][15] + kernel[4][3] ~^ image[15][16] + kernel[4][4] ~^ image[15][17];
assign xor_sum[11][14] = kernel[0][0] ~^ image[11][14] + kernel[0][1] ~^ image[11][15] + kernel[0][2] ~^ image[11][16] + kernel[0][3] ~^ image[11][17] + kernel[0][4] ~^ image[11][18] + kernel[1][0] ~^ image[12][14] + kernel[1][1] ~^ image[12][15] + kernel[1][2] ~^ image[12][16] + kernel[1][3] ~^ image[12][17] + kernel[1][4] ~^ image[12][18] + kernel[2][0] ~^ image[13][14] + kernel[2][1] ~^ image[13][15] + kernel[2][2] ~^ image[13][16] + kernel[2][3] ~^ image[13][17] + kernel[2][4] ~^ image[13][18] + kernel[3][0] ~^ image[14][14] + kernel[3][1] ~^ image[14][15] + kernel[3][2] ~^ image[14][16] + kernel[3][3] ~^ image[14][17] + kernel[3][4] ~^ image[14][18] + kernel[4][0] ~^ image[15][14] + kernel[4][1] ~^ image[15][15] + kernel[4][2] ~^ image[15][16] + kernel[4][3] ~^ image[15][17] + kernel[4][4] ~^ image[15][18];
assign xor_sum[11][15] = kernel[0][0] ~^ image[11][15] + kernel[0][1] ~^ image[11][16] + kernel[0][2] ~^ image[11][17] + kernel[0][3] ~^ image[11][18] + kernel[0][4] ~^ image[11][19] + kernel[1][0] ~^ image[12][15] + kernel[1][1] ~^ image[12][16] + kernel[1][2] ~^ image[12][17] + kernel[1][3] ~^ image[12][18] + kernel[1][4] ~^ image[12][19] + kernel[2][0] ~^ image[13][15] + kernel[2][1] ~^ image[13][16] + kernel[2][2] ~^ image[13][17] + kernel[2][3] ~^ image[13][18] + kernel[2][4] ~^ image[13][19] + kernel[3][0] ~^ image[14][15] + kernel[3][1] ~^ image[14][16] + kernel[3][2] ~^ image[14][17] + kernel[3][3] ~^ image[14][18] + kernel[3][4] ~^ image[14][19] + kernel[4][0] ~^ image[15][15] + kernel[4][1] ~^ image[15][16] + kernel[4][2] ~^ image[15][17] + kernel[4][3] ~^ image[15][18] + kernel[4][4] ~^ image[15][19];
assign xor_sum[11][16] = kernel[0][0] ~^ image[11][16] + kernel[0][1] ~^ image[11][17] + kernel[0][2] ~^ image[11][18] + kernel[0][3] ~^ image[11][19] + kernel[0][4] ~^ image[11][20] + kernel[1][0] ~^ image[12][16] + kernel[1][1] ~^ image[12][17] + kernel[1][2] ~^ image[12][18] + kernel[1][3] ~^ image[12][19] + kernel[1][4] ~^ image[12][20] + kernel[2][0] ~^ image[13][16] + kernel[2][1] ~^ image[13][17] + kernel[2][2] ~^ image[13][18] + kernel[2][3] ~^ image[13][19] + kernel[2][4] ~^ image[13][20] + kernel[3][0] ~^ image[14][16] + kernel[3][1] ~^ image[14][17] + kernel[3][2] ~^ image[14][18] + kernel[3][3] ~^ image[14][19] + kernel[3][4] ~^ image[14][20] + kernel[4][0] ~^ image[15][16] + kernel[4][1] ~^ image[15][17] + kernel[4][2] ~^ image[15][18] + kernel[4][3] ~^ image[15][19] + kernel[4][4] ~^ image[15][20];
assign xor_sum[11][17] = kernel[0][0] ~^ image[11][17] + kernel[0][1] ~^ image[11][18] + kernel[0][2] ~^ image[11][19] + kernel[0][3] ~^ image[11][20] + kernel[0][4] ~^ image[11][21] + kernel[1][0] ~^ image[12][17] + kernel[1][1] ~^ image[12][18] + kernel[1][2] ~^ image[12][19] + kernel[1][3] ~^ image[12][20] + kernel[1][4] ~^ image[12][21] + kernel[2][0] ~^ image[13][17] + kernel[2][1] ~^ image[13][18] + kernel[2][2] ~^ image[13][19] + kernel[2][3] ~^ image[13][20] + kernel[2][4] ~^ image[13][21] + kernel[3][0] ~^ image[14][17] + kernel[3][1] ~^ image[14][18] + kernel[3][2] ~^ image[14][19] + kernel[3][3] ~^ image[14][20] + kernel[3][4] ~^ image[14][21] + kernel[4][0] ~^ image[15][17] + kernel[4][1] ~^ image[15][18] + kernel[4][2] ~^ image[15][19] + kernel[4][3] ~^ image[15][20] + kernel[4][4] ~^ image[15][21];
assign xor_sum[11][18] = kernel[0][0] ~^ image[11][18] + kernel[0][1] ~^ image[11][19] + kernel[0][2] ~^ image[11][20] + kernel[0][3] ~^ image[11][21] + kernel[0][4] ~^ image[11][22] + kernel[1][0] ~^ image[12][18] + kernel[1][1] ~^ image[12][19] + kernel[1][2] ~^ image[12][20] + kernel[1][3] ~^ image[12][21] + kernel[1][4] ~^ image[12][22] + kernel[2][0] ~^ image[13][18] + kernel[2][1] ~^ image[13][19] + kernel[2][2] ~^ image[13][20] + kernel[2][3] ~^ image[13][21] + kernel[2][4] ~^ image[13][22] + kernel[3][0] ~^ image[14][18] + kernel[3][1] ~^ image[14][19] + kernel[3][2] ~^ image[14][20] + kernel[3][3] ~^ image[14][21] + kernel[3][4] ~^ image[14][22] + kernel[4][0] ~^ image[15][18] + kernel[4][1] ~^ image[15][19] + kernel[4][2] ~^ image[15][20] + kernel[4][3] ~^ image[15][21] + kernel[4][4] ~^ image[15][22];
assign xor_sum[11][19] = kernel[0][0] ~^ image[11][19] + kernel[0][1] ~^ image[11][20] + kernel[0][2] ~^ image[11][21] + kernel[0][3] ~^ image[11][22] + kernel[0][4] ~^ image[11][23] + kernel[1][0] ~^ image[12][19] + kernel[1][1] ~^ image[12][20] + kernel[1][2] ~^ image[12][21] + kernel[1][3] ~^ image[12][22] + kernel[1][4] ~^ image[12][23] + kernel[2][0] ~^ image[13][19] + kernel[2][1] ~^ image[13][20] + kernel[2][2] ~^ image[13][21] + kernel[2][3] ~^ image[13][22] + kernel[2][4] ~^ image[13][23] + kernel[3][0] ~^ image[14][19] + kernel[3][1] ~^ image[14][20] + kernel[3][2] ~^ image[14][21] + kernel[3][3] ~^ image[14][22] + kernel[3][4] ~^ image[14][23] + kernel[4][0] ~^ image[15][19] + kernel[4][1] ~^ image[15][20] + kernel[4][2] ~^ image[15][21] + kernel[4][3] ~^ image[15][22] + kernel[4][4] ~^ image[15][23];
assign xor_sum[11][20] = kernel[0][0] ~^ image[11][20] + kernel[0][1] ~^ image[11][21] + kernel[0][2] ~^ image[11][22] + kernel[0][3] ~^ image[11][23] + kernel[0][4] ~^ image[11][24] + kernel[1][0] ~^ image[12][20] + kernel[1][1] ~^ image[12][21] + kernel[1][2] ~^ image[12][22] + kernel[1][3] ~^ image[12][23] + kernel[1][4] ~^ image[12][24] + kernel[2][0] ~^ image[13][20] + kernel[2][1] ~^ image[13][21] + kernel[2][2] ~^ image[13][22] + kernel[2][3] ~^ image[13][23] + kernel[2][4] ~^ image[13][24] + kernel[3][0] ~^ image[14][20] + kernel[3][1] ~^ image[14][21] + kernel[3][2] ~^ image[14][22] + kernel[3][3] ~^ image[14][23] + kernel[3][4] ~^ image[14][24] + kernel[4][0] ~^ image[15][20] + kernel[4][1] ~^ image[15][21] + kernel[4][2] ~^ image[15][22] + kernel[4][3] ~^ image[15][23] + kernel[4][4] ~^ image[15][24];
assign xor_sum[11][21] = kernel[0][0] ~^ image[11][21] + kernel[0][1] ~^ image[11][22] + kernel[0][2] ~^ image[11][23] + kernel[0][3] ~^ image[11][24] + kernel[0][4] ~^ image[11][25] + kernel[1][0] ~^ image[12][21] + kernel[1][1] ~^ image[12][22] + kernel[1][2] ~^ image[12][23] + kernel[1][3] ~^ image[12][24] + kernel[1][4] ~^ image[12][25] + kernel[2][0] ~^ image[13][21] + kernel[2][1] ~^ image[13][22] + kernel[2][2] ~^ image[13][23] + kernel[2][3] ~^ image[13][24] + kernel[2][4] ~^ image[13][25] + kernel[3][0] ~^ image[14][21] + kernel[3][1] ~^ image[14][22] + kernel[3][2] ~^ image[14][23] + kernel[3][3] ~^ image[14][24] + kernel[3][4] ~^ image[14][25] + kernel[4][0] ~^ image[15][21] + kernel[4][1] ~^ image[15][22] + kernel[4][2] ~^ image[15][23] + kernel[4][3] ~^ image[15][24] + kernel[4][4] ~^ image[15][25];
assign xor_sum[11][22] = kernel[0][0] ~^ image[11][22] + kernel[0][1] ~^ image[11][23] + kernel[0][2] ~^ image[11][24] + kernel[0][3] ~^ image[11][25] + kernel[0][4] ~^ image[11][26] + kernel[1][0] ~^ image[12][22] + kernel[1][1] ~^ image[12][23] + kernel[1][2] ~^ image[12][24] + kernel[1][3] ~^ image[12][25] + kernel[1][4] ~^ image[12][26] + kernel[2][0] ~^ image[13][22] + kernel[2][1] ~^ image[13][23] + kernel[2][2] ~^ image[13][24] + kernel[2][3] ~^ image[13][25] + kernel[2][4] ~^ image[13][26] + kernel[3][0] ~^ image[14][22] + kernel[3][1] ~^ image[14][23] + kernel[3][2] ~^ image[14][24] + kernel[3][3] ~^ image[14][25] + kernel[3][4] ~^ image[14][26] + kernel[4][0] ~^ image[15][22] + kernel[4][1] ~^ image[15][23] + kernel[4][2] ~^ image[15][24] + kernel[4][3] ~^ image[15][25] + kernel[4][4] ~^ image[15][26];
assign xor_sum[11][23] = kernel[0][0] ~^ image[11][23] + kernel[0][1] ~^ image[11][24] + kernel[0][2] ~^ image[11][25] + kernel[0][3] ~^ image[11][26] + kernel[0][4] ~^ image[11][27] + kernel[1][0] ~^ image[12][23] + kernel[1][1] ~^ image[12][24] + kernel[1][2] ~^ image[12][25] + kernel[1][3] ~^ image[12][26] + kernel[1][4] ~^ image[12][27] + kernel[2][0] ~^ image[13][23] + kernel[2][1] ~^ image[13][24] + kernel[2][2] ~^ image[13][25] + kernel[2][3] ~^ image[13][26] + kernel[2][4] ~^ image[13][27] + kernel[3][0] ~^ image[14][23] + kernel[3][1] ~^ image[14][24] + kernel[3][2] ~^ image[14][25] + kernel[3][3] ~^ image[14][26] + kernel[3][4] ~^ image[14][27] + kernel[4][0] ~^ image[15][23] + kernel[4][1] ~^ image[15][24] + kernel[4][2] ~^ image[15][25] + kernel[4][3] ~^ image[15][26] + kernel[4][4] ~^ image[15][27];
assign xor_sum[12][0] = kernel[0][0] ~^ image[12][0] + kernel[0][1] ~^ image[12][1] + kernel[0][2] ~^ image[12][2] + kernel[0][3] ~^ image[12][3] + kernel[0][4] ~^ image[12][4] + kernel[1][0] ~^ image[13][0] + kernel[1][1] ~^ image[13][1] + kernel[1][2] ~^ image[13][2] + kernel[1][3] ~^ image[13][3] + kernel[1][4] ~^ image[13][4] + kernel[2][0] ~^ image[14][0] + kernel[2][1] ~^ image[14][1] + kernel[2][2] ~^ image[14][2] + kernel[2][3] ~^ image[14][3] + kernel[2][4] ~^ image[14][4] + kernel[3][0] ~^ image[15][0] + kernel[3][1] ~^ image[15][1] + kernel[3][2] ~^ image[15][2] + kernel[3][3] ~^ image[15][3] + kernel[3][4] ~^ image[15][4] + kernel[4][0] ~^ image[16][0] + kernel[4][1] ~^ image[16][1] + kernel[4][2] ~^ image[16][2] + kernel[4][3] ~^ image[16][3] + kernel[4][4] ~^ image[16][4];
assign xor_sum[12][1] = kernel[0][0] ~^ image[12][1] + kernel[0][1] ~^ image[12][2] + kernel[0][2] ~^ image[12][3] + kernel[0][3] ~^ image[12][4] + kernel[0][4] ~^ image[12][5] + kernel[1][0] ~^ image[13][1] + kernel[1][1] ~^ image[13][2] + kernel[1][2] ~^ image[13][3] + kernel[1][3] ~^ image[13][4] + kernel[1][4] ~^ image[13][5] + kernel[2][0] ~^ image[14][1] + kernel[2][1] ~^ image[14][2] + kernel[2][2] ~^ image[14][3] + kernel[2][3] ~^ image[14][4] + kernel[2][4] ~^ image[14][5] + kernel[3][0] ~^ image[15][1] + kernel[3][1] ~^ image[15][2] + kernel[3][2] ~^ image[15][3] + kernel[3][3] ~^ image[15][4] + kernel[3][4] ~^ image[15][5] + kernel[4][0] ~^ image[16][1] + kernel[4][1] ~^ image[16][2] + kernel[4][2] ~^ image[16][3] + kernel[4][3] ~^ image[16][4] + kernel[4][4] ~^ image[16][5];
assign xor_sum[12][2] = kernel[0][0] ~^ image[12][2] + kernel[0][1] ~^ image[12][3] + kernel[0][2] ~^ image[12][4] + kernel[0][3] ~^ image[12][5] + kernel[0][4] ~^ image[12][6] + kernel[1][0] ~^ image[13][2] + kernel[1][1] ~^ image[13][3] + kernel[1][2] ~^ image[13][4] + kernel[1][3] ~^ image[13][5] + kernel[1][4] ~^ image[13][6] + kernel[2][0] ~^ image[14][2] + kernel[2][1] ~^ image[14][3] + kernel[2][2] ~^ image[14][4] + kernel[2][3] ~^ image[14][5] + kernel[2][4] ~^ image[14][6] + kernel[3][0] ~^ image[15][2] + kernel[3][1] ~^ image[15][3] + kernel[3][2] ~^ image[15][4] + kernel[3][3] ~^ image[15][5] + kernel[3][4] ~^ image[15][6] + kernel[4][0] ~^ image[16][2] + kernel[4][1] ~^ image[16][3] + kernel[4][2] ~^ image[16][4] + kernel[4][3] ~^ image[16][5] + kernel[4][4] ~^ image[16][6];
assign xor_sum[12][3] = kernel[0][0] ~^ image[12][3] + kernel[0][1] ~^ image[12][4] + kernel[0][2] ~^ image[12][5] + kernel[0][3] ~^ image[12][6] + kernel[0][4] ~^ image[12][7] + kernel[1][0] ~^ image[13][3] + kernel[1][1] ~^ image[13][4] + kernel[1][2] ~^ image[13][5] + kernel[1][3] ~^ image[13][6] + kernel[1][4] ~^ image[13][7] + kernel[2][0] ~^ image[14][3] + kernel[2][1] ~^ image[14][4] + kernel[2][2] ~^ image[14][5] + kernel[2][3] ~^ image[14][6] + kernel[2][4] ~^ image[14][7] + kernel[3][0] ~^ image[15][3] + kernel[3][1] ~^ image[15][4] + kernel[3][2] ~^ image[15][5] + kernel[3][3] ~^ image[15][6] + kernel[3][4] ~^ image[15][7] + kernel[4][0] ~^ image[16][3] + kernel[4][1] ~^ image[16][4] + kernel[4][2] ~^ image[16][5] + kernel[4][3] ~^ image[16][6] + kernel[4][4] ~^ image[16][7];
assign xor_sum[12][4] = kernel[0][0] ~^ image[12][4] + kernel[0][1] ~^ image[12][5] + kernel[0][2] ~^ image[12][6] + kernel[0][3] ~^ image[12][7] + kernel[0][4] ~^ image[12][8] + kernel[1][0] ~^ image[13][4] + kernel[1][1] ~^ image[13][5] + kernel[1][2] ~^ image[13][6] + kernel[1][3] ~^ image[13][7] + kernel[1][4] ~^ image[13][8] + kernel[2][0] ~^ image[14][4] + kernel[2][1] ~^ image[14][5] + kernel[2][2] ~^ image[14][6] + kernel[2][3] ~^ image[14][7] + kernel[2][4] ~^ image[14][8] + kernel[3][0] ~^ image[15][4] + kernel[3][1] ~^ image[15][5] + kernel[3][2] ~^ image[15][6] + kernel[3][3] ~^ image[15][7] + kernel[3][4] ~^ image[15][8] + kernel[4][0] ~^ image[16][4] + kernel[4][1] ~^ image[16][5] + kernel[4][2] ~^ image[16][6] + kernel[4][3] ~^ image[16][7] + kernel[4][4] ~^ image[16][8];
assign xor_sum[12][5] = kernel[0][0] ~^ image[12][5] + kernel[0][1] ~^ image[12][6] + kernel[0][2] ~^ image[12][7] + kernel[0][3] ~^ image[12][8] + kernel[0][4] ~^ image[12][9] + kernel[1][0] ~^ image[13][5] + kernel[1][1] ~^ image[13][6] + kernel[1][2] ~^ image[13][7] + kernel[1][3] ~^ image[13][8] + kernel[1][4] ~^ image[13][9] + kernel[2][0] ~^ image[14][5] + kernel[2][1] ~^ image[14][6] + kernel[2][2] ~^ image[14][7] + kernel[2][3] ~^ image[14][8] + kernel[2][4] ~^ image[14][9] + kernel[3][0] ~^ image[15][5] + kernel[3][1] ~^ image[15][6] + kernel[3][2] ~^ image[15][7] + kernel[3][3] ~^ image[15][8] + kernel[3][4] ~^ image[15][9] + kernel[4][0] ~^ image[16][5] + kernel[4][1] ~^ image[16][6] + kernel[4][2] ~^ image[16][7] + kernel[4][3] ~^ image[16][8] + kernel[4][4] ~^ image[16][9];
assign xor_sum[12][6] = kernel[0][0] ~^ image[12][6] + kernel[0][1] ~^ image[12][7] + kernel[0][2] ~^ image[12][8] + kernel[0][3] ~^ image[12][9] + kernel[0][4] ~^ image[12][10] + kernel[1][0] ~^ image[13][6] + kernel[1][1] ~^ image[13][7] + kernel[1][2] ~^ image[13][8] + kernel[1][3] ~^ image[13][9] + kernel[1][4] ~^ image[13][10] + kernel[2][0] ~^ image[14][6] + kernel[2][1] ~^ image[14][7] + kernel[2][2] ~^ image[14][8] + kernel[2][3] ~^ image[14][9] + kernel[2][4] ~^ image[14][10] + kernel[3][0] ~^ image[15][6] + kernel[3][1] ~^ image[15][7] + kernel[3][2] ~^ image[15][8] + kernel[3][3] ~^ image[15][9] + kernel[3][4] ~^ image[15][10] + kernel[4][0] ~^ image[16][6] + kernel[4][1] ~^ image[16][7] + kernel[4][2] ~^ image[16][8] + kernel[4][3] ~^ image[16][9] + kernel[4][4] ~^ image[16][10];
assign xor_sum[12][7] = kernel[0][0] ~^ image[12][7] + kernel[0][1] ~^ image[12][8] + kernel[0][2] ~^ image[12][9] + kernel[0][3] ~^ image[12][10] + kernel[0][4] ~^ image[12][11] + kernel[1][0] ~^ image[13][7] + kernel[1][1] ~^ image[13][8] + kernel[1][2] ~^ image[13][9] + kernel[1][3] ~^ image[13][10] + kernel[1][4] ~^ image[13][11] + kernel[2][0] ~^ image[14][7] + kernel[2][1] ~^ image[14][8] + kernel[2][2] ~^ image[14][9] + kernel[2][3] ~^ image[14][10] + kernel[2][4] ~^ image[14][11] + kernel[3][0] ~^ image[15][7] + kernel[3][1] ~^ image[15][8] + kernel[3][2] ~^ image[15][9] + kernel[3][3] ~^ image[15][10] + kernel[3][4] ~^ image[15][11] + kernel[4][0] ~^ image[16][7] + kernel[4][1] ~^ image[16][8] + kernel[4][2] ~^ image[16][9] + kernel[4][3] ~^ image[16][10] + kernel[4][4] ~^ image[16][11];
assign xor_sum[12][8] = kernel[0][0] ~^ image[12][8] + kernel[0][1] ~^ image[12][9] + kernel[0][2] ~^ image[12][10] + kernel[0][3] ~^ image[12][11] + kernel[0][4] ~^ image[12][12] + kernel[1][0] ~^ image[13][8] + kernel[1][1] ~^ image[13][9] + kernel[1][2] ~^ image[13][10] + kernel[1][3] ~^ image[13][11] + kernel[1][4] ~^ image[13][12] + kernel[2][0] ~^ image[14][8] + kernel[2][1] ~^ image[14][9] + kernel[2][2] ~^ image[14][10] + kernel[2][3] ~^ image[14][11] + kernel[2][4] ~^ image[14][12] + kernel[3][0] ~^ image[15][8] + kernel[3][1] ~^ image[15][9] + kernel[3][2] ~^ image[15][10] + kernel[3][3] ~^ image[15][11] + kernel[3][4] ~^ image[15][12] + kernel[4][0] ~^ image[16][8] + kernel[4][1] ~^ image[16][9] + kernel[4][2] ~^ image[16][10] + kernel[4][3] ~^ image[16][11] + kernel[4][4] ~^ image[16][12];
assign xor_sum[12][9] = kernel[0][0] ~^ image[12][9] + kernel[0][1] ~^ image[12][10] + kernel[0][2] ~^ image[12][11] + kernel[0][3] ~^ image[12][12] + kernel[0][4] ~^ image[12][13] + kernel[1][0] ~^ image[13][9] + kernel[1][1] ~^ image[13][10] + kernel[1][2] ~^ image[13][11] + kernel[1][3] ~^ image[13][12] + kernel[1][4] ~^ image[13][13] + kernel[2][0] ~^ image[14][9] + kernel[2][1] ~^ image[14][10] + kernel[2][2] ~^ image[14][11] + kernel[2][3] ~^ image[14][12] + kernel[2][4] ~^ image[14][13] + kernel[3][0] ~^ image[15][9] + kernel[3][1] ~^ image[15][10] + kernel[3][2] ~^ image[15][11] + kernel[3][3] ~^ image[15][12] + kernel[3][4] ~^ image[15][13] + kernel[4][0] ~^ image[16][9] + kernel[4][1] ~^ image[16][10] + kernel[4][2] ~^ image[16][11] + kernel[4][3] ~^ image[16][12] + kernel[4][4] ~^ image[16][13];
assign xor_sum[12][10] = kernel[0][0] ~^ image[12][10] + kernel[0][1] ~^ image[12][11] + kernel[0][2] ~^ image[12][12] + kernel[0][3] ~^ image[12][13] + kernel[0][4] ~^ image[12][14] + kernel[1][0] ~^ image[13][10] + kernel[1][1] ~^ image[13][11] + kernel[1][2] ~^ image[13][12] + kernel[1][3] ~^ image[13][13] + kernel[1][4] ~^ image[13][14] + kernel[2][0] ~^ image[14][10] + kernel[2][1] ~^ image[14][11] + kernel[2][2] ~^ image[14][12] + kernel[2][3] ~^ image[14][13] + kernel[2][4] ~^ image[14][14] + kernel[3][0] ~^ image[15][10] + kernel[3][1] ~^ image[15][11] + kernel[3][2] ~^ image[15][12] + kernel[3][3] ~^ image[15][13] + kernel[3][4] ~^ image[15][14] + kernel[4][0] ~^ image[16][10] + kernel[4][1] ~^ image[16][11] + kernel[4][2] ~^ image[16][12] + kernel[4][3] ~^ image[16][13] + kernel[4][4] ~^ image[16][14];
assign xor_sum[12][11] = kernel[0][0] ~^ image[12][11] + kernel[0][1] ~^ image[12][12] + kernel[0][2] ~^ image[12][13] + kernel[0][3] ~^ image[12][14] + kernel[0][4] ~^ image[12][15] + kernel[1][0] ~^ image[13][11] + kernel[1][1] ~^ image[13][12] + kernel[1][2] ~^ image[13][13] + kernel[1][3] ~^ image[13][14] + kernel[1][4] ~^ image[13][15] + kernel[2][0] ~^ image[14][11] + kernel[2][1] ~^ image[14][12] + kernel[2][2] ~^ image[14][13] + kernel[2][3] ~^ image[14][14] + kernel[2][4] ~^ image[14][15] + kernel[3][0] ~^ image[15][11] + kernel[3][1] ~^ image[15][12] + kernel[3][2] ~^ image[15][13] + kernel[3][3] ~^ image[15][14] + kernel[3][4] ~^ image[15][15] + kernel[4][0] ~^ image[16][11] + kernel[4][1] ~^ image[16][12] + kernel[4][2] ~^ image[16][13] + kernel[4][3] ~^ image[16][14] + kernel[4][4] ~^ image[16][15];
assign xor_sum[12][12] = kernel[0][0] ~^ image[12][12] + kernel[0][1] ~^ image[12][13] + kernel[0][2] ~^ image[12][14] + kernel[0][3] ~^ image[12][15] + kernel[0][4] ~^ image[12][16] + kernel[1][0] ~^ image[13][12] + kernel[1][1] ~^ image[13][13] + kernel[1][2] ~^ image[13][14] + kernel[1][3] ~^ image[13][15] + kernel[1][4] ~^ image[13][16] + kernel[2][0] ~^ image[14][12] + kernel[2][1] ~^ image[14][13] + kernel[2][2] ~^ image[14][14] + kernel[2][3] ~^ image[14][15] + kernel[2][4] ~^ image[14][16] + kernel[3][0] ~^ image[15][12] + kernel[3][1] ~^ image[15][13] + kernel[3][2] ~^ image[15][14] + kernel[3][3] ~^ image[15][15] + kernel[3][4] ~^ image[15][16] + kernel[4][0] ~^ image[16][12] + kernel[4][1] ~^ image[16][13] + kernel[4][2] ~^ image[16][14] + kernel[4][3] ~^ image[16][15] + kernel[4][4] ~^ image[16][16];
assign xor_sum[12][13] = kernel[0][0] ~^ image[12][13] + kernel[0][1] ~^ image[12][14] + kernel[0][2] ~^ image[12][15] + kernel[0][3] ~^ image[12][16] + kernel[0][4] ~^ image[12][17] + kernel[1][0] ~^ image[13][13] + kernel[1][1] ~^ image[13][14] + kernel[1][2] ~^ image[13][15] + kernel[1][3] ~^ image[13][16] + kernel[1][4] ~^ image[13][17] + kernel[2][0] ~^ image[14][13] + kernel[2][1] ~^ image[14][14] + kernel[2][2] ~^ image[14][15] + kernel[2][3] ~^ image[14][16] + kernel[2][4] ~^ image[14][17] + kernel[3][0] ~^ image[15][13] + kernel[3][1] ~^ image[15][14] + kernel[3][2] ~^ image[15][15] + kernel[3][3] ~^ image[15][16] + kernel[3][4] ~^ image[15][17] + kernel[4][0] ~^ image[16][13] + kernel[4][1] ~^ image[16][14] + kernel[4][2] ~^ image[16][15] + kernel[4][3] ~^ image[16][16] + kernel[4][4] ~^ image[16][17];
assign xor_sum[12][14] = kernel[0][0] ~^ image[12][14] + kernel[0][1] ~^ image[12][15] + kernel[0][2] ~^ image[12][16] + kernel[0][3] ~^ image[12][17] + kernel[0][4] ~^ image[12][18] + kernel[1][0] ~^ image[13][14] + kernel[1][1] ~^ image[13][15] + kernel[1][2] ~^ image[13][16] + kernel[1][3] ~^ image[13][17] + kernel[1][4] ~^ image[13][18] + kernel[2][0] ~^ image[14][14] + kernel[2][1] ~^ image[14][15] + kernel[2][2] ~^ image[14][16] + kernel[2][3] ~^ image[14][17] + kernel[2][4] ~^ image[14][18] + kernel[3][0] ~^ image[15][14] + kernel[3][1] ~^ image[15][15] + kernel[3][2] ~^ image[15][16] + kernel[3][3] ~^ image[15][17] + kernel[3][4] ~^ image[15][18] + kernel[4][0] ~^ image[16][14] + kernel[4][1] ~^ image[16][15] + kernel[4][2] ~^ image[16][16] + kernel[4][3] ~^ image[16][17] + kernel[4][4] ~^ image[16][18];
assign xor_sum[12][15] = kernel[0][0] ~^ image[12][15] + kernel[0][1] ~^ image[12][16] + kernel[0][2] ~^ image[12][17] + kernel[0][3] ~^ image[12][18] + kernel[0][4] ~^ image[12][19] + kernel[1][0] ~^ image[13][15] + kernel[1][1] ~^ image[13][16] + kernel[1][2] ~^ image[13][17] + kernel[1][3] ~^ image[13][18] + kernel[1][4] ~^ image[13][19] + kernel[2][0] ~^ image[14][15] + kernel[2][1] ~^ image[14][16] + kernel[2][2] ~^ image[14][17] + kernel[2][3] ~^ image[14][18] + kernel[2][4] ~^ image[14][19] + kernel[3][0] ~^ image[15][15] + kernel[3][1] ~^ image[15][16] + kernel[3][2] ~^ image[15][17] + kernel[3][3] ~^ image[15][18] + kernel[3][4] ~^ image[15][19] + kernel[4][0] ~^ image[16][15] + kernel[4][1] ~^ image[16][16] + kernel[4][2] ~^ image[16][17] + kernel[4][3] ~^ image[16][18] + kernel[4][4] ~^ image[16][19];
assign xor_sum[12][16] = kernel[0][0] ~^ image[12][16] + kernel[0][1] ~^ image[12][17] + kernel[0][2] ~^ image[12][18] + kernel[0][3] ~^ image[12][19] + kernel[0][4] ~^ image[12][20] + kernel[1][0] ~^ image[13][16] + kernel[1][1] ~^ image[13][17] + kernel[1][2] ~^ image[13][18] + kernel[1][3] ~^ image[13][19] + kernel[1][4] ~^ image[13][20] + kernel[2][0] ~^ image[14][16] + kernel[2][1] ~^ image[14][17] + kernel[2][2] ~^ image[14][18] + kernel[2][3] ~^ image[14][19] + kernel[2][4] ~^ image[14][20] + kernel[3][0] ~^ image[15][16] + kernel[3][1] ~^ image[15][17] + kernel[3][2] ~^ image[15][18] + kernel[3][3] ~^ image[15][19] + kernel[3][4] ~^ image[15][20] + kernel[4][0] ~^ image[16][16] + kernel[4][1] ~^ image[16][17] + kernel[4][2] ~^ image[16][18] + kernel[4][3] ~^ image[16][19] + kernel[4][4] ~^ image[16][20];
assign xor_sum[12][17] = kernel[0][0] ~^ image[12][17] + kernel[0][1] ~^ image[12][18] + kernel[0][2] ~^ image[12][19] + kernel[0][3] ~^ image[12][20] + kernel[0][4] ~^ image[12][21] + kernel[1][0] ~^ image[13][17] + kernel[1][1] ~^ image[13][18] + kernel[1][2] ~^ image[13][19] + kernel[1][3] ~^ image[13][20] + kernel[1][4] ~^ image[13][21] + kernel[2][0] ~^ image[14][17] + kernel[2][1] ~^ image[14][18] + kernel[2][2] ~^ image[14][19] + kernel[2][3] ~^ image[14][20] + kernel[2][4] ~^ image[14][21] + kernel[3][0] ~^ image[15][17] + kernel[3][1] ~^ image[15][18] + kernel[3][2] ~^ image[15][19] + kernel[3][3] ~^ image[15][20] + kernel[3][4] ~^ image[15][21] + kernel[4][0] ~^ image[16][17] + kernel[4][1] ~^ image[16][18] + kernel[4][2] ~^ image[16][19] + kernel[4][3] ~^ image[16][20] + kernel[4][4] ~^ image[16][21];
assign xor_sum[12][18] = kernel[0][0] ~^ image[12][18] + kernel[0][1] ~^ image[12][19] + kernel[0][2] ~^ image[12][20] + kernel[0][3] ~^ image[12][21] + kernel[0][4] ~^ image[12][22] + kernel[1][0] ~^ image[13][18] + kernel[1][1] ~^ image[13][19] + kernel[1][2] ~^ image[13][20] + kernel[1][3] ~^ image[13][21] + kernel[1][4] ~^ image[13][22] + kernel[2][0] ~^ image[14][18] + kernel[2][1] ~^ image[14][19] + kernel[2][2] ~^ image[14][20] + kernel[2][3] ~^ image[14][21] + kernel[2][4] ~^ image[14][22] + kernel[3][0] ~^ image[15][18] + kernel[3][1] ~^ image[15][19] + kernel[3][2] ~^ image[15][20] + kernel[3][3] ~^ image[15][21] + kernel[3][4] ~^ image[15][22] + kernel[4][0] ~^ image[16][18] + kernel[4][1] ~^ image[16][19] + kernel[4][2] ~^ image[16][20] + kernel[4][3] ~^ image[16][21] + kernel[4][4] ~^ image[16][22];
assign xor_sum[12][19] = kernel[0][0] ~^ image[12][19] + kernel[0][1] ~^ image[12][20] + kernel[0][2] ~^ image[12][21] + kernel[0][3] ~^ image[12][22] + kernel[0][4] ~^ image[12][23] + kernel[1][0] ~^ image[13][19] + kernel[1][1] ~^ image[13][20] + kernel[1][2] ~^ image[13][21] + kernel[1][3] ~^ image[13][22] + kernel[1][4] ~^ image[13][23] + kernel[2][0] ~^ image[14][19] + kernel[2][1] ~^ image[14][20] + kernel[2][2] ~^ image[14][21] + kernel[2][3] ~^ image[14][22] + kernel[2][4] ~^ image[14][23] + kernel[3][0] ~^ image[15][19] + kernel[3][1] ~^ image[15][20] + kernel[3][2] ~^ image[15][21] + kernel[3][3] ~^ image[15][22] + kernel[3][4] ~^ image[15][23] + kernel[4][0] ~^ image[16][19] + kernel[4][1] ~^ image[16][20] + kernel[4][2] ~^ image[16][21] + kernel[4][3] ~^ image[16][22] + kernel[4][4] ~^ image[16][23];
assign xor_sum[12][20] = kernel[0][0] ~^ image[12][20] + kernel[0][1] ~^ image[12][21] + kernel[0][2] ~^ image[12][22] + kernel[0][3] ~^ image[12][23] + kernel[0][4] ~^ image[12][24] + kernel[1][0] ~^ image[13][20] + kernel[1][1] ~^ image[13][21] + kernel[1][2] ~^ image[13][22] + kernel[1][3] ~^ image[13][23] + kernel[1][4] ~^ image[13][24] + kernel[2][0] ~^ image[14][20] + kernel[2][1] ~^ image[14][21] + kernel[2][2] ~^ image[14][22] + kernel[2][3] ~^ image[14][23] + kernel[2][4] ~^ image[14][24] + kernel[3][0] ~^ image[15][20] + kernel[3][1] ~^ image[15][21] + kernel[3][2] ~^ image[15][22] + kernel[3][3] ~^ image[15][23] + kernel[3][4] ~^ image[15][24] + kernel[4][0] ~^ image[16][20] + kernel[4][1] ~^ image[16][21] + kernel[4][2] ~^ image[16][22] + kernel[4][3] ~^ image[16][23] + kernel[4][4] ~^ image[16][24];
assign xor_sum[12][21] = kernel[0][0] ~^ image[12][21] + kernel[0][1] ~^ image[12][22] + kernel[0][2] ~^ image[12][23] + kernel[0][3] ~^ image[12][24] + kernel[0][4] ~^ image[12][25] + kernel[1][0] ~^ image[13][21] + kernel[1][1] ~^ image[13][22] + kernel[1][2] ~^ image[13][23] + kernel[1][3] ~^ image[13][24] + kernel[1][4] ~^ image[13][25] + kernel[2][0] ~^ image[14][21] + kernel[2][1] ~^ image[14][22] + kernel[2][2] ~^ image[14][23] + kernel[2][3] ~^ image[14][24] + kernel[2][4] ~^ image[14][25] + kernel[3][0] ~^ image[15][21] + kernel[3][1] ~^ image[15][22] + kernel[3][2] ~^ image[15][23] + kernel[3][3] ~^ image[15][24] + kernel[3][4] ~^ image[15][25] + kernel[4][0] ~^ image[16][21] + kernel[4][1] ~^ image[16][22] + kernel[4][2] ~^ image[16][23] + kernel[4][3] ~^ image[16][24] + kernel[4][4] ~^ image[16][25];
assign xor_sum[12][22] = kernel[0][0] ~^ image[12][22] + kernel[0][1] ~^ image[12][23] + kernel[0][2] ~^ image[12][24] + kernel[0][3] ~^ image[12][25] + kernel[0][4] ~^ image[12][26] + kernel[1][0] ~^ image[13][22] + kernel[1][1] ~^ image[13][23] + kernel[1][2] ~^ image[13][24] + kernel[1][3] ~^ image[13][25] + kernel[1][4] ~^ image[13][26] + kernel[2][0] ~^ image[14][22] + kernel[2][1] ~^ image[14][23] + kernel[2][2] ~^ image[14][24] + kernel[2][3] ~^ image[14][25] + kernel[2][4] ~^ image[14][26] + kernel[3][0] ~^ image[15][22] + kernel[3][1] ~^ image[15][23] + kernel[3][2] ~^ image[15][24] + kernel[3][3] ~^ image[15][25] + kernel[3][4] ~^ image[15][26] + kernel[4][0] ~^ image[16][22] + kernel[4][1] ~^ image[16][23] + kernel[4][2] ~^ image[16][24] + kernel[4][3] ~^ image[16][25] + kernel[4][4] ~^ image[16][26];
assign xor_sum[12][23] = kernel[0][0] ~^ image[12][23] + kernel[0][1] ~^ image[12][24] + kernel[0][2] ~^ image[12][25] + kernel[0][3] ~^ image[12][26] + kernel[0][4] ~^ image[12][27] + kernel[1][0] ~^ image[13][23] + kernel[1][1] ~^ image[13][24] + kernel[1][2] ~^ image[13][25] + kernel[1][3] ~^ image[13][26] + kernel[1][4] ~^ image[13][27] + kernel[2][0] ~^ image[14][23] + kernel[2][1] ~^ image[14][24] + kernel[2][2] ~^ image[14][25] + kernel[2][3] ~^ image[14][26] + kernel[2][4] ~^ image[14][27] + kernel[3][0] ~^ image[15][23] + kernel[3][1] ~^ image[15][24] + kernel[3][2] ~^ image[15][25] + kernel[3][3] ~^ image[15][26] + kernel[3][4] ~^ image[15][27] + kernel[4][0] ~^ image[16][23] + kernel[4][1] ~^ image[16][24] + kernel[4][2] ~^ image[16][25] + kernel[4][3] ~^ image[16][26] + kernel[4][4] ~^ image[16][27];
assign xor_sum[13][0] = kernel[0][0] ~^ image[13][0] + kernel[0][1] ~^ image[13][1] + kernel[0][2] ~^ image[13][2] + kernel[0][3] ~^ image[13][3] + kernel[0][4] ~^ image[13][4] + kernel[1][0] ~^ image[14][0] + kernel[1][1] ~^ image[14][1] + kernel[1][2] ~^ image[14][2] + kernel[1][3] ~^ image[14][3] + kernel[1][4] ~^ image[14][4] + kernel[2][0] ~^ image[15][0] + kernel[2][1] ~^ image[15][1] + kernel[2][2] ~^ image[15][2] + kernel[2][3] ~^ image[15][3] + kernel[2][4] ~^ image[15][4] + kernel[3][0] ~^ image[16][0] + kernel[3][1] ~^ image[16][1] + kernel[3][2] ~^ image[16][2] + kernel[3][3] ~^ image[16][3] + kernel[3][4] ~^ image[16][4] + kernel[4][0] ~^ image[17][0] + kernel[4][1] ~^ image[17][1] + kernel[4][2] ~^ image[17][2] + kernel[4][3] ~^ image[17][3] + kernel[4][4] ~^ image[17][4];
assign xor_sum[13][1] = kernel[0][0] ~^ image[13][1] + kernel[0][1] ~^ image[13][2] + kernel[0][2] ~^ image[13][3] + kernel[0][3] ~^ image[13][4] + kernel[0][4] ~^ image[13][5] + kernel[1][0] ~^ image[14][1] + kernel[1][1] ~^ image[14][2] + kernel[1][2] ~^ image[14][3] + kernel[1][3] ~^ image[14][4] + kernel[1][4] ~^ image[14][5] + kernel[2][0] ~^ image[15][1] + kernel[2][1] ~^ image[15][2] + kernel[2][2] ~^ image[15][3] + kernel[2][3] ~^ image[15][4] + kernel[2][4] ~^ image[15][5] + kernel[3][0] ~^ image[16][1] + kernel[3][1] ~^ image[16][2] + kernel[3][2] ~^ image[16][3] + kernel[3][3] ~^ image[16][4] + kernel[3][4] ~^ image[16][5] + kernel[4][0] ~^ image[17][1] + kernel[4][1] ~^ image[17][2] + kernel[4][2] ~^ image[17][3] + kernel[4][3] ~^ image[17][4] + kernel[4][4] ~^ image[17][5];
assign xor_sum[13][2] = kernel[0][0] ~^ image[13][2] + kernel[0][1] ~^ image[13][3] + kernel[0][2] ~^ image[13][4] + kernel[0][3] ~^ image[13][5] + kernel[0][4] ~^ image[13][6] + kernel[1][0] ~^ image[14][2] + kernel[1][1] ~^ image[14][3] + kernel[1][2] ~^ image[14][4] + kernel[1][3] ~^ image[14][5] + kernel[1][4] ~^ image[14][6] + kernel[2][0] ~^ image[15][2] + kernel[2][1] ~^ image[15][3] + kernel[2][2] ~^ image[15][4] + kernel[2][3] ~^ image[15][5] + kernel[2][4] ~^ image[15][6] + kernel[3][0] ~^ image[16][2] + kernel[3][1] ~^ image[16][3] + kernel[3][2] ~^ image[16][4] + kernel[3][3] ~^ image[16][5] + kernel[3][4] ~^ image[16][6] + kernel[4][0] ~^ image[17][2] + kernel[4][1] ~^ image[17][3] + kernel[4][2] ~^ image[17][4] + kernel[4][3] ~^ image[17][5] + kernel[4][4] ~^ image[17][6];
assign xor_sum[13][3] = kernel[0][0] ~^ image[13][3] + kernel[0][1] ~^ image[13][4] + kernel[0][2] ~^ image[13][5] + kernel[0][3] ~^ image[13][6] + kernel[0][4] ~^ image[13][7] + kernel[1][0] ~^ image[14][3] + kernel[1][1] ~^ image[14][4] + kernel[1][2] ~^ image[14][5] + kernel[1][3] ~^ image[14][6] + kernel[1][4] ~^ image[14][7] + kernel[2][0] ~^ image[15][3] + kernel[2][1] ~^ image[15][4] + kernel[2][2] ~^ image[15][5] + kernel[2][3] ~^ image[15][6] + kernel[2][4] ~^ image[15][7] + kernel[3][0] ~^ image[16][3] + kernel[3][1] ~^ image[16][4] + kernel[3][2] ~^ image[16][5] + kernel[3][3] ~^ image[16][6] + kernel[3][4] ~^ image[16][7] + kernel[4][0] ~^ image[17][3] + kernel[4][1] ~^ image[17][4] + kernel[4][2] ~^ image[17][5] + kernel[4][3] ~^ image[17][6] + kernel[4][4] ~^ image[17][7];
assign xor_sum[13][4] = kernel[0][0] ~^ image[13][4] + kernel[0][1] ~^ image[13][5] + kernel[0][2] ~^ image[13][6] + kernel[0][3] ~^ image[13][7] + kernel[0][4] ~^ image[13][8] + kernel[1][0] ~^ image[14][4] + kernel[1][1] ~^ image[14][5] + kernel[1][2] ~^ image[14][6] + kernel[1][3] ~^ image[14][7] + kernel[1][4] ~^ image[14][8] + kernel[2][0] ~^ image[15][4] + kernel[2][1] ~^ image[15][5] + kernel[2][2] ~^ image[15][6] + kernel[2][3] ~^ image[15][7] + kernel[2][4] ~^ image[15][8] + kernel[3][0] ~^ image[16][4] + kernel[3][1] ~^ image[16][5] + kernel[3][2] ~^ image[16][6] + kernel[3][3] ~^ image[16][7] + kernel[3][4] ~^ image[16][8] + kernel[4][0] ~^ image[17][4] + kernel[4][1] ~^ image[17][5] + kernel[4][2] ~^ image[17][6] + kernel[4][3] ~^ image[17][7] + kernel[4][4] ~^ image[17][8];
assign xor_sum[13][5] = kernel[0][0] ~^ image[13][5] + kernel[0][1] ~^ image[13][6] + kernel[0][2] ~^ image[13][7] + kernel[0][3] ~^ image[13][8] + kernel[0][4] ~^ image[13][9] + kernel[1][0] ~^ image[14][5] + kernel[1][1] ~^ image[14][6] + kernel[1][2] ~^ image[14][7] + kernel[1][3] ~^ image[14][8] + kernel[1][4] ~^ image[14][9] + kernel[2][0] ~^ image[15][5] + kernel[2][1] ~^ image[15][6] + kernel[2][2] ~^ image[15][7] + kernel[2][3] ~^ image[15][8] + kernel[2][4] ~^ image[15][9] + kernel[3][0] ~^ image[16][5] + kernel[3][1] ~^ image[16][6] + kernel[3][2] ~^ image[16][7] + kernel[3][3] ~^ image[16][8] + kernel[3][4] ~^ image[16][9] + kernel[4][0] ~^ image[17][5] + kernel[4][1] ~^ image[17][6] + kernel[4][2] ~^ image[17][7] + kernel[4][3] ~^ image[17][8] + kernel[4][4] ~^ image[17][9];
assign xor_sum[13][6] = kernel[0][0] ~^ image[13][6] + kernel[0][1] ~^ image[13][7] + kernel[0][2] ~^ image[13][8] + kernel[0][3] ~^ image[13][9] + kernel[0][4] ~^ image[13][10] + kernel[1][0] ~^ image[14][6] + kernel[1][1] ~^ image[14][7] + kernel[1][2] ~^ image[14][8] + kernel[1][3] ~^ image[14][9] + kernel[1][4] ~^ image[14][10] + kernel[2][0] ~^ image[15][6] + kernel[2][1] ~^ image[15][7] + kernel[2][2] ~^ image[15][8] + kernel[2][3] ~^ image[15][9] + kernel[2][4] ~^ image[15][10] + kernel[3][0] ~^ image[16][6] + kernel[3][1] ~^ image[16][7] + kernel[3][2] ~^ image[16][8] + kernel[3][3] ~^ image[16][9] + kernel[3][4] ~^ image[16][10] + kernel[4][0] ~^ image[17][6] + kernel[4][1] ~^ image[17][7] + kernel[4][2] ~^ image[17][8] + kernel[4][3] ~^ image[17][9] + kernel[4][4] ~^ image[17][10];
assign xor_sum[13][7] = kernel[0][0] ~^ image[13][7] + kernel[0][1] ~^ image[13][8] + kernel[0][2] ~^ image[13][9] + kernel[0][3] ~^ image[13][10] + kernel[0][4] ~^ image[13][11] + kernel[1][0] ~^ image[14][7] + kernel[1][1] ~^ image[14][8] + kernel[1][2] ~^ image[14][9] + kernel[1][3] ~^ image[14][10] + kernel[1][4] ~^ image[14][11] + kernel[2][0] ~^ image[15][7] + kernel[2][1] ~^ image[15][8] + kernel[2][2] ~^ image[15][9] + kernel[2][3] ~^ image[15][10] + kernel[2][4] ~^ image[15][11] + kernel[3][0] ~^ image[16][7] + kernel[3][1] ~^ image[16][8] + kernel[3][2] ~^ image[16][9] + kernel[3][3] ~^ image[16][10] + kernel[3][4] ~^ image[16][11] + kernel[4][0] ~^ image[17][7] + kernel[4][1] ~^ image[17][8] + kernel[4][2] ~^ image[17][9] + kernel[4][3] ~^ image[17][10] + kernel[4][4] ~^ image[17][11];
assign xor_sum[13][8] = kernel[0][0] ~^ image[13][8] + kernel[0][1] ~^ image[13][9] + kernel[0][2] ~^ image[13][10] + kernel[0][3] ~^ image[13][11] + kernel[0][4] ~^ image[13][12] + kernel[1][0] ~^ image[14][8] + kernel[1][1] ~^ image[14][9] + kernel[1][2] ~^ image[14][10] + kernel[1][3] ~^ image[14][11] + kernel[1][4] ~^ image[14][12] + kernel[2][0] ~^ image[15][8] + kernel[2][1] ~^ image[15][9] + kernel[2][2] ~^ image[15][10] + kernel[2][3] ~^ image[15][11] + kernel[2][4] ~^ image[15][12] + kernel[3][0] ~^ image[16][8] + kernel[3][1] ~^ image[16][9] + kernel[3][2] ~^ image[16][10] + kernel[3][3] ~^ image[16][11] + kernel[3][4] ~^ image[16][12] + kernel[4][0] ~^ image[17][8] + kernel[4][1] ~^ image[17][9] + kernel[4][2] ~^ image[17][10] + kernel[4][3] ~^ image[17][11] + kernel[4][4] ~^ image[17][12];
assign xor_sum[13][9] = kernel[0][0] ~^ image[13][9] + kernel[0][1] ~^ image[13][10] + kernel[0][2] ~^ image[13][11] + kernel[0][3] ~^ image[13][12] + kernel[0][4] ~^ image[13][13] + kernel[1][0] ~^ image[14][9] + kernel[1][1] ~^ image[14][10] + kernel[1][2] ~^ image[14][11] + kernel[1][3] ~^ image[14][12] + kernel[1][4] ~^ image[14][13] + kernel[2][0] ~^ image[15][9] + kernel[2][1] ~^ image[15][10] + kernel[2][2] ~^ image[15][11] + kernel[2][3] ~^ image[15][12] + kernel[2][4] ~^ image[15][13] + kernel[3][0] ~^ image[16][9] + kernel[3][1] ~^ image[16][10] + kernel[3][2] ~^ image[16][11] + kernel[3][3] ~^ image[16][12] + kernel[3][4] ~^ image[16][13] + kernel[4][0] ~^ image[17][9] + kernel[4][1] ~^ image[17][10] + kernel[4][2] ~^ image[17][11] + kernel[4][3] ~^ image[17][12] + kernel[4][4] ~^ image[17][13];
assign xor_sum[13][10] = kernel[0][0] ~^ image[13][10] + kernel[0][1] ~^ image[13][11] + kernel[0][2] ~^ image[13][12] + kernel[0][3] ~^ image[13][13] + kernel[0][4] ~^ image[13][14] + kernel[1][0] ~^ image[14][10] + kernel[1][1] ~^ image[14][11] + kernel[1][2] ~^ image[14][12] + kernel[1][3] ~^ image[14][13] + kernel[1][4] ~^ image[14][14] + kernel[2][0] ~^ image[15][10] + kernel[2][1] ~^ image[15][11] + kernel[2][2] ~^ image[15][12] + kernel[2][3] ~^ image[15][13] + kernel[2][4] ~^ image[15][14] + kernel[3][0] ~^ image[16][10] + kernel[3][1] ~^ image[16][11] + kernel[3][2] ~^ image[16][12] + kernel[3][3] ~^ image[16][13] + kernel[3][4] ~^ image[16][14] + kernel[4][0] ~^ image[17][10] + kernel[4][1] ~^ image[17][11] + kernel[4][2] ~^ image[17][12] + kernel[4][3] ~^ image[17][13] + kernel[4][4] ~^ image[17][14];
assign xor_sum[13][11] = kernel[0][0] ~^ image[13][11] + kernel[0][1] ~^ image[13][12] + kernel[0][2] ~^ image[13][13] + kernel[0][3] ~^ image[13][14] + kernel[0][4] ~^ image[13][15] + kernel[1][0] ~^ image[14][11] + kernel[1][1] ~^ image[14][12] + kernel[1][2] ~^ image[14][13] + kernel[1][3] ~^ image[14][14] + kernel[1][4] ~^ image[14][15] + kernel[2][0] ~^ image[15][11] + kernel[2][1] ~^ image[15][12] + kernel[2][2] ~^ image[15][13] + kernel[2][3] ~^ image[15][14] + kernel[2][4] ~^ image[15][15] + kernel[3][0] ~^ image[16][11] + kernel[3][1] ~^ image[16][12] + kernel[3][2] ~^ image[16][13] + kernel[3][3] ~^ image[16][14] + kernel[3][4] ~^ image[16][15] + kernel[4][0] ~^ image[17][11] + kernel[4][1] ~^ image[17][12] + kernel[4][2] ~^ image[17][13] + kernel[4][3] ~^ image[17][14] + kernel[4][4] ~^ image[17][15];
assign xor_sum[13][12] = kernel[0][0] ~^ image[13][12] + kernel[0][1] ~^ image[13][13] + kernel[0][2] ~^ image[13][14] + kernel[0][3] ~^ image[13][15] + kernel[0][4] ~^ image[13][16] + kernel[1][0] ~^ image[14][12] + kernel[1][1] ~^ image[14][13] + kernel[1][2] ~^ image[14][14] + kernel[1][3] ~^ image[14][15] + kernel[1][4] ~^ image[14][16] + kernel[2][0] ~^ image[15][12] + kernel[2][1] ~^ image[15][13] + kernel[2][2] ~^ image[15][14] + kernel[2][3] ~^ image[15][15] + kernel[2][4] ~^ image[15][16] + kernel[3][0] ~^ image[16][12] + kernel[3][1] ~^ image[16][13] + kernel[3][2] ~^ image[16][14] + kernel[3][3] ~^ image[16][15] + kernel[3][4] ~^ image[16][16] + kernel[4][0] ~^ image[17][12] + kernel[4][1] ~^ image[17][13] + kernel[4][2] ~^ image[17][14] + kernel[4][3] ~^ image[17][15] + kernel[4][4] ~^ image[17][16];
assign xor_sum[13][13] = kernel[0][0] ~^ image[13][13] + kernel[0][1] ~^ image[13][14] + kernel[0][2] ~^ image[13][15] + kernel[0][3] ~^ image[13][16] + kernel[0][4] ~^ image[13][17] + kernel[1][0] ~^ image[14][13] + kernel[1][1] ~^ image[14][14] + kernel[1][2] ~^ image[14][15] + kernel[1][3] ~^ image[14][16] + kernel[1][4] ~^ image[14][17] + kernel[2][0] ~^ image[15][13] + kernel[2][1] ~^ image[15][14] + kernel[2][2] ~^ image[15][15] + kernel[2][3] ~^ image[15][16] + kernel[2][4] ~^ image[15][17] + kernel[3][0] ~^ image[16][13] + kernel[3][1] ~^ image[16][14] + kernel[3][2] ~^ image[16][15] + kernel[3][3] ~^ image[16][16] + kernel[3][4] ~^ image[16][17] + kernel[4][0] ~^ image[17][13] + kernel[4][1] ~^ image[17][14] + kernel[4][2] ~^ image[17][15] + kernel[4][3] ~^ image[17][16] + kernel[4][4] ~^ image[17][17];
assign xor_sum[13][14] = kernel[0][0] ~^ image[13][14] + kernel[0][1] ~^ image[13][15] + kernel[0][2] ~^ image[13][16] + kernel[0][3] ~^ image[13][17] + kernel[0][4] ~^ image[13][18] + kernel[1][0] ~^ image[14][14] + kernel[1][1] ~^ image[14][15] + kernel[1][2] ~^ image[14][16] + kernel[1][3] ~^ image[14][17] + kernel[1][4] ~^ image[14][18] + kernel[2][0] ~^ image[15][14] + kernel[2][1] ~^ image[15][15] + kernel[2][2] ~^ image[15][16] + kernel[2][3] ~^ image[15][17] + kernel[2][4] ~^ image[15][18] + kernel[3][0] ~^ image[16][14] + kernel[3][1] ~^ image[16][15] + kernel[3][2] ~^ image[16][16] + kernel[3][3] ~^ image[16][17] + kernel[3][4] ~^ image[16][18] + kernel[4][0] ~^ image[17][14] + kernel[4][1] ~^ image[17][15] + kernel[4][2] ~^ image[17][16] + kernel[4][3] ~^ image[17][17] + kernel[4][4] ~^ image[17][18];
assign xor_sum[13][15] = kernel[0][0] ~^ image[13][15] + kernel[0][1] ~^ image[13][16] + kernel[0][2] ~^ image[13][17] + kernel[0][3] ~^ image[13][18] + kernel[0][4] ~^ image[13][19] + kernel[1][0] ~^ image[14][15] + kernel[1][1] ~^ image[14][16] + kernel[1][2] ~^ image[14][17] + kernel[1][3] ~^ image[14][18] + kernel[1][4] ~^ image[14][19] + kernel[2][0] ~^ image[15][15] + kernel[2][1] ~^ image[15][16] + kernel[2][2] ~^ image[15][17] + kernel[2][3] ~^ image[15][18] + kernel[2][4] ~^ image[15][19] + kernel[3][0] ~^ image[16][15] + kernel[3][1] ~^ image[16][16] + kernel[3][2] ~^ image[16][17] + kernel[3][3] ~^ image[16][18] + kernel[3][4] ~^ image[16][19] + kernel[4][0] ~^ image[17][15] + kernel[4][1] ~^ image[17][16] + kernel[4][2] ~^ image[17][17] + kernel[4][3] ~^ image[17][18] + kernel[4][4] ~^ image[17][19];
assign xor_sum[13][16] = kernel[0][0] ~^ image[13][16] + kernel[0][1] ~^ image[13][17] + kernel[0][2] ~^ image[13][18] + kernel[0][3] ~^ image[13][19] + kernel[0][4] ~^ image[13][20] + kernel[1][0] ~^ image[14][16] + kernel[1][1] ~^ image[14][17] + kernel[1][2] ~^ image[14][18] + kernel[1][3] ~^ image[14][19] + kernel[1][4] ~^ image[14][20] + kernel[2][0] ~^ image[15][16] + kernel[2][1] ~^ image[15][17] + kernel[2][2] ~^ image[15][18] + kernel[2][3] ~^ image[15][19] + kernel[2][4] ~^ image[15][20] + kernel[3][0] ~^ image[16][16] + kernel[3][1] ~^ image[16][17] + kernel[3][2] ~^ image[16][18] + kernel[3][3] ~^ image[16][19] + kernel[3][4] ~^ image[16][20] + kernel[4][0] ~^ image[17][16] + kernel[4][1] ~^ image[17][17] + kernel[4][2] ~^ image[17][18] + kernel[4][3] ~^ image[17][19] + kernel[4][4] ~^ image[17][20];
assign xor_sum[13][17] = kernel[0][0] ~^ image[13][17] + kernel[0][1] ~^ image[13][18] + kernel[0][2] ~^ image[13][19] + kernel[0][3] ~^ image[13][20] + kernel[0][4] ~^ image[13][21] + kernel[1][0] ~^ image[14][17] + kernel[1][1] ~^ image[14][18] + kernel[1][2] ~^ image[14][19] + kernel[1][3] ~^ image[14][20] + kernel[1][4] ~^ image[14][21] + kernel[2][0] ~^ image[15][17] + kernel[2][1] ~^ image[15][18] + kernel[2][2] ~^ image[15][19] + kernel[2][3] ~^ image[15][20] + kernel[2][4] ~^ image[15][21] + kernel[3][0] ~^ image[16][17] + kernel[3][1] ~^ image[16][18] + kernel[3][2] ~^ image[16][19] + kernel[3][3] ~^ image[16][20] + kernel[3][4] ~^ image[16][21] + kernel[4][0] ~^ image[17][17] + kernel[4][1] ~^ image[17][18] + kernel[4][2] ~^ image[17][19] + kernel[4][3] ~^ image[17][20] + kernel[4][4] ~^ image[17][21];
assign xor_sum[13][18] = kernel[0][0] ~^ image[13][18] + kernel[0][1] ~^ image[13][19] + kernel[0][2] ~^ image[13][20] + kernel[0][3] ~^ image[13][21] + kernel[0][4] ~^ image[13][22] + kernel[1][0] ~^ image[14][18] + kernel[1][1] ~^ image[14][19] + kernel[1][2] ~^ image[14][20] + kernel[1][3] ~^ image[14][21] + kernel[1][4] ~^ image[14][22] + kernel[2][0] ~^ image[15][18] + kernel[2][1] ~^ image[15][19] + kernel[2][2] ~^ image[15][20] + kernel[2][3] ~^ image[15][21] + kernel[2][4] ~^ image[15][22] + kernel[3][0] ~^ image[16][18] + kernel[3][1] ~^ image[16][19] + kernel[3][2] ~^ image[16][20] + kernel[3][3] ~^ image[16][21] + kernel[3][4] ~^ image[16][22] + kernel[4][0] ~^ image[17][18] + kernel[4][1] ~^ image[17][19] + kernel[4][2] ~^ image[17][20] + kernel[4][3] ~^ image[17][21] + kernel[4][4] ~^ image[17][22];
assign xor_sum[13][19] = kernel[0][0] ~^ image[13][19] + kernel[0][1] ~^ image[13][20] + kernel[0][2] ~^ image[13][21] + kernel[0][3] ~^ image[13][22] + kernel[0][4] ~^ image[13][23] + kernel[1][0] ~^ image[14][19] + kernel[1][1] ~^ image[14][20] + kernel[1][2] ~^ image[14][21] + kernel[1][3] ~^ image[14][22] + kernel[1][4] ~^ image[14][23] + kernel[2][0] ~^ image[15][19] + kernel[2][1] ~^ image[15][20] + kernel[2][2] ~^ image[15][21] + kernel[2][3] ~^ image[15][22] + kernel[2][4] ~^ image[15][23] + kernel[3][0] ~^ image[16][19] + kernel[3][1] ~^ image[16][20] + kernel[3][2] ~^ image[16][21] + kernel[3][3] ~^ image[16][22] + kernel[3][4] ~^ image[16][23] + kernel[4][0] ~^ image[17][19] + kernel[4][1] ~^ image[17][20] + kernel[4][2] ~^ image[17][21] + kernel[4][3] ~^ image[17][22] + kernel[4][4] ~^ image[17][23];
assign xor_sum[13][20] = kernel[0][0] ~^ image[13][20] + kernel[0][1] ~^ image[13][21] + kernel[0][2] ~^ image[13][22] + kernel[0][3] ~^ image[13][23] + kernel[0][4] ~^ image[13][24] + kernel[1][0] ~^ image[14][20] + kernel[1][1] ~^ image[14][21] + kernel[1][2] ~^ image[14][22] + kernel[1][3] ~^ image[14][23] + kernel[1][4] ~^ image[14][24] + kernel[2][0] ~^ image[15][20] + kernel[2][1] ~^ image[15][21] + kernel[2][2] ~^ image[15][22] + kernel[2][3] ~^ image[15][23] + kernel[2][4] ~^ image[15][24] + kernel[3][0] ~^ image[16][20] + kernel[3][1] ~^ image[16][21] + kernel[3][2] ~^ image[16][22] + kernel[3][3] ~^ image[16][23] + kernel[3][4] ~^ image[16][24] + kernel[4][0] ~^ image[17][20] + kernel[4][1] ~^ image[17][21] + kernel[4][2] ~^ image[17][22] + kernel[4][3] ~^ image[17][23] + kernel[4][4] ~^ image[17][24];
assign xor_sum[13][21] = kernel[0][0] ~^ image[13][21] + kernel[0][1] ~^ image[13][22] + kernel[0][2] ~^ image[13][23] + kernel[0][3] ~^ image[13][24] + kernel[0][4] ~^ image[13][25] + kernel[1][0] ~^ image[14][21] + kernel[1][1] ~^ image[14][22] + kernel[1][2] ~^ image[14][23] + kernel[1][3] ~^ image[14][24] + kernel[1][4] ~^ image[14][25] + kernel[2][0] ~^ image[15][21] + kernel[2][1] ~^ image[15][22] + kernel[2][2] ~^ image[15][23] + kernel[2][3] ~^ image[15][24] + kernel[2][4] ~^ image[15][25] + kernel[3][0] ~^ image[16][21] + kernel[3][1] ~^ image[16][22] + kernel[3][2] ~^ image[16][23] + kernel[3][3] ~^ image[16][24] + kernel[3][4] ~^ image[16][25] + kernel[4][0] ~^ image[17][21] + kernel[4][1] ~^ image[17][22] + kernel[4][2] ~^ image[17][23] + kernel[4][3] ~^ image[17][24] + kernel[4][4] ~^ image[17][25];
assign xor_sum[13][22] = kernel[0][0] ~^ image[13][22] + kernel[0][1] ~^ image[13][23] + kernel[0][2] ~^ image[13][24] + kernel[0][3] ~^ image[13][25] + kernel[0][4] ~^ image[13][26] + kernel[1][0] ~^ image[14][22] + kernel[1][1] ~^ image[14][23] + kernel[1][2] ~^ image[14][24] + kernel[1][3] ~^ image[14][25] + kernel[1][4] ~^ image[14][26] + kernel[2][0] ~^ image[15][22] + kernel[2][1] ~^ image[15][23] + kernel[2][2] ~^ image[15][24] + kernel[2][3] ~^ image[15][25] + kernel[2][4] ~^ image[15][26] + kernel[3][0] ~^ image[16][22] + kernel[3][1] ~^ image[16][23] + kernel[3][2] ~^ image[16][24] + kernel[3][3] ~^ image[16][25] + kernel[3][4] ~^ image[16][26] + kernel[4][0] ~^ image[17][22] + kernel[4][1] ~^ image[17][23] + kernel[4][2] ~^ image[17][24] + kernel[4][3] ~^ image[17][25] + kernel[4][4] ~^ image[17][26];
assign xor_sum[13][23] = kernel[0][0] ~^ image[13][23] + kernel[0][1] ~^ image[13][24] + kernel[0][2] ~^ image[13][25] + kernel[0][3] ~^ image[13][26] + kernel[0][4] ~^ image[13][27] + kernel[1][0] ~^ image[14][23] + kernel[1][1] ~^ image[14][24] + kernel[1][2] ~^ image[14][25] + kernel[1][3] ~^ image[14][26] + kernel[1][4] ~^ image[14][27] + kernel[2][0] ~^ image[15][23] + kernel[2][1] ~^ image[15][24] + kernel[2][2] ~^ image[15][25] + kernel[2][3] ~^ image[15][26] + kernel[2][4] ~^ image[15][27] + kernel[3][0] ~^ image[16][23] + kernel[3][1] ~^ image[16][24] + kernel[3][2] ~^ image[16][25] + kernel[3][3] ~^ image[16][26] + kernel[3][4] ~^ image[16][27] + kernel[4][0] ~^ image[17][23] + kernel[4][1] ~^ image[17][24] + kernel[4][2] ~^ image[17][25] + kernel[4][3] ~^ image[17][26] + kernel[4][4] ~^ image[17][27];
assign xor_sum[14][0] = kernel[0][0] ~^ image[14][0] + kernel[0][1] ~^ image[14][1] + kernel[0][2] ~^ image[14][2] + kernel[0][3] ~^ image[14][3] + kernel[0][4] ~^ image[14][4] + kernel[1][0] ~^ image[15][0] + kernel[1][1] ~^ image[15][1] + kernel[1][2] ~^ image[15][2] + kernel[1][3] ~^ image[15][3] + kernel[1][4] ~^ image[15][4] + kernel[2][0] ~^ image[16][0] + kernel[2][1] ~^ image[16][1] + kernel[2][2] ~^ image[16][2] + kernel[2][3] ~^ image[16][3] + kernel[2][4] ~^ image[16][4] + kernel[3][0] ~^ image[17][0] + kernel[3][1] ~^ image[17][1] + kernel[3][2] ~^ image[17][2] + kernel[3][3] ~^ image[17][3] + kernel[3][4] ~^ image[17][4] + kernel[4][0] ~^ image[18][0] + kernel[4][1] ~^ image[18][1] + kernel[4][2] ~^ image[18][2] + kernel[4][3] ~^ image[18][3] + kernel[4][4] ~^ image[18][4];
assign xor_sum[14][1] = kernel[0][0] ~^ image[14][1] + kernel[0][1] ~^ image[14][2] + kernel[0][2] ~^ image[14][3] + kernel[0][3] ~^ image[14][4] + kernel[0][4] ~^ image[14][5] + kernel[1][0] ~^ image[15][1] + kernel[1][1] ~^ image[15][2] + kernel[1][2] ~^ image[15][3] + kernel[1][3] ~^ image[15][4] + kernel[1][4] ~^ image[15][5] + kernel[2][0] ~^ image[16][1] + kernel[2][1] ~^ image[16][2] + kernel[2][2] ~^ image[16][3] + kernel[2][3] ~^ image[16][4] + kernel[2][4] ~^ image[16][5] + kernel[3][0] ~^ image[17][1] + kernel[3][1] ~^ image[17][2] + kernel[3][2] ~^ image[17][3] + kernel[3][3] ~^ image[17][4] + kernel[3][4] ~^ image[17][5] + kernel[4][0] ~^ image[18][1] + kernel[4][1] ~^ image[18][2] + kernel[4][2] ~^ image[18][3] + kernel[4][3] ~^ image[18][4] + kernel[4][4] ~^ image[18][5];
assign xor_sum[14][2] = kernel[0][0] ~^ image[14][2] + kernel[0][1] ~^ image[14][3] + kernel[0][2] ~^ image[14][4] + kernel[0][3] ~^ image[14][5] + kernel[0][4] ~^ image[14][6] + kernel[1][0] ~^ image[15][2] + kernel[1][1] ~^ image[15][3] + kernel[1][2] ~^ image[15][4] + kernel[1][3] ~^ image[15][5] + kernel[1][4] ~^ image[15][6] + kernel[2][0] ~^ image[16][2] + kernel[2][1] ~^ image[16][3] + kernel[2][2] ~^ image[16][4] + kernel[2][3] ~^ image[16][5] + kernel[2][4] ~^ image[16][6] + kernel[3][0] ~^ image[17][2] + kernel[3][1] ~^ image[17][3] + kernel[3][2] ~^ image[17][4] + kernel[3][3] ~^ image[17][5] + kernel[3][4] ~^ image[17][6] + kernel[4][0] ~^ image[18][2] + kernel[4][1] ~^ image[18][3] + kernel[4][2] ~^ image[18][4] + kernel[4][3] ~^ image[18][5] + kernel[4][4] ~^ image[18][6];
assign xor_sum[14][3] = kernel[0][0] ~^ image[14][3] + kernel[0][1] ~^ image[14][4] + kernel[0][2] ~^ image[14][5] + kernel[0][3] ~^ image[14][6] + kernel[0][4] ~^ image[14][7] + kernel[1][0] ~^ image[15][3] + kernel[1][1] ~^ image[15][4] + kernel[1][2] ~^ image[15][5] + kernel[1][3] ~^ image[15][6] + kernel[1][4] ~^ image[15][7] + kernel[2][0] ~^ image[16][3] + kernel[2][1] ~^ image[16][4] + kernel[2][2] ~^ image[16][5] + kernel[2][3] ~^ image[16][6] + kernel[2][4] ~^ image[16][7] + kernel[3][0] ~^ image[17][3] + kernel[3][1] ~^ image[17][4] + kernel[3][2] ~^ image[17][5] + kernel[3][3] ~^ image[17][6] + kernel[3][4] ~^ image[17][7] + kernel[4][0] ~^ image[18][3] + kernel[4][1] ~^ image[18][4] + kernel[4][2] ~^ image[18][5] + kernel[4][3] ~^ image[18][6] + kernel[4][4] ~^ image[18][7];
assign xor_sum[14][4] = kernel[0][0] ~^ image[14][4] + kernel[0][1] ~^ image[14][5] + kernel[0][2] ~^ image[14][6] + kernel[0][3] ~^ image[14][7] + kernel[0][4] ~^ image[14][8] + kernel[1][0] ~^ image[15][4] + kernel[1][1] ~^ image[15][5] + kernel[1][2] ~^ image[15][6] + kernel[1][3] ~^ image[15][7] + kernel[1][4] ~^ image[15][8] + kernel[2][0] ~^ image[16][4] + kernel[2][1] ~^ image[16][5] + kernel[2][2] ~^ image[16][6] + kernel[2][3] ~^ image[16][7] + kernel[2][4] ~^ image[16][8] + kernel[3][0] ~^ image[17][4] + kernel[3][1] ~^ image[17][5] + kernel[3][2] ~^ image[17][6] + kernel[3][3] ~^ image[17][7] + kernel[3][4] ~^ image[17][8] + kernel[4][0] ~^ image[18][4] + kernel[4][1] ~^ image[18][5] + kernel[4][2] ~^ image[18][6] + kernel[4][3] ~^ image[18][7] + kernel[4][4] ~^ image[18][8];
assign xor_sum[14][5] = kernel[0][0] ~^ image[14][5] + kernel[0][1] ~^ image[14][6] + kernel[0][2] ~^ image[14][7] + kernel[0][3] ~^ image[14][8] + kernel[0][4] ~^ image[14][9] + kernel[1][0] ~^ image[15][5] + kernel[1][1] ~^ image[15][6] + kernel[1][2] ~^ image[15][7] + kernel[1][3] ~^ image[15][8] + kernel[1][4] ~^ image[15][9] + kernel[2][0] ~^ image[16][5] + kernel[2][1] ~^ image[16][6] + kernel[2][2] ~^ image[16][7] + kernel[2][3] ~^ image[16][8] + kernel[2][4] ~^ image[16][9] + kernel[3][0] ~^ image[17][5] + kernel[3][1] ~^ image[17][6] + kernel[3][2] ~^ image[17][7] + kernel[3][3] ~^ image[17][8] + kernel[3][4] ~^ image[17][9] + kernel[4][0] ~^ image[18][5] + kernel[4][1] ~^ image[18][6] + kernel[4][2] ~^ image[18][7] + kernel[4][3] ~^ image[18][8] + kernel[4][4] ~^ image[18][9];
assign xor_sum[14][6] = kernel[0][0] ~^ image[14][6] + kernel[0][1] ~^ image[14][7] + kernel[0][2] ~^ image[14][8] + kernel[0][3] ~^ image[14][9] + kernel[0][4] ~^ image[14][10] + kernel[1][0] ~^ image[15][6] + kernel[1][1] ~^ image[15][7] + kernel[1][2] ~^ image[15][8] + kernel[1][3] ~^ image[15][9] + kernel[1][4] ~^ image[15][10] + kernel[2][0] ~^ image[16][6] + kernel[2][1] ~^ image[16][7] + kernel[2][2] ~^ image[16][8] + kernel[2][3] ~^ image[16][9] + kernel[2][4] ~^ image[16][10] + kernel[3][0] ~^ image[17][6] + kernel[3][1] ~^ image[17][7] + kernel[3][2] ~^ image[17][8] + kernel[3][3] ~^ image[17][9] + kernel[3][4] ~^ image[17][10] + kernel[4][0] ~^ image[18][6] + kernel[4][1] ~^ image[18][7] + kernel[4][2] ~^ image[18][8] + kernel[4][3] ~^ image[18][9] + kernel[4][4] ~^ image[18][10];
assign xor_sum[14][7] = kernel[0][0] ~^ image[14][7] + kernel[0][1] ~^ image[14][8] + kernel[0][2] ~^ image[14][9] + kernel[0][3] ~^ image[14][10] + kernel[0][4] ~^ image[14][11] + kernel[1][0] ~^ image[15][7] + kernel[1][1] ~^ image[15][8] + kernel[1][2] ~^ image[15][9] + kernel[1][3] ~^ image[15][10] + kernel[1][4] ~^ image[15][11] + kernel[2][0] ~^ image[16][7] + kernel[2][1] ~^ image[16][8] + kernel[2][2] ~^ image[16][9] + kernel[2][3] ~^ image[16][10] + kernel[2][4] ~^ image[16][11] + kernel[3][0] ~^ image[17][7] + kernel[3][1] ~^ image[17][8] + kernel[3][2] ~^ image[17][9] + kernel[3][3] ~^ image[17][10] + kernel[3][4] ~^ image[17][11] + kernel[4][0] ~^ image[18][7] + kernel[4][1] ~^ image[18][8] + kernel[4][2] ~^ image[18][9] + kernel[4][3] ~^ image[18][10] + kernel[4][4] ~^ image[18][11];
assign xor_sum[14][8] = kernel[0][0] ~^ image[14][8] + kernel[0][1] ~^ image[14][9] + kernel[0][2] ~^ image[14][10] + kernel[0][3] ~^ image[14][11] + kernel[0][4] ~^ image[14][12] + kernel[1][0] ~^ image[15][8] + kernel[1][1] ~^ image[15][9] + kernel[1][2] ~^ image[15][10] + kernel[1][3] ~^ image[15][11] + kernel[1][4] ~^ image[15][12] + kernel[2][0] ~^ image[16][8] + kernel[2][1] ~^ image[16][9] + kernel[2][2] ~^ image[16][10] + kernel[2][3] ~^ image[16][11] + kernel[2][4] ~^ image[16][12] + kernel[3][0] ~^ image[17][8] + kernel[3][1] ~^ image[17][9] + kernel[3][2] ~^ image[17][10] + kernel[3][3] ~^ image[17][11] + kernel[3][4] ~^ image[17][12] + kernel[4][0] ~^ image[18][8] + kernel[4][1] ~^ image[18][9] + kernel[4][2] ~^ image[18][10] + kernel[4][3] ~^ image[18][11] + kernel[4][4] ~^ image[18][12];
assign xor_sum[14][9] = kernel[0][0] ~^ image[14][9] + kernel[0][1] ~^ image[14][10] + kernel[0][2] ~^ image[14][11] + kernel[0][3] ~^ image[14][12] + kernel[0][4] ~^ image[14][13] + kernel[1][0] ~^ image[15][9] + kernel[1][1] ~^ image[15][10] + kernel[1][2] ~^ image[15][11] + kernel[1][3] ~^ image[15][12] + kernel[1][4] ~^ image[15][13] + kernel[2][0] ~^ image[16][9] + kernel[2][1] ~^ image[16][10] + kernel[2][2] ~^ image[16][11] + kernel[2][3] ~^ image[16][12] + kernel[2][4] ~^ image[16][13] + kernel[3][0] ~^ image[17][9] + kernel[3][1] ~^ image[17][10] + kernel[3][2] ~^ image[17][11] + kernel[3][3] ~^ image[17][12] + kernel[3][4] ~^ image[17][13] + kernel[4][0] ~^ image[18][9] + kernel[4][1] ~^ image[18][10] + kernel[4][2] ~^ image[18][11] + kernel[4][3] ~^ image[18][12] + kernel[4][4] ~^ image[18][13];
assign xor_sum[14][10] = kernel[0][0] ~^ image[14][10] + kernel[0][1] ~^ image[14][11] + kernel[0][2] ~^ image[14][12] + kernel[0][3] ~^ image[14][13] + kernel[0][4] ~^ image[14][14] + kernel[1][0] ~^ image[15][10] + kernel[1][1] ~^ image[15][11] + kernel[1][2] ~^ image[15][12] + kernel[1][3] ~^ image[15][13] + kernel[1][4] ~^ image[15][14] + kernel[2][0] ~^ image[16][10] + kernel[2][1] ~^ image[16][11] + kernel[2][2] ~^ image[16][12] + kernel[2][3] ~^ image[16][13] + kernel[2][4] ~^ image[16][14] + kernel[3][0] ~^ image[17][10] + kernel[3][1] ~^ image[17][11] + kernel[3][2] ~^ image[17][12] + kernel[3][3] ~^ image[17][13] + kernel[3][4] ~^ image[17][14] + kernel[4][0] ~^ image[18][10] + kernel[4][1] ~^ image[18][11] + kernel[4][2] ~^ image[18][12] + kernel[4][3] ~^ image[18][13] + kernel[4][4] ~^ image[18][14];
assign xor_sum[14][11] = kernel[0][0] ~^ image[14][11] + kernel[0][1] ~^ image[14][12] + kernel[0][2] ~^ image[14][13] + kernel[0][3] ~^ image[14][14] + kernel[0][4] ~^ image[14][15] + kernel[1][0] ~^ image[15][11] + kernel[1][1] ~^ image[15][12] + kernel[1][2] ~^ image[15][13] + kernel[1][3] ~^ image[15][14] + kernel[1][4] ~^ image[15][15] + kernel[2][0] ~^ image[16][11] + kernel[2][1] ~^ image[16][12] + kernel[2][2] ~^ image[16][13] + kernel[2][3] ~^ image[16][14] + kernel[2][4] ~^ image[16][15] + kernel[3][0] ~^ image[17][11] + kernel[3][1] ~^ image[17][12] + kernel[3][2] ~^ image[17][13] + kernel[3][3] ~^ image[17][14] + kernel[3][4] ~^ image[17][15] + kernel[4][0] ~^ image[18][11] + kernel[4][1] ~^ image[18][12] + kernel[4][2] ~^ image[18][13] + kernel[4][3] ~^ image[18][14] + kernel[4][4] ~^ image[18][15];
assign xor_sum[14][12] = kernel[0][0] ~^ image[14][12] + kernel[0][1] ~^ image[14][13] + kernel[0][2] ~^ image[14][14] + kernel[0][3] ~^ image[14][15] + kernel[0][4] ~^ image[14][16] + kernel[1][0] ~^ image[15][12] + kernel[1][1] ~^ image[15][13] + kernel[1][2] ~^ image[15][14] + kernel[1][3] ~^ image[15][15] + kernel[1][4] ~^ image[15][16] + kernel[2][0] ~^ image[16][12] + kernel[2][1] ~^ image[16][13] + kernel[2][2] ~^ image[16][14] + kernel[2][3] ~^ image[16][15] + kernel[2][4] ~^ image[16][16] + kernel[3][0] ~^ image[17][12] + kernel[3][1] ~^ image[17][13] + kernel[3][2] ~^ image[17][14] + kernel[3][3] ~^ image[17][15] + kernel[3][4] ~^ image[17][16] + kernel[4][0] ~^ image[18][12] + kernel[4][1] ~^ image[18][13] + kernel[4][2] ~^ image[18][14] + kernel[4][3] ~^ image[18][15] + kernel[4][4] ~^ image[18][16];
assign xor_sum[14][13] = kernel[0][0] ~^ image[14][13] + kernel[0][1] ~^ image[14][14] + kernel[0][2] ~^ image[14][15] + kernel[0][3] ~^ image[14][16] + kernel[0][4] ~^ image[14][17] + kernel[1][0] ~^ image[15][13] + kernel[1][1] ~^ image[15][14] + kernel[1][2] ~^ image[15][15] + kernel[1][3] ~^ image[15][16] + kernel[1][4] ~^ image[15][17] + kernel[2][0] ~^ image[16][13] + kernel[2][1] ~^ image[16][14] + kernel[2][2] ~^ image[16][15] + kernel[2][3] ~^ image[16][16] + kernel[2][4] ~^ image[16][17] + kernel[3][0] ~^ image[17][13] + kernel[3][1] ~^ image[17][14] + kernel[3][2] ~^ image[17][15] + kernel[3][3] ~^ image[17][16] + kernel[3][4] ~^ image[17][17] + kernel[4][0] ~^ image[18][13] + kernel[4][1] ~^ image[18][14] + kernel[4][2] ~^ image[18][15] + kernel[4][3] ~^ image[18][16] + kernel[4][4] ~^ image[18][17];
assign xor_sum[14][14] = kernel[0][0] ~^ image[14][14] + kernel[0][1] ~^ image[14][15] + kernel[0][2] ~^ image[14][16] + kernel[0][3] ~^ image[14][17] + kernel[0][4] ~^ image[14][18] + kernel[1][0] ~^ image[15][14] + kernel[1][1] ~^ image[15][15] + kernel[1][2] ~^ image[15][16] + kernel[1][3] ~^ image[15][17] + kernel[1][4] ~^ image[15][18] + kernel[2][0] ~^ image[16][14] + kernel[2][1] ~^ image[16][15] + kernel[2][2] ~^ image[16][16] + kernel[2][3] ~^ image[16][17] + kernel[2][4] ~^ image[16][18] + kernel[3][0] ~^ image[17][14] + kernel[3][1] ~^ image[17][15] + kernel[3][2] ~^ image[17][16] + kernel[3][3] ~^ image[17][17] + kernel[3][4] ~^ image[17][18] + kernel[4][0] ~^ image[18][14] + kernel[4][1] ~^ image[18][15] + kernel[4][2] ~^ image[18][16] + kernel[4][3] ~^ image[18][17] + kernel[4][4] ~^ image[18][18];
assign xor_sum[14][15] = kernel[0][0] ~^ image[14][15] + kernel[0][1] ~^ image[14][16] + kernel[0][2] ~^ image[14][17] + kernel[0][3] ~^ image[14][18] + kernel[0][4] ~^ image[14][19] + kernel[1][0] ~^ image[15][15] + kernel[1][1] ~^ image[15][16] + kernel[1][2] ~^ image[15][17] + kernel[1][3] ~^ image[15][18] + kernel[1][4] ~^ image[15][19] + kernel[2][0] ~^ image[16][15] + kernel[2][1] ~^ image[16][16] + kernel[2][2] ~^ image[16][17] + kernel[2][3] ~^ image[16][18] + kernel[2][4] ~^ image[16][19] + kernel[3][0] ~^ image[17][15] + kernel[3][1] ~^ image[17][16] + kernel[3][2] ~^ image[17][17] + kernel[3][3] ~^ image[17][18] + kernel[3][4] ~^ image[17][19] + kernel[4][0] ~^ image[18][15] + kernel[4][1] ~^ image[18][16] + kernel[4][2] ~^ image[18][17] + kernel[4][3] ~^ image[18][18] + kernel[4][4] ~^ image[18][19];
assign xor_sum[14][16] = kernel[0][0] ~^ image[14][16] + kernel[0][1] ~^ image[14][17] + kernel[0][2] ~^ image[14][18] + kernel[0][3] ~^ image[14][19] + kernel[0][4] ~^ image[14][20] + kernel[1][0] ~^ image[15][16] + kernel[1][1] ~^ image[15][17] + kernel[1][2] ~^ image[15][18] + kernel[1][3] ~^ image[15][19] + kernel[1][4] ~^ image[15][20] + kernel[2][0] ~^ image[16][16] + kernel[2][1] ~^ image[16][17] + kernel[2][2] ~^ image[16][18] + kernel[2][3] ~^ image[16][19] + kernel[2][4] ~^ image[16][20] + kernel[3][0] ~^ image[17][16] + kernel[3][1] ~^ image[17][17] + kernel[3][2] ~^ image[17][18] + kernel[3][3] ~^ image[17][19] + kernel[3][4] ~^ image[17][20] + kernel[4][0] ~^ image[18][16] + kernel[4][1] ~^ image[18][17] + kernel[4][2] ~^ image[18][18] + kernel[4][3] ~^ image[18][19] + kernel[4][4] ~^ image[18][20];
assign xor_sum[14][17] = kernel[0][0] ~^ image[14][17] + kernel[0][1] ~^ image[14][18] + kernel[0][2] ~^ image[14][19] + kernel[0][3] ~^ image[14][20] + kernel[0][4] ~^ image[14][21] + kernel[1][0] ~^ image[15][17] + kernel[1][1] ~^ image[15][18] + kernel[1][2] ~^ image[15][19] + kernel[1][3] ~^ image[15][20] + kernel[1][4] ~^ image[15][21] + kernel[2][0] ~^ image[16][17] + kernel[2][1] ~^ image[16][18] + kernel[2][2] ~^ image[16][19] + kernel[2][3] ~^ image[16][20] + kernel[2][4] ~^ image[16][21] + kernel[3][0] ~^ image[17][17] + kernel[3][1] ~^ image[17][18] + kernel[3][2] ~^ image[17][19] + kernel[3][3] ~^ image[17][20] + kernel[3][4] ~^ image[17][21] + kernel[4][0] ~^ image[18][17] + kernel[4][1] ~^ image[18][18] + kernel[4][2] ~^ image[18][19] + kernel[4][3] ~^ image[18][20] + kernel[4][4] ~^ image[18][21];
assign xor_sum[14][18] = kernel[0][0] ~^ image[14][18] + kernel[0][1] ~^ image[14][19] + kernel[0][2] ~^ image[14][20] + kernel[0][3] ~^ image[14][21] + kernel[0][4] ~^ image[14][22] + kernel[1][0] ~^ image[15][18] + kernel[1][1] ~^ image[15][19] + kernel[1][2] ~^ image[15][20] + kernel[1][3] ~^ image[15][21] + kernel[1][4] ~^ image[15][22] + kernel[2][0] ~^ image[16][18] + kernel[2][1] ~^ image[16][19] + kernel[2][2] ~^ image[16][20] + kernel[2][3] ~^ image[16][21] + kernel[2][4] ~^ image[16][22] + kernel[3][0] ~^ image[17][18] + kernel[3][1] ~^ image[17][19] + kernel[3][2] ~^ image[17][20] + kernel[3][3] ~^ image[17][21] + kernel[3][4] ~^ image[17][22] + kernel[4][0] ~^ image[18][18] + kernel[4][1] ~^ image[18][19] + kernel[4][2] ~^ image[18][20] + kernel[4][3] ~^ image[18][21] + kernel[4][4] ~^ image[18][22];
assign xor_sum[14][19] = kernel[0][0] ~^ image[14][19] + kernel[0][1] ~^ image[14][20] + kernel[0][2] ~^ image[14][21] + kernel[0][3] ~^ image[14][22] + kernel[0][4] ~^ image[14][23] + kernel[1][0] ~^ image[15][19] + kernel[1][1] ~^ image[15][20] + kernel[1][2] ~^ image[15][21] + kernel[1][3] ~^ image[15][22] + kernel[1][4] ~^ image[15][23] + kernel[2][0] ~^ image[16][19] + kernel[2][1] ~^ image[16][20] + kernel[2][2] ~^ image[16][21] + kernel[2][3] ~^ image[16][22] + kernel[2][4] ~^ image[16][23] + kernel[3][0] ~^ image[17][19] + kernel[3][1] ~^ image[17][20] + kernel[3][2] ~^ image[17][21] + kernel[3][3] ~^ image[17][22] + kernel[3][4] ~^ image[17][23] + kernel[4][0] ~^ image[18][19] + kernel[4][1] ~^ image[18][20] + kernel[4][2] ~^ image[18][21] + kernel[4][3] ~^ image[18][22] + kernel[4][4] ~^ image[18][23];
assign xor_sum[14][20] = kernel[0][0] ~^ image[14][20] + kernel[0][1] ~^ image[14][21] + kernel[0][2] ~^ image[14][22] + kernel[0][3] ~^ image[14][23] + kernel[0][4] ~^ image[14][24] + kernel[1][0] ~^ image[15][20] + kernel[1][1] ~^ image[15][21] + kernel[1][2] ~^ image[15][22] + kernel[1][3] ~^ image[15][23] + kernel[1][4] ~^ image[15][24] + kernel[2][0] ~^ image[16][20] + kernel[2][1] ~^ image[16][21] + kernel[2][2] ~^ image[16][22] + kernel[2][3] ~^ image[16][23] + kernel[2][4] ~^ image[16][24] + kernel[3][0] ~^ image[17][20] + kernel[3][1] ~^ image[17][21] + kernel[3][2] ~^ image[17][22] + kernel[3][3] ~^ image[17][23] + kernel[3][4] ~^ image[17][24] + kernel[4][0] ~^ image[18][20] + kernel[4][1] ~^ image[18][21] + kernel[4][2] ~^ image[18][22] + kernel[4][3] ~^ image[18][23] + kernel[4][4] ~^ image[18][24];
assign xor_sum[14][21] = kernel[0][0] ~^ image[14][21] + kernel[0][1] ~^ image[14][22] + kernel[0][2] ~^ image[14][23] + kernel[0][3] ~^ image[14][24] + kernel[0][4] ~^ image[14][25] + kernel[1][0] ~^ image[15][21] + kernel[1][1] ~^ image[15][22] + kernel[1][2] ~^ image[15][23] + kernel[1][3] ~^ image[15][24] + kernel[1][4] ~^ image[15][25] + kernel[2][0] ~^ image[16][21] + kernel[2][1] ~^ image[16][22] + kernel[2][2] ~^ image[16][23] + kernel[2][3] ~^ image[16][24] + kernel[2][4] ~^ image[16][25] + kernel[3][0] ~^ image[17][21] + kernel[3][1] ~^ image[17][22] + kernel[3][2] ~^ image[17][23] + kernel[3][3] ~^ image[17][24] + kernel[3][4] ~^ image[17][25] + kernel[4][0] ~^ image[18][21] + kernel[4][1] ~^ image[18][22] + kernel[4][2] ~^ image[18][23] + kernel[4][3] ~^ image[18][24] + kernel[4][4] ~^ image[18][25];
assign xor_sum[14][22] = kernel[0][0] ~^ image[14][22] + kernel[0][1] ~^ image[14][23] + kernel[0][2] ~^ image[14][24] + kernel[0][3] ~^ image[14][25] + kernel[0][4] ~^ image[14][26] + kernel[1][0] ~^ image[15][22] + kernel[1][1] ~^ image[15][23] + kernel[1][2] ~^ image[15][24] + kernel[1][3] ~^ image[15][25] + kernel[1][4] ~^ image[15][26] + kernel[2][0] ~^ image[16][22] + kernel[2][1] ~^ image[16][23] + kernel[2][2] ~^ image[16][24] + kernel[2][3] ~^ image[16][25] + kernel[2][4] ~^ image[16][26] + kernel[3][0] ~^ image[17][22] + kernel[3][1] ~^ image[17][23] + kernel[3][2] ~^ image[17][24] + kernel[3][3] ~^ image[17][25] + kernel[3][4] ~^ image[17][26] + kernel[4][0] ~^ image[18][22] + kernel[4][1] ~^ image[18][23] + kernel[4][2] ~^ image[18][24] + kernel[4][3] ~^ image[18][25] + kernel[4][4] ~^ image[18][26];
assign xor_sum[14][23] = kernel[0][0] ~^ image[14][23] + kernel[0][1] ~^ image[14][24] + kernel[0][2] ~^ image[14][25] + kernel[0][3] ~^ image[14][26] + kernel[0][4] ~^ image[14][27] + kernel[1][0] ~^ image[15][23] + kernel[1][1] ~^ image[15][24] + kernel[1][2] ~^ image[15][25] + kernel[1][3] ~^ image[15][26] + kernel[1][4] ~^ image[15][27] + kernel[2][0] ~^ image[16][23] + kernel[2][1] ~^ image[16][24] + kernel[2][2] ~^ image[16][25] + kernel[2][3] ~^ image[16][26] + kernel[2][4] ~^ image[16][27] + kernel[3][0] ~^ image[17][23] + kernel[3][1] ~^ image[17][24] + kernel[3][2] ~^ image[17][25] + kernel[3][3] ~^ image[17][26] + kernel[3][4] ~^ image[17][27] + kernel[4][0] ~^ image[18][23] + kernel[4][1] ~^ image[18][24] + kernel[4][2] ~^ image[18][25] + kernel[4][3] ~^ image[18][26] + kernel[4][4] ~^ image[18][27];
assign xor_sum[15][0] = kernel[0][0] ~^ image[15][0] + kernel[0][1] ~^ image[15][1] + kernel[0][2] ~^ image[15][2] + kernel[0][3] ~^ image[15][3] + kernel[0][4] ~^ image[15][4] + kernel[1][0] ~^ image[16][0] + kernel[1][1] ~^ image[16][1] + kernel[1][2] ~^ image[16][2] + kernel[1][3] ~^ image[16][3] + kernel[1][4] ~^ image[16][4] + kernel[2][0] ~^ image[17][0] + kernel[2][1] ~^ image[17][1] + kernel[2][2] ~^ image[17][2] + kernel[2][3] ~^ image[17][3] + kernel[2][4] ~^ image[17][4] + kernel[3][0] ~^ image[18][0] + kernel[3][1] ~^ image[18][1] + kernel[3][2] ~^ image[18][2] + kernel[3][3] ~^ image[18][3] + kernel[3][4] ~^ image[18][4] + kernel[4][0] ~^ image[19][0] + kernel[4][1] ~^ image[19][1] + kernel[4][2] ~^ image[19][2] + kernel[4][3] ~^ image[19][3] + kernel[4][4] ~^ image[19][4];
assign xor_sum[15][1] = kernel[0][0] ~^ image[15][1] + kernel[0][1] ~^ image[15][2] + kernel[0][2] ~^ image[15][3] + kernel[0][3] ~^ image[15][4] + kernel[0][4] ~^ image[15][5] + kernel[1][0] ~^ image[16][1] + kernel[1][1] ~^ image[16][2] + kernel[1][2] ~^ image[16][3] + kernel[1][3] ~^ image[16][4] + kernel[1][4] ~^ image[16][5] + kernel[2][0] ~^ image[17][1] + kernel[2][1] ~^ image[17][2] + kernel[2][2] ~^ image[17][3] + kernel[2][3] ~^ image[17][4] + kernel[2][4] ~^ image[17][5] + kernel[3][0] ~^ image[18][1] + kernel[3][1] ~^ image[18][2] + kernel[3][2] ~^ image[18][3] + kernel[3][3] ~^ image[18][4] + kernel[3][4] ~^ image[18][5] + kernel[4][0] ~^ image[19][1] + kernel[4][1] ~^ image[19][2] + kernel[4][2] ~^ image[19][3] + kernel[4][3] ~^ image[19][4] + kernel[4][4] ~^ image[19][5];
assign xor_sum[15][2] = kernel[0][0] ~^ image[15][2] + kernel[0][1] ~^ image[15][3] + kernel[0][2] ~^ image[15][4] + kernel[0][3] ~^ image[15][5] + kernel[0][4] ~^ image[15][6] + kernel[1][0] ~^ image[16][2] + kernel[1][1] ~^ image[16][3] + kernel[1][2] ~^ image[16][4] + kernel[1][3] ~^ image[16][5] + kernel[1][4] ~^ image[16][6] + kernel[2][0] ~^ image[17][2] + kernel[2][1] ~^ image[17][3] + kernel[2][2] ~^ image[17][4] + kernel[2][3] ~^ image[17][5] + kernel[2][4] ~^ image[17][6] + kernel[3][0] ~^ image[18][2] + kernel[3][1] ~^ image[18][3] + kernel[3][2] ~^ image[18][4] + kernel[3][3] ~^ image[18][5] + kernel[3][4] ~^ image[18][6] + kernel[4][0] ~^ image[19][2] + kernel[4][1] ~^ image[19][3] + kernel[4][2] ~^ image[19][4] + kernel[4][3] ~^ image[19][5] + kernel[4][4] ~^ image[19][6];
assign xor_sum[15][3] = kernel[0][0] ~^ image[15][3] + kernel[0][1] ~^ image[15][4] + kernel[0][2] ~^ image[15][5] + kernel[0][3] ~^ image[15][6] + kernel[0][4] ~^ image[15][7] + kernel[1][0] ~^ image[16][3] + kernel[1][1] ~^ image[16][4] + kernel[1][2] ~^ image[16][5] + kernel[1][3] ~^ image[16][6] + kernel[1][4] ~^ image[16][7] + kernel[2][0] ~^ image[17][3] + kernel[2][1] ~^ image[17][4] + kernel[2][2] ~^ image[17][5] + kernel[2][3] ~^ image[17][6] + kernel[2][4] ~^ image[17][7] + kernel[3][0] ~^ image[18][3] + kernel[3][1] ~^ image[18][4] + kernel[3][2] ~^ image[18][5] + kernel[3][3] ~^ image[18][6] + kernel[3][4] ~^ image[18][7] + kernel[4][0] ~^ image[19][3] + kernel[4][1] ~^ image[19][4] + kernel[4][2] ~^ image[19][5] + kernel[4][3] ~^ image[19][6] + kernel[4][4] ~^ image[19][7];
assign xor_sum[15][4] = kernel[0][0] ~^ image[15][4] + kernel[0][1] ~^ image[15][5] + kernel[0][2] ~^ image[15][6] + kernel[0][3] ~^ image[15][7] + kernel[0][4] ~^ image[15][8] + kernel[1][0] ~^ image[16][4] + kernel[1][1] ~^ image[16][5] + kernel[1][2] ~^ image[16][6] + kernel[1][3] ~^ image[16][7] + kernel[1][4] ~^ image[16][8] + kernel[2][0] ~^ image[17][4] + kernel[2][1] ~^ image[17][5] + kernel[2][2] ~^ image[17][6] + kernel[2][3] ~^ image[17][7] + kernel[2][4] ~^ image[17][8] + kernel[3][0] ~^ image[18][4] + kernel[3][1] ~^ image[18][5] + kernel[3][2] ~^ image[18][6] + kernel[3][3] ~^ image[18][7] + kernel[3][4] ~^ image[18][8] + kernel[4][0] ~^ image[19][4] + kernel[4][1] ~^ image[19][5] + kernel[4][2] ~^ image[19][6] + kernel[4][3] ~^ image[19][7] + kernel[4][4] ~^ image[19][8];
assign xor_sum[15][5] = kernel[0][0] ~^ image[15][5] + kernel[0][1] ~^ image[15][6] + kernel[0][2] ~^ image[15][7] + kernel[0][3] ~^ image[15][8] + kernel[0][4] ~^ image[15][9] + kernel[1][0] ~^ image[16][5] + kernel[1][1] ~^ image[16][6] + kernel[1][2] ~^ image[16][7] + kernel[1][3] ~^ image[16][8] + kernel[1][4] ~^ image[16][9] + kernel[2][0] ~^ image[17][5] + kernel[2][1] ~^ image[17][6] + kernel[2][2] ~^ image[17][7] + kernel[2][3] ~^ image[17][8] + kernel[2][4] ~^ image[17][9] + kernel[3][0] ~^ image[18][5] + kernel[3][1] ~^ image[18][6] + kernel[3][2] ~^ image[18][7] + kernel[3][3] ~^ image[18][8] + kernel[3][4] ~^ image[18][9] + kernel[4][0] ~^ image[19][5] + kernel[4][1] ~^ image[19][6] + kernel[4][2] ~^ image[19][7] + kernel[4][3] ~^ image[19][8] + kernel[4][4] ~^ image[19][9];
assign xor_sum[15][6] = kernel[0][0] ~^ image[15][6] + kernel[0][1] ~^ image[15][7] + kernel[0][2] ~^ image[15][8] + kernel[0][3] ~^ image[15][9] + kernel[0][4] ~^ image[15][10] + kernel[1][0] ~^ image[16][6] + kernel[1][1] ~^ image[16][7] + kernel[1][2] ~^ image[16][8] + kernel[1][3] ~^ image[16][9] + kernel[1][4] ~^ image[16][10] + kernel[2][0] ~^ image[17][6] + kernel[2][1] ~^ image[17][7] + kernel[2][2] ~^ image[17][8] + kernel[2][3] ~^ image[17][9] + kernel[2][4] ~^ image[17][10] + kernel[3][0] ~^ image[18][6] + kernel[3][1] ~^ image[18][7] + kernel[3][2] ~^ image[18][8] + kernel[3][3] ~^ image[18][9] + kernel[3][4] ~^ image[18][10] + kernel[4][0] ~^ image[19][6] + kernel[4][1] ~^ image[19][7] + kernel[4][2] ~^ image[19][8] + kernel[4][3] ~^ image[19][9] + kernel[4][4] ~^ image[19][10];
assign xor_sum[15][7] = kernel[0][0] ~^ image[15][7] + kernel[0][1] ~^ image[15][8] + kernel[0][2] ~^ image[15][9] + kernel[0][3] ~^ image[15][10] + kernel[0][4] ~^ image[15][11] + kernel[1][0] ~^ image[16][7] + kernel[1][1] ~^ image[16][8] + kernel[1][2] ~^ image[16][9] + kernel[1][3] ~^ image[16][10] + kernel[1][4] ~^ image[16][11] + kernel[2][0] ~^ image[17][7] + kernel[2][1] ~^ image[17][8] + kernel[2][2] ~^ image[17][9] + kernel[2][3] ~^ image[17][10] + kernel[2][4] ~^ image[17][11] + kernel[3][0] ~^ image[18][7] + kernel[3][1] ~^ image[18][8] + kernel[3][2] ~^ image[18][9] + kernel[3][3] ~^ image[18][10] + kernel[3][4] ~^ image[18][11] + kernel[4][0] ~^ image[19][7] + kernel[4][1] ~^ image[19][8] + kernel[4][2] ~^ image[19][9] + kernel[4][3] ~^ image[19][10] + kernel[4][4] ~^ image[19][11];
assign xor_sum[15][8] = kernel[0][0] ~^ image[15][8] + kernel[0][1] ~^ image[15][9] + kernel[0][2] ~^ image[15][10] + kernel[0][3] ~^ image[15][11] + kernel[0][4] ~^ image[15][12] + kernel[1][0] ~^ image[16][8] + kernel[1][1] ~^ image[16][9] + kernel[1][2] ~^ image[16][10] + kernel[1][3] ~^ image[16][11] + kernel[1][4] ~^ image[16][12] + kernel[2][0] ~^ image[17][8] + kernel[2][1] ~^ image[17][9] + kernel[2][2] ~^ image[17][10] + kernel[2][3] ~^ image[17][11] + kernel[2][4] ~^ image[17][12] + kernel[3][0] ~^ image[18][8] + kernel[3][1] ~^ image[18][9] + kernel[3][2] ~^ image[18][10] + kernel[3][3] ~^ image[18][11] + kernel[3][4] ~^ image[18][12] + kernel[4][0] ~^ image[19][8] + kernel[4][1] ~^ image[19][9] + kernel[4][2] ~^ image[19][10] + kernel[4][3] ~^ image[19][11] + kernel[4][4] ~^ image[19][12];
assign xor_sum[15][9] = kernel[0][0] ~^ image[15][9] + kernel[0][1] ~^ image[15][10] + kernel[0][2] ~^ image[15][11] + kernel[0][3] ~^ image[15][12] + kernel[0][4] ~^ image[15][13] + kernel[1][0] ~^ image[16][9] + kernel[1][1] ~^ image[16][10] + kernel[1][2] ~^ image[16][11] + kernel[1][3] ~^ image[16][12] + kernel[1][4] ~^ image[16][13] + kernel[2][0] ~^ image[17][9] + kernel[2][1] ~^ image[17][10] + kernel[2][2] ~^ image[17][11] + kernel[2][3] ~^ image[17][12] + kernel[2][4] ~^ image[17][13] + kernel[3][0] ~^ image[18][9] + kernel[3][1] ~^ image[18][10] + kernel[3][2] ~^ image[18][11] + kernel[3][3] ~^ image[18][12] + kernel[3][4] ~^ image[18][13] + kernel[4][0] ~^ image[19][9] + kernel[4][1] ~^ image[19][10] + kernel[4][2] ~^ image[19][11] + kernel[4][3] ~^ image[19][12] + kernel[4][4] ~^ image[19][13];
assign xor_sum[15][10] = kernel[0][0] ~^ image[15][10] + kernel[0][1] ~^ image[15][11] + kernel[0][2] ~^ image[15][12] + kernel[0][3] ~^ image[15][13] + kernel[0][4] ~^ image[15][14] + kernel[1][0] ~^ image[16][10] + kernel[1][1] ~^ image[16][11] + kernel[1][2] ~^ image[16][12] + kernel[1][3] ~^ image[16][13] + kernel[1][4] ~^ image[16][14] + kernel[2][0] ~^ image[17][10] + kernel[2][1] ~^ image[17][11] + kernel[2][2] ~^ image[17][12] + kernel[2][3] ~^ image[17][13] + kernel[2][4] ~^ image[17][14] + kernel[3][0] ~^ image[18][10] + kernel[3][1] ~^ image[18][11] + kernel[3][2] ~^ image[18][12] + kernel[3][3] ~^ image[18][13] + kernel[3][4] ~^ image[18][14] + kernel[4][0] ~^ image[19][10] + kernel[4][1] ~^ image[19][11] + kernel[4][2] ~^ image[19][12] + kernel[4][3] ~^ image[19][13] + kernel[4][4] ~^ image[19][14];
assign xor_sum[15][11] = kernel[0][0] ~^ image[15][11] + kernel[0][1] ~^ image[15][12] + kernel[0][2] ~^ image[15][13] + kernel[0][3] ~^ image[15][14] + kernel[0][4] ~^ image[15][15] + kernel[1][0] ~^ image[16][11] + kernel[1][1] ~^ image[16][12] + kernel[1][2] ~^ image[16][13] + kernel[1][3] ~^ image[16][14] + kernel[1][4] ~^ image[16][15] + kernel[2][0] ~^ image[17][11] + kernel[2][1] ~^ image[17][12] + kernel[2][2] ~^ image[17][13] + kernel[2][3] ~^ image[17][14] + kernel[2][4] ~^ image[17][15] + kernel[3][0] ~^ image[18][11] + kernel[3][1] ~^ image[18][12] + kernel[3][2] ~^ image[18][13] + kernel[3][3] ~^ image[18][14] + kernel[3][4] ~^ image[18][15] + kernel[4][0] ~^ image[19][11] + kernel[4][1] ~^ image[19][12] + kernel[4][2] ~^ image[19][13] + kernel[4][3] ~^ image[19][14] + kernel[4][4] ~^ image[19][15];
assign xor_sum[15][12] = kernel[0][0] ~^ image[15][12] + kernel[0][1] ~^ image[15][13] + kernel[0][2] ~^ image[15][14] + kernel[0][3] ~^ image[15][15] + kernel[0][4] ~^ image[15][16] + kernel[1][0] ~^ image[16][12] + kernel[1][1] ~^ image[16][13] + kernel[1][2] ~^ image[16][14] + kernel[1][3] ~^ image[16][15] + kernel[1][4] ~^ image[16][16] + kernel[2][0] ~^ image[17][12] + kernel[2][1] ~^ image[17][13] + kernel[2][2] ~^ image[17][14] + kernel[2][3] ~^ image[17][15] + kernel[2][4] ~^ image[17][16] + kernel[3][0] ~^ image[18][12] + kernel[3][1] ~^ image[18][13] + kernel[3][2] ~^ image[18][14] + kernel[3][3] ~^ image[18][15] + kernel[3][4] ~^ image[18][16] + kernel[4][0] ~^ image[19][12] + kernel[4][1] ~^ image[19][13] + kernel[4][2] ~^ image[19][14] + kernel[4][3] ~^ image[19][15] + kernel[4][4] ~^ image[19][16];
assign xor_sum[15][13] = kernel[0][0] ~^ image[15][13] + kernel[0][1] ~^ image[15][14] + kernel[0][2] ~^ image[15][15] + kernel[0][3] ~^ image[15][16] + kernel[0][4] ~^ image[15][17] + kernel[1][0] ~^ image[16][13] + kernel[1][1] ~^ image[16][14] + kernel[1][2] ~^ image[16][15] + kernel[1][3] ~^ image[16][16] + kernel[1][4] ~^ image[16][17] + kernel[2][0] ~^ image[17][13] + kernel[2][1] ~^ image[17][14] + kernel[2][2] ~^ image[17][15] + kernel[2][3] ~^ image[17][16] + kernel[2][4] ~^ image[17][17] + kernel[3][0] ~^ image[18][13] + kernel[3][1] ~^ image[18][14] + kernel[3][2] ~^ image[18][15] + kernel[3][3] ~^ image[18][16] + kernel[3][4] ~^ image[18][17] + kernel[4][0] ~^ image[19][13] + kernel[4][1] ~^ image[19][14] + kernel[4][2] ~^ image[19][15] + kernel[4][3] ~^ image[19][16] + kernel[4][4] ~^ image[19][17];
assign xor_sum[15][14] = kernel[0][0] ~^ image[15][14] + kernel[0][1] ~^ image[15][15] + kernel[0][2] ~^ image[15][16] + kernel[0][3] ~^ image[15][17] + kernel[0][4] ~^ image[15][18] + kernel[1][0] ~^ image[16][14] + kernel[1][1] ~^ image[16][15] + kernel[1][2] ~^ image[16][16] + kernel[1][3] ~^ image[16][17] + kernel[1][4] ~^ image[16][18] + kernel[2][0] ~^ image[17][14] + kernel[2][1] ~^ image[17][15] + kernel[2][2] ~^ image[17][16] + kernel[2][3] ~^ image[17][17] + kernel[2][4] ~^ image[17][18] + kernel[3][0] ~^ image[18][14] + kernel[3][1] ~^ image[18][15] + kernel[3][2] ~^ image[18][16] + kernel[3][3] ~^ image[18][17] + kernel[3][4] ~^ image[18][18] + kernel[4][0] ~^ image[19][14] + kernel[4][1] ~^ image[19][15] + kernel[4][2] ~^ image[19][16] + kernel[4][3] ~^ image[19][17] + kernel[4][4] ~^ image[19][18];
assign xor_sum[15][15] = kernel[0][0] ~^ image[15][15] + kernel[0][1] ~^ image[15][16] + kernel[0][2] ~^ image[15][17] + kernel[0][3] ~^ image[15][18] + kernel[0][4] ~^ image[15][19] + kernel[1][0] ~^ image[16][15] + kernel[1][1] ~^ image[16][16] + kernel[1][2] ~^ image[16][17] + kernel[1][3] ~^ image[16][18] + kernel[1][4] ~^ image[16][19] + kernel[2][0] ~^ image[17][15] + kernel[2][1] ~^ image[17][16] + kernel[2][2] ~^ image[17][17] + kernel[2][3] ~^ image[17][18] + kernel[2][4] ~^ image[17][19] + kernel[3][0] ~^ image[18][15] + kernel[3][1] ~^ image[18][16] + kernel[3][2] ~^ image[18][17] + kernel[3][3] ~^ image[18][18] + kernel[3][4] ~^ image[18][19] + kernel[4][0] ~^ image[19][15] + kernel[4][1] ~^ image[19][16] + kernel[4][2] ~^ image[19][17] + kernel[4][3] ~^ image[19][18] + kernel[4][4] ~^ image[19][19];
assign xor_sum[15][16] = kernel[0][0] ~^ image[15][16] + kernel[0][1] ~^ image[15][17] + kernel[0][2] ~^ image[15][18] + kernel[0][3] ~^ image[15][19] + kernel[0][4] ~^ image[15][20] + kernel[1][0] ~^ image[16][16] + kernel[1][1] ~^ image[16][17] + kernel[1][2] ~^ image[16][18] + kernel[1][3] ~^ image[16][19] + kernel[1][4] ~^ image[16][20] + kernel[2][0] ~^ image[17][16] + kernel[2][1] ~^ image[17][17] + kernel[2][2] ~^ image[17][18] + kernel[2][3] ~^ image[17][19] + kernel[2][4] ~^ image[17][20] + kernel[3][0] ~^ image[18][16] + kernel[3][1] ~^ image[18][17] + kernel[3][2] ~^ image[18][18] + kernel[3][3] ~^ image[18][19] + kernel[3][4] ~^ image[18][20] + kernel[4][0] ~^ image[19][16] + kernel[4][1] ~^ image[19][17] + kernel[4][2] ~^ image[19][18] + kernel[4][3] ~^ image[19][19] + kernel[4][4] ~^ image[19][20];
assign xor_sum[15][17] = kernel[0][0] ~^ image[15][17] + kernel[0][1] ~^ image[15][18] + kernel[0][2] ~^ image[15][19] + kernel[0][3] ~^ image[15][20] + kernel[0][4] ~^ image[15][21] + kernel[1][0] ~^ image[16][17] + kernel[1][1] ~^ image[16][18] + kernel[1][2] ~^ image[16][19] + kernel[1][3] ~^ image[16][20] + kernel[1][4] ~^ image[16][21] + kernel[2][0] ~^ image[17][17] + kernel[2][1] ~^ image[17][18] + kernel[2][2] ~^ image[17][19] + kernel[2][3] ~^ image[17][20] + kernel[2][4] ~^ image[17][21] + kernel[3][0] ~^ image[18][17] + kernel[3][1] ~^ image[18][18] + kernel[3][2] ~^ image[18][19] + kernel[3][3] ~^ image[18][20] + kernel[3][4] ~^ image[18][21] + kernel[4][0] ~^ image[19][17] + kernel[4][1] ~^ image[19][18] + kernel[4][2] ~^ image[19][19] + kernel[4][3] ~^ image[19][20] + kernel[4][4] ~^ image[19][21];
assign xor_sum[15][18] = kernel[0][0] ~^ image[15][18] + kernel[0][1] ~^ image[15][19] + kernel[0][2] ~^ image[15][20] + kernel[0][3] ~^ image[15][21] + kernel[0][4] ~^ image[15][22] + kernel[1][0] ~^ image[16][18] + kernel[1][1] ~^ image[16][19] + kernel[1][2] ~^ image[16][20] + kernel[1][3] ~^ image[16][21] + kernel[1][4] ~^ image[16][22] + kernel[2][0] ~^ image[17][18] + kernel[2][1] ~^ image[17][19] + kernel[2][2] ~^ image[17][20] + kernel[2][3] ~^ image[17][21] + kernel[2][4] ~^ image[17][22] + kernel[3][0] ~^ image[18][18] + kernel[3][1] ~^ image[18][19] + kernel[3][2] ~^ image[18][20] + kernel[3][3] ~^ image[18][21] + kernel[3][4] ~^ image[18][22] + kernel[4][0] ~^ image[19][18] + kernel[4][1] ~^ image[19][19] + kernel[4][2] ~^ image[19][20] + kernel[4][3] ~^ image[19][21] + kernel[4][4] ~^ image[19][22];
assign xor_sum[15][19] = kernel[0][0] ~^ image[15][19] + kernel[0][1] ~^ image[15][20] + kernel[0][2] ~^ image[15][21] + kernel[0][3] ~^ image[15][22] + kernel[0][4] ~^ image[15][23] + kernel[1][0] ~^ image[16][19] + kernel[1][1] ~^ image[16][20] + kernel[1][2] ~^ image[16][21] + kernel[1][3] ~^ image[16][22] + kernel[1][4] ~^ image[16][23] + kernel[2][0] ~^ image[17][19] + kernel[2][1] ~^ image[17][20] + kernel[2][2] ~^ image[17][21] + kernel[2][3] ~^ image[17][22] + kernel[2][4] ~^ image[17][23] + kernel[3][0] ~^ image[18][19] + kernel[3][1] ~^ image[18][20] + kernel[3][2] ~^ image[18][21] + kernel[3][3] ~^ image[18][22] + kernel[3][4] ~^ image[18][23] + kernel[4][0] ~^ image[19][19] + kernel[4][1] ~^ image[19][20] + kernel[4][2] ~^ image[19][21] + kernel[4][3] ~^ image[19][22] + kernel[4][4] ~^ image[19][23];
assign xor_sum[15][20] = kernel[0][0] ~^ image[15][20] + kernel[0][1] ~^ image[15][21] + kernel[0][2] ~^ image[15][22] + kernel[0][3] ~^ image[15][23] + kernel[0][4] ~^ image[15][24] + kernel[1][0] ~^ image[16][20] + kernel[1][1] ~^ image[16][21] + kernel[1][2] ~^ image[16][22] + kernel[1][3] ~^ image[16][23] + kernel[1][4] ~^ image[16][24] + kernel[2][0] ~^ image[17][20] + kernel[2][1] ~^ image[17][21] + kernel[2][2] ~^ image[17][22] + kernel[2][3] ~^ image[17][23] + kernel[2][4] ~^ image[17][24] + kernel[3][0] ~^ image[18][20] + kernel[3][1] ~^ image[18][21] + kernel[3][2] ~^ image[18][22] + kernel[3][3] ~^ image[18][23] + kernel[3][4] ~^ image[18][24] + kernel[4][0] ~^ image[19][20] + kernel[4][1] ~^ image[19][21] + kernel[4][2] ~^ image[19][22] + kernel[4][3] ~^ image[19][23] + kernel[4][4] ~^ image[19][24];
assign xor_sum[15][21] = kernel[0][0] ~^ image[15][21] + kernel[0][1] ~^ image[15][22] + kernel[0][2] ~^ image[15][23] + kernel[0][3] ~^ image[15][24] + kernel[0][4] ~^ image[15][25] + kernel[1][0] ~^ image[16][21] + kernel[1][1] ~^ image[16][22] + kernel[1][2] ~^ image[16][23] + kernel[1][3] ~^ image[16][24] + kernel[1][4] ~^ image[16][25] + kernel[2][0] ~^ image[17][21] + kernel[2][1] ~^ image[17][22] + kernel[2][2] ~^ image[17][23] + kernel[2][3] ~^ image[17][24] + kernel[2][4] ~^ image[17][25] + kernel[3][0] ~^ image[18][21] + kernel[3][1] ~^ image[18][22] + kernel[3][2] ~^ image[18][23] + kernel[3][3] ~^ image[18][24] + kernel[3][4] ~^ image[18][25] + kernel[4][0] ~^ image[19][21] + kernel[4][1] ~^ image[19][22] + kernel[4][2] ~^ image[19][23] + kernel[4][3] ~^ image[19][24] + kernel[4][4] ~^ image[19][25];
assign xor_sum[15][22] = kernel[0][0] ~^ image[15][22] + kernel[0][1] ~^ image[15][23] + kernel[0][2] ~^ image[15][24] + kernel[0][3] ~^ image[15][25] + kernel[0][4] ~^ image[15][26] + kernel[1][0] ~^ image[16][22] + kernel[1][1] ~^ image[16][23] + kernel[1][2] ~^ image[16][24] + kernel[1][3] ~^ image[16][25] + kernel[1][4] ~^ image[16][26] + kernel[2][0] ~^ image[17][22] + kernel[2][1] ~^ image[17][23] + kernel[2][2] ~^ image[17][24] + kernel[2][3] ~^ image[17][25] + kernel[2][4] ~^ image[17][26] + kernel[3][0] ~^ image[18][22] + kernel[3][1] ~^ image[18][23] + kernel[3][2] ~^ image[18][24] + kernel[3][3] ~^ image[18][25] + kernel[3][4] ~^ image[18][26] + kernel[4][0] ~^ image[19][22] + kernel[4][1] ~^ image[19][23] + kernel[4][2] ~^ image[19][24] + kernel[4][3] ~^ image[19][25] + kernel[4][4] ~^ image[19][26];
assign xor_sum[15][23] = kernel[0][0] ~^ image[15][23] + kernel[0][1] ~^ image[15][24] + kernel[0][2] ~^ image[15][25] + kernel[0][3] ~^ image[15][26] + kernel[0][4] ~^ image[15][27] + kernel[1][0] ~^ image[16][23] + kernel[1][1] ~^ image[16][24] + kernel[1][2] ~^ image[16][25] + kernel[1][3] ~^ image[16][26] + kernel[1][4] ~^ image[16][27] + kernel[2][0] ~^ image[17][23] + kernel[2][1] ~^ image[17][24] + kernel[2][2] ~^ image[17][25] + kernel[2][3] ~^ image[17][26] + kernel[2][4] ~^ image[17][27] + kernel[3][0] ~^ image[18][23] + kernel[3][1] ~^ image[18][24] + kernel[3][2] ~^ image[18][25] + kernel[3][3] ~^ image[18][26] + kernel[3][4] ~^ image[18][27] + kernel[4][0] ~^ image[19][23] + kernel[4][1] ~^ image[19][24] + kernel[4][2] ~^ image[19][25] + kernel[4][3] ~^ image[19][26] + kernel[4][4] ~^ image[19][27];
assign xor_sum[16][0] = kernel[0][0] ~^ image[16][0] + kernel[0][1] ~^ image[16][1] + kernel[0][2] ~^ image[16][2] + kernel[0][3] ~^ image[16][3] + kernel[0][4] ~^ image[16][4] + kernel[1][0] ~^ image[17][0] + kernel[1][1] ~^ image[17][1] + kernel[1][2] ~^ image[17][2] + kernel[1][3] ~^ image[17][3] + kernel[1][4] ~^ image[17][4] + kernel[2][0] ~^ image[18][0] + kernel[2][1] ~^ image[18][1] + kernel[2][2] ~^ image[18][2] + kernel[2][3] ~^ image[18][3] + kernel[2][4] ~^ image[18][4] + kernel[3][0] ~^ image[19][0] + kernel[3][1] ~^ image[19][1] + kernel[3][2] ~^ image[19][2] + kernel[3][3] ~^ image[19][3] + kernel[3][4] ~^ image[19][4] + kernel[4][0] ~^ image[20][0] + kernel[4][1] ~^ image[20][1] + kernel[4][2] ~^ image[20][2] + kernel[4][3] ~^ image[20][3] + kernel[4][4] ~^ image[20][4];
assign xor_sum[16][1] = kernel[0][0] ~^ image[16][1] + kernel[0][1] ~^ image[16][2] + kernel[0][2] ~^ image[16][3] + kernel[0][3] ~^ image[16][4] + kernel[0][4] ~^ image[16][5] + kernel[1][0] ~^ image[17][1] + kernel[1][1] ~^ image[17][2] + kernel[1][2] ~^ image[17][3] + kernel[1][3] ~^ image[17][4] + kernel[1][4] ~^ image[17][5] + kernel[2][0] ~^ image[18][1] + kernel[2][1] ~^ image[18][2] + kernel[2][2] ~^ image[18][3] + kernel[2][3] ~^ image[18][4] + kernel[2][4] ~^ image[18][5] + kernel[3][0] ~^ image[19][1] + kernel[3][1] ~^ image[19][2] + kernel[3][2] ~^ image[19][3] + kernel[3][3] ~^ image[19][4] + kernel[3][4] ~^ image[19][5] + kernel[4][0] ~^ image[20][1] + kernel[4][1] ~^ image[20][2] + kernel[4][2] ~^ image[20][3] + kernel[4][3] ~^ image[20][4] + kernel[4][4] ~^ image[20][5];
assign xor_sum[16][2] = kernel[0][0] ~^ image[16][2] + kernel[0][1] ~^ image[16][3] + kernel[0][2] ~^ image[16][4] + kernel[0][3] ~^ image[16][5] + kernel[0][4] ~^ image[16][6] + kernel[1][0] ~^ image[17][2] + kernel[1][1] ~^ image[17][3] + kernel[1][2] ~^ image[17][4] + kernel[1][3] ~^ image[17][5] + kernel[1][4] ~^ image[17][6] + kernel[2][0] ~^ image[18][2] + kernel[2][1] ~^ image[18][3] + kernel[2][2] ~^ image[18][4] + kernel[2][3] ~^ image[18][5] + kernel[2][4] ~^ image[18][6] + kernel[3][0] ~^ image[19][2] + kernel[3][1] ~^ image[19][3] + kernel[3][2] ~^ image[19][4] + kernel[3][3] ~^ image[19][5] + kernel[3][4] ~^ image[19][6] + kernel[4][0] ~^ image[20][2] + kernel[4][1] ~^ image[20][3] + kernel[4][2] ~^ image[20][4] + kernel[4][3] ~^ image[20][5] + kernel[4][4] ~^ image[20][6];
assign xor_sum[16][3] = kernel[0][0] ~^ image[16][3] + kernel[0][1] ~^ image[16][4] + kernel[0][2] ~^ image[16][5] + kernel[0][3] ~^ image[16][6] + kernel[0][4] ~^ image[16][7] + kernel[1][0] ~^ image[17][3] + kernel[1][1] ~^ image[17][4] + kernel[1][2] ~^ image[17][5] + kernel[1][3] ~^ image[17][6] + kernel[1][4] ~^ image[17][7] + kernel[2][0] ~^ image[18][3] + kernel[2][1] ~^ image[18][4] + kernel[2][2] ~^ image[18][5] + kernel[2][3] ~^ image[18][6] + kernel[2][4] ~^ image[18][7] + kernel[3][0] ~^ image[19][3] + kernel[3][1] ~^ image[19][4] + kernel[3][2] ~^ image[19][5] + kernel[3][3] ~^ image[19][6] + kernel[3][4] ~^ image[19][7] + kernel[4][0] ~^ image[20][3] + kernel[4][1] ~^ image[20][4] + kernel[4][2] ~^ image[20][5] + kernel[4][3] ~^ image[20][6] + kernel[4][4] ~^ image[20][7];
assign xor_sum[16][4] = kernel[0][0] ~^ image[16][4] + kernel[0][1] ~^ image[16][5] + kernel[0][2] ~^ image[16][6] + kernel[0][3] ~^ image[16][7] + kernel[0][4] ~^ image[16][8] + kernel[1][0] ~^ image[17][4] + kernel[1][1] ~^ image[17][5] + kernel[1][2] ~^ image[17][6] + kernel[1][3] ~^ image[17][7] + kernel[1][4] ~^ image[17][8] + kernel[2][0] ~^ image[18][4] + kernel[2][1] ~^ image[18][5] + kernel[2][2] ~^ image[18][6] + kernel[2][3] ~^ image[18][7] + kernel[2][4] ~^ image[18][8] + kernel[3][0] ~^ image[19][4] + kernel[3][1] ~^ image[19][5] + kernel[3][2] ~^ image[19][6] + kernel[3][3] ~^ image[19][7] + kernel[3][4] ~^ image[19][8] + kernel[4][0] ~^ image[20][4] + kernel[4][1] ~^ image[20][5] + kernel[4][2] ~^ image[20][6] + kernel[4][3] ~^ image[20][7] + kernel[4][4] ~^ image[20][8];
assign xor_sum[16][5] = kernel[0][0] ~^ image[16][5] + kernel[0][1] ~^ image[16][6] + kernel[0][2] ~^ image[16][7] + kernel[0][3] ~^ image[16][8] + kernel[0][4] ~^ image[16][9] + kernel[1][0] ~^ image[17][5] + kernel[1][1] ~^ image[17][6] + kernel[1][2] ~^ image[17][7] + kernel[1][3] ~^ image[17][8] + kernel[1][4] ~^ image[17][9] + kernel[2][0] ~^ image[18][5] + kernel[2][1] ~^ image[18][6] + kernel[2][2] ~^ image[18][7] + kernel[2][3] ~^ image[18][8] + kernel[2][4] ~^ image[18][9] + kernel[3][0] ~^ image[19][5] + kernel[3][1] ~^ image[19][6] + kernel[3][2] ~^ image[19][7] + kernel[3][3] ~^ image[19][8] + kernel[3][4] ~^ image[19][9] + kernel[4][0] ~^ image[20][5] + kernel[4][1] ~^ image[20][6] + kernel[4][2] ~^ image[20][7] + kernel[4][3] ~^ image[20][8] + kernel[4][4] ~^ image[20][9];
assign xor_sum[16][6] = kernel[0][0] ~^ image[16][6] + kernel[0][1] ~^ image[16][7] + kernel[0][2] ~^ image[16][8] + kernel[0][3] ~^ image[16][9] + kernel[0][4] ~^ image[16][10] + kernel[1][0] ~^ image[17][6] + kernel[1][1] ~^ image[17][7] + kernel[1][2] ~^ image[17][8] + kernel[1][3] ~^ image[17][9] + kernel[1][4] ~^ image[17][10] + kernel[2][0] ~^ image[18][6] + kernel[2][1] ~^ image[18][7] + kernel[2][2] ~^ image[18][8] + kernel[2][3] ~^ image[18][9] + kernel[2][4] ~^ image[18][10] + kernel[3][0] ~^ image[19][6] + kernel[3][1] ~^ image[19][7] + kernel[3][2] ~^ image[19][8] + kernel[3][3] ~^ image[19][9] + kernel[3][4] ~^ image[19][10] + kernel[4][0] ~^ image[20][6] + kernel[4][1] ~^ image[20][7] + kernel[4][2] ~^ image[20][8] + kernel[4][3] ~^ image[20][9] + kernel[4][4] ~^ image[20][10];
assign xor_sum[16][7] = kernel[0][0] ~^ image[16][7] + kernel[0][1] ~^ image[16][8] + kernel[0][2] ~^ image[16][9] + kernel[0][3] ~^ image[16][10] + kernel[0][4] ~^ image[16][11] + kernel[1][0] ~^ image[17][7] + kernel[1][1] ~^ image[17][8] + kernel[1][2] ~^ image[17][9] + kernel[1][3] ~^ image[17][10] + kernel[1][4] ~^ image[17][11] + kernel[2][0] ~^ image[18][7] + kernel[2][1] ~^ image[18][8] + kernel[2][2] ~^ image[18][9] + kernel[2][3] ~^ image[18][10] + kernel[2][4] ~^ image[18][11] + kernel[3][0] ~^ image[19][7] + kernel[3][1] ~^ image[19][8] + kernel[3][2] ~^ image[19][9] + kernel[3][3] ~^ image[19][10] + kernel[3][4] ~^ image[19][11] + kernel[4][0] ~^ image[20][7] + kernel[4][1] ~^ image[20][8] + kernel[4][2] ~^ image[20][9] + kernel[4][3] ~^ image[20][10] + kernel[4][4] ~^ image[20][11];
assign xor_sum[16][8] = kernel[0][0] ~^ image[16][8] + kernel[0][1] ~^ image[16][9] + kernel[0][2] ~^ image[16][10] + kernel[0][3] ~^ image[16][11] + kernel[0][4] ~^ image[16][12] + kernel[1][0] ~^ image[17][8] + kernel[1][1] ~^ image[17][9] + kernel[1][2] ~^ image[17][10] + kernel[1][3] ~^ image[17][11] + kernel[1][4] ~^ image[17][12] + kernel[2][0] ~^ image[18][8] + kernel[2][1] ~^ image[18][9] + kernel[2][2] ~^ image[18][10] + kernel[2][3] ~^ image[18][11] + kernel[2][4] ~^ image[18][12] + kernel[3][0] ~^ image[19][8] + kernel[3][1] ~^ image[19][9] + kernel[3][2] ~^ image[19][10] + kernel[3][3] ~^ image[19][11] + kernel[3][4] ~^ image[19][12] + kernel[4][0] ~^ image[20][8] + kernel[4][1] ~^ image[20][9] + kernel[4][2] ~^ image[20][10] + kernel[4][3] ~^ image[20][11] + kernel[4][4] ~^ image[20][12];
assign xor_sum[16][9] = kernel[0][0] ~^ image[16][9] + kernel[0][1] ~^ image[16][10] + kernel[0][2] ~^ image[16][11] + kernel[0][3] ~^ image[16][12] + kernel[0][4] ~^ image[16][13] + kernel[1][0] ~^ image[17][9] + kernel[1][1] ~^ image[17][10] + kernel[1][2] ~^ image[17][11] + kernel[1][3] ~^ image[17][12] + kernel[1][4] ~^ image[17][13] + kernel[2][0] ~^ image[18][9] + kernel[2][1] ~^ image[18][10] + kernel[2][2] ~^ image[18][11] + kernel[2][3] ~^ image[18][12] + kernel[2][4] ~^ image[18][13] + kernel[3][0] ~^ image[19][9] + kernel[3][1] ~^ image[19][10] + kernel[3][2] ~^ image[19][11] + kernel[3][3] ~^ image[19][12] + kernel[3][4] ~^ image[19][13] + kernel[4][0] ~^ image[20][9] + kernel[4][1] ~^ image[20][10] + kernel[4][2] ~^ image[20][11] + kernel[4][3] ~^ image[20][12] + kernel[4][4] ~^ image[20][13];
assign xor_sum[16][10] = kernel[0][0] ~^ image[16][10] + kernel[0][1] ~^ image[16][11] + kernel[0][2] ~^ image[16][12] + kernel[0][3] ~^ image[16][13] + kernel[0][4] ~^ image[16][14] + kernel[1][0] ~^ image[17][10] + kernel[1][1] ~^ image[17][11] + kernel[1][2] ~^ image[17][12] + kernel[1][3] ~^ image[17][13] + kernel[1][4] ~^ image[17][14] + kernel[2][0] ~^ image[18][10] + kernel[2][1] ~^ image[18][11] + kernel[2][2] ~^ image[18][12] + kernel[2][3] ~^ image[18][13] + kernel[2][4] ~^ image[18][14] + kernel[3][0] ~^ image[19][10] + kernel[3][1] ~^ image[19][11] + kernel[3][2] ~^ image[19][12] + kernel[3][3] ~^ image[19][13] + kernel[3][4] ~^ image[19][14] + kernel[4][0] ~^ image[20][10] + kernel[4][1] ~^ image[20][11] + kernel[4][2] ~^ image[20][12] + kernel[4][3] ~^ image[20][13] + kernel[4][4] ~^ image[20][14];
assign xor_sum[16][11] = kernel[0][0] ~^ image[16][11] + kernel[0][1] ~^ image[16][12] + kernel[0][2] ~^ image[16][13] + kernel[0][3] ~^ image[16][14] + kernel[0][4] ~^ image[16][15] + kernel[1][0] ~^ image[17][11] + kernel[1][1] ~^ image[17][12] + kernel[1][2] ~^ image[17][13] + kernel[1][3] ~^ image[17][14] + kernel[1][4] ~^ image[17][15] + kernel[2][0] ~^ image[18][11] + kernel[2][1] ~^ image[18][12] + kernel[2][2] ~^ image[18][13] + kernel[2][3] ~^ image[18][14] + kernel[2][4] ~^ image[18][15] + kernel[3][0] ~^ image[19][11] + kernel[3][1] ~^ image[19][12] + kernel[3][2] ~^ image[19][13] + kernel[3][3] ~^ image[19][14] + kernel[3][4] ~^ image[19][15] + kernel[4][0] ~^ image[20][11] + kernel[4][1] ~^ image[20][12] + kernel[4][2] ~^ image[20][13] + kernel[4][3] ~^ image[20][14] + kernel[4][4] ~^ image[20][15];
assign xor_sum[16][12] = kernel[0][0] ~^ image[16][12] + kernel[0][1] ~^ image[16][13] + kernel[0][2] ~^ image[16][14] + kernel[0][3] ~^ image[16][15] + kernel[0][4] ~^ image[16][16] + kernel[1][0] ~^ image[17][12] + kernel[1][1] ~^ image[17][13] + kernel[1][2] ~^ image[17][14] + kernel[1][3] ~^ image[17][15] + kernel[1][4] ~^ image[17][16] + kernel[2][0] ~^ image[18][12] + kernel[2][1] ~^ image[18][13] + kernel[2][2] ~^ image[18][14] + kernel[2][3] ~^ image[18][15] + kernel[2][4] ~^ image[18][16] + kernel[3][0] ~^ image[19][12] + kernel[3][1] ~^ image[19][13] + kernel[3][2] ~^ image[19][14] + kernel[3][3] ~^ image[19][15] + kernel[3][4] ~^ image[19][16] + kernel[4][0] ~^ image[20][12] + kernel[4][1] ~^ image[20][13] + kernel[4][2] ~^ image[20][14] + kernel[4][3] ~^ image[20][15] + kernel[4][4] ~^ image[20][16];
assign xor_sum[16][13] = kernel[0][0] ~^ image[16][13] + kernel[0][1] ~^ image[16][14] + kernel[0][2] ~^ image[16][15] + kernel[0][3] ~^ image[16][16] + kernel[0][4] ~^ image[16][17] + kernel[1][0] ~^ image[17][13] + kernel[1][1] ~^ image[17][14] + kernel[1][2] ~^ image[17][15] + kernel[1][3] ~^ image[17][16] + kernel[1][4] ~^ image[17][17] + kernel[2][0] ~^ image[18][13] + kernel[2][1] ~^ image[18][14] + kernel[2][2] ~^ image[18][15] + kernel[2][3] ~^ image[18][16] + kernel[2][4] ~^ image[18][17] + kernel[3][0] ~^ image[19][13] + kernel[3][1] ~^ image[19][14] + kernel[3][2] ~^ image[19][15] + kernel[3][3] ~^ image[19][16] + kernel[3][4] ~^ image[19][17] + kernel[4][0] ~^ image[20][13] + kernel[4][1] ~^ image[20][14] + kernel[4][2] ~^ image[20][15] + kernel[4][3] ~^ image[20][16] + kernel[4][4] ~^ image[20][17];
assign xor_sum[16][14] = kernel[0][0] ~^ image[16][14] + kernel[0][1] ~^ image[16][15] + kernel[0][2] ~^ image[16][16] + kernel[0][3] ~^ image[16][17] + kernel[0][4] ~^ image[16][18] + kernel[1][0] ~^ image[17][14] + kernel[1][1] ~^ image[17][15] + kernel[1][2] ~^ image[17][16] + kernel[1][3] ~^ image[17][17] + kernel[1][4] ~^ image[17][18] + kernel[2][0] ~^ image[18][14] + kernel[2][1] ~^ image[18][15] + kernel[2][2] ~^ image[18][16] + kernel[2][3] ~^ image[18][17] + kernel[2][4] ~^ image[18][18] + kernel[3][0] ~^ image[19][14] + kernel[3][1] ~^ image[19][15] + kernel[3][2] ~^ image[19][16] + kernel[3][3] ~^ image[19][17] + kernel[3][4] ~^ image[19][18] + kernel[4][0] ~^ image[20][14] + kernel[4][1] ~^ image[20][15] + kernel[4][2] ~^ image[20][16] + kernel[4][3] ~^ image[20][17] + kernel[4][4] ~^ image[20][18];
assign xor_sum[16][15] = kernel[0][0] ~^ image[16][15] + kernel[0][1] ~^ image[16][16] + kernel[0][2] ~^ image[16][17] + kernel[0][3] ~^ image[16][18] + kernel[0][4] ~^ image[16][19] + kernel[1][0] ~^ image[17][15] + kernel[1][1] ~^ image[17][16] + kernel[1][2] ~^ image[17][17] + kernel[1][3] ~^ image[17][18] + kernel[1][4] ~^ image[17][19] + kernel[2][0] ~^ image[18][15] + kernel[2][1] ~^ image[18][16] + kernel[2][2] ~^ image[18][17] + kernel[2][3] ~^ image[18][18] + kernel[2][4] ~^ image[18][19] + kernel[3][0] ~^ image[19][15] + kernel[3][1] ~^ image[19][16] + kernel[3][2] ~^ image[19][17] + kernel[3][3] ~^ image[19][18] + kernel[3][4] ~^ image[19][19] + kernel[4][0] ~^ image[20][15] + kernel[4][1] ~^ image[20][16] + kernel[4][2] ~^ image[20][17] + kernel[4][3] ~^ image[20][18] + kernel[4][4] ~^ image[20][19];
assign xor_sum[16][16] = kernel[0][0] ~^ image[16][16] + kernel[0][1] ~^ image[16][17] + kernel[0][2] ~^ image[16][18] + kernel[0][3] ~^ image[16][19] + kernel[0][4] ~^ image[16][20] + kernel[1][0] ~^ image[17][16] + kernel[1][1] ~^ image[17][17] + kernel[1][2] ~^ image[17][18] + kernel[1][3] ~^ image[17][19] + kernel[1][4] ~^ image[17][20] + kernel[2][0] ~^ image[18][16] + kernel[2][1] ~^ image[18][17] + kernel[2][2] ~^ image[18][18] + kernel[2][3] ~^ image[18][19] + kernel[2][4] ~^ image[18][20] + kernel[3][0] ~^ image[19][16] + kernel[3][1] ~^ image[19][17] + kernel[3][2] ~^ image[19][18] + kernel[3][3] ~^ image[19][19] + kernel[3][4] ~^ image[19][20] + kernel[4][0] ~^ image[20][16] + kernel[4][1] ~^ image[20][17] + kernel[4][2] ~^ image[20][18] + kernel[4][3] ~^ image[20][19] + kernel[4][4] ~^ image[20][20];
assign xor_sum[16][17] = kernel[0][0] ~^ image[16][17] + kernel[0][1] ~^ image[16][18] + kernel[0][2] ~^ image[16][19] + kernel[0][3] ~^ image[16][20] + kernel[0][4] ~^ image[16][21] + kernel[1][0] ~^ image[17][17] + kernel[1][1] ~^ image[17][18] + kernel[1][2] ~^ image[17][19] + kernel[1][3] ~^ image[17][20] + kernel[1][4] ~^ image[17][21] + kernel[2][0] ~^ image[18][17] + kernel[2][1] ~^ image[18][18] + kernel[2][2] ~^ image[18][19] + kernel[2][3] ~^ image[18][20] + kernel[2][4] ~^ image[18][21] + kernel[3][0] ~^ image[19][17] + kernel[3][1] ~^ image[19][18] + kernel[3][2] ~^ image[19][19] + kernel[3][3] ~^ image[19][20] + kernel[3][4] ~^ image[19][21] + kernel[4][0] ~^ image[20][17] + kernel[4][1] ~^ image[20][18] + kernel[4][2] ~^ image[20][19] + kernel[4][3] ~^ image[20][20] + kernel[4][4] ~^ image[20][21];
assign xor_sum[16][18] = kernel[0][0] ~^ image[16][18] + kernel[0][1] ~^ image[16][19] + kernel[0][2] ~^ image[16][20] + kernel[0][3] ~^ image[16][21] + kernel[0][4] ~^ image[16][22] + kernel[1][0] ~^ image[17][18] + kernel[1][1] ~^ image[17][19] + kernel[1][2] ~^ image[17][20] + kernel[1][3] ~^ image[17][21] + kernel[1][4] ~^ image[17][22] + kernel[2][0] ~^ image[18][18] + kernel[2][1] ~^ image[18][19] + kernel[2][2] ~^ image[18][20] + kernel[2][3] ~^ image[18][21] + kernel[2][4] ~^ image[18][22] + kernel[3][0] ~^ image[19][18] + kernel[3][1] ~^ image[19][19] + kernel[3][2] ~^ image[19][20] + kernel[3][3] ~^ image[19][21] + kernel[3][4] ~^ image[19][22] + kernel[4][0] ~^ image[20][18] + kernel[4][1] ~^ image[20][19] + kernel[4][2] ~^ image[20][20] + kernel[4][3] ~^ image[20][21] + kernel[4][4] ~^ image[20][22];
assign xor_sum[16][19] = kernel[0][0] ~^ image[16][19] + kernel[0][1] ~^ image[16][20] + kernel[0][2] ~^ image[16][21] + kernel[0][3] ~^ image[16][22] + kernel[0][4] ~^ image[16][23] + kernel[1][0] ~^ image[17][19] + kernel[1][1] ~^ image[17][20] + kernel[1][2] ~^ image[17][21] + kernel[1][3] ~^ image[17][22] + kernel[1][4] ~^ image[17][23] + kernel[2][0] ~^ image[18][19] + kernel[2][1] ~^ image[18][20] + kernel[2][2] ~^ image[18][21] + kernel[2][3] ~^ image[18][22] + kernel[2][4] ~^ image[18][23] + kernel[3][0] ~^ image[19][19] + kernel[3][1] ~^ image[19][20] + kernel[3][2] ~^ image[19][21] + kernel[3][3] ~^ image[19][22] + kernel[3][4] ~^ image[19][23] + kernel[4][0] ~^ image[20][19] + kernel[4][1] ~^ image[20][20] + kernel[4][2] ~^ image[20][21] + kernel[4][3] ~^ image[20][22] + kernel[4][4] ~^ image[20][23];
assign xor_sum[16][20] = kernel[0][0] ~^ image[16][20] + kernel[0][1] ~^ image[16][21] + kernel[0][2] ~^ image[16][22] + kernel[0][3] ~^ image[16][23] + kernel[0][4] ~^ image[16][24] + kernel[1][0] ~^ image[17][20] + kernel[1][1] ~^ image[17][21] + kernel[1][2] ~^ image[17][22] + kernel[1][3] ~^ image[17][23] + kernel[1][4] ~^ image[17][24] + kernel[2][0] ~^ image[18][20] + kernel[2][1] ~^ image[18][21] + kernel[2][2] ~^ image[18][22] + kernel[2][3] ~^ image[18][23] + kernel[2][4] ~^ image[18][24] + kernel[3][0] ~^ image[19][20] + kernel[3][1] ~^ image[19][21] + kernel[3][2] ~^ image[19][22] + kernel[3][3] ~^ image[19][23] + kernel[3][4] ~^ image[19][24] + kernel[4][0] ~^ image[20][20] + kernel[4][1] ~^ image[20][21] + kernel[4][2] ~^ image[20][22] + kernel[4][3] ~^ image[20][23] + kernel[4][4] ~^ image[20][24];
assign xor_sum[16][21] = kernel[0][0] ~^ image[16][21] + kernel[0][1] ~^ image[16][22] + kernel[0][2] ~^ image[16][23] + kernel[0][3] ~^ image[16][24] + kernel[0][4] ~^ image[16][25] + kernel[1][0] ~^ image[17][21] + kernel[1][1] ~^ image[17][22] + kernel[1][2] ~^ image[17][23] + kernel[1][3] ~^ image[17][24] + kernel[1][4] ~^ image[17][25] + kernel[2][0] ~^ image[18][21] + kernel[2][1] ~^ image[18][22] + kernel[2][2] ~^ image[18][23] + kernel[2][3] ~^ image[18][24] + kernel[2][4] ~^ image[18][25] + kernel[3][0] ~^ image[19][21] + kernel[3][1] ~^ image[19][22] + kernel[3][2] ~^ image[19][23] + kernel[3][3] ~^ image[19][24] + kernel[3][4] ~^ image[19][25] + kernel[4][0] ~^ image[20][21] + kernel[4][1] ~^ image[20][22] + kernel[4][2] ~^ image[20][23] + kernel[4][3] ~^ image[20][24] + kernel[4][4] ~^ image[20][25];
assign xor_sum[16][22] = kernel[0][0] ~^ image[16][22] + kernel[0][1] ~^ image[16][23] + kernel[0][2] ~^ image[16][24] + kernel[0][3] ~^ image[16][25] + kernel[0][4] ~^ image[16][26] + kernel[1][0] ~^ image[17][22] + kernel[1][1] ~^ image[17][23] + kernel[1][2] ~^ image[17][24] + kernel[1][3] ~^ image[17][25] + kernel[1][4] ~^ image[17][26] + kernel[2][0] ~^ image[18][22] + kernel[2][1] ~^ image[18][23] + kernel[2][2] ~^ image[18][24] + kernel[2][3] ~^ image[18][25] + kernel[2][4] ~^ image[18][26] + kernel[3][0] ~^ image[19][22] + kernel[3][1] ~^ image[19][23] + kernel[3][2] ~^ image[19][24] + kernel[3][3] ~^ image[19][25] + kernel[3][4] ~^ image[19][26] + kernel[4][0] ~^ image[20][22] + kernel[4][1] ~^ image[20][23] + kernel[4][2] ~^ image[20][24] + kernel[4][3] ~^ image[20][25] + kernel[4][4] ~^ image[20][26];
assign xor_sum[16][23] = kernel[0][0] ~^ image[16][23] + kernel[0][1] ~^ image[16][24] + kernel[0][2] ~^ image[16][25] + kernel[0][3] ~^ image[16][26] + kernel[0][4] ~^ image[16][27] + kernel[1][0] ~^ image[17][23] + kernel[1][1] ~^ image[17][24] + kernel[1][2] ~^ image[17][25] + kernel[1][3] ~^ image[17][26] + kernel[1][4] ~^ image[17][27] + kernel[2][0] ~^ image[18][23] + kernel[2][1] ~^ image[18][24] + kernel[2][2] ~^ image[18][25] + kernel[2][3] ~^ image[18][26] + kernel[2][4] ~^ image[18][27] + kernel[3][0] ~^ image[19][23] + kernel[3][1] ~^ image[19][24] + kernel[3][2] ~^ image[19][25] + kernel[3][3] ~^ image[19][26] + kernel[3][4] ~^ image[19][27] + kernel[4][0] ~^ image[20][23] + kernel[4][1] ~^ image[20][24] + kernel[4][2] ~^ image[20][25] + kernel[4][3] ~^ image[20][26] + kernel[4][4] ~^ image[20][27];
assign xor_sum[17][0] = kernel[0][0] ~^ image[17][0] + kernel[0][1] ~^ image[17][1] + kernel[0][2] ~^ image[17][2] + kernel[0][3] ~^ image[17][3] + kernel[0][4] ~^ image[17][4] + kernel[1][0] ~^ image[18][0] + kernel[1][1] ~^ image[18][1] + kernel[1][2] ~^ image[18][2] + kernel[1][3] ~^ image[18][3] + kernel[1][4] ~^ image[18][4] + kernel[2][0] ~^ image[19][0] + kernel[2][1] ~^ image[19][1] + kernel[2][2] ~^ image[19][2] + kernel[2][3] ~^ image[19][3] + kernel[2][4] ~^ image[19][4] + kernel[3][0] ~^ image[20][0] + kernel[3][1] ~^ image[20][1] + kernel[3][2] ~^ image[20][2] + kernel[3][3] ~^ image[20][3] + kernel[3][4] ~^ image[20][4] + kernel[4][0] ~^ image[21][0] + kernel[4][1] ~^ image[21][1] + kernel[4][2] ~^ image[21][2] + kernel[4][3] ~^ image[21][3] + kernel[4][4] ~^ image[21][4];
assign xor_sum[17][1] = kernel[0][0] ~^ image[17][1] + kernel[0][1] ~^ image[17][2] + kernel[0][2] ~^ image[17][3] + kernel[0][3] ~^ image[17][4] + kernel[0][4] ~^ image[17][5] + kernel[1][0] ~^ image[18][1] + kernel[1][1] ~^ image[18][2] + kernel[1][2] ~^ image[18][3] + kernel[1][3] ~^ image[18][4] + kernel[1][4] ~^ image[18][5] + kernel[2][0] ~^ image[19][1] + kernel[2][1] ~^ image[19][2] + kernel[2][2] ~^ image[19][3] + kernel[2][3] ~^ image[19][4] + kernel[2][4] ~^ image[19][5] + kernel[3][0] ~^ image[20][1] + kernel[3][1] ~^ image[20][2] + kernel[3][2] ~^ image[20][3] + kernel[3][3] ~^ image[20][4] + kernel[3][4] ~^ image[20][5] + kernel[4][0] ~^ image[21][1] + kernel[4][1] ~^ image[21][2] + kernel[4][2] ~^ image[21][3] + kernel[4][3] ~^ image[21][4] + kernel[4][4] ~^ image[21][5];
assign xor_sum[17][2] = kernel[0][0] ~^ image[17][2] + kernel[0][1] ~^ image[17][3] + kernel[0][2] ~^ image[17][4] + kernel[0][3] ~^ image[17][5] + kernel[0][4] ~^ image[17][6] + kernel[1][0] ~^ image[18][2] + kernel[1][1] ~^ image[18][3] + kernel[1][2] ~^ image[18][4] + kernel[1][3] ~^ image[18][5] + kernel[1][4] ~^ image[18][6] + kernel[2][0] ~^ image[19][2] + kernel[2][1] ~^ image[19][3] + kernel[2][2] ~^ image[19][4] + kernel[2][3] ~^ image[19][5] + kernel[2][4] ~^ image[19][6] + kernel[3][0] ~^ image[20][2] + kernel[3][1] ~^ image[20][3] + kernel[3][2] ~^ image[20][4] + kernel[3][3] ~^ image[20][5] + kernel[3][4] ~^ image[20][6] + kernel[4][0] ~^ image[21][2] + kernel[4][1] ~^ image[21][3] + kernel[4][2] ~^ image[21][4] + kernel[4][3] ~^ image[21][5] + kernel[4][4] ~^ image[21][6];
assign xor_sum[17][3] = kernel[0][0] ~^ image[17][3] + kernel[0][1] ~^ image[17][4] + kernel[0][2] ~^ image[17][5] + kernel[0][3] ~^ image[17][6] + kernel[0][4] ~^ image[17][7] + kernel[1][0] ~^ image[18][3] + kernel[1][1] ~^ image[18][4] + kernel[1][2] ~^ image[18][5] + kernel[1][3] ~^ image[18][6] + kernel[1][4] ~^ image[18][7] + kernel[2][0] ~^ image[19][3] + kernel[2][1] ~^ image[19][4] + kernel[2][2] ~^ image[19][5] + kernel[2][3] ~^ image[19][6] + kernel[2][4] ~^ image[19][7] + kernel[3][0] ~^ image[20][3] + kernel[3][1] ~^ image[20][4] + kernel[3][2] ~^ image[20][5] + kernel[3][3] ~^ image[20][6] + kernel[3][4] ~^ image[20][7] + kernel[4][0] ~^ image[21][3] + kernel[4][1] ~^ image[21][4] + kernel[4][2] ~^ image[21][5] + kernel[4][3] ~^ image[21][6] + kernel[4][4] ~^ image[21][7];
assign xor_sum[17][4] = kernel[0][0] ~^ image[17][4] + kernel[0][1] ~^ image[17][5] + kernel[0][2] ~^ image[17][6] + kernel[0][3] ~^ image[17][7] + kernel[0][4] ~^ image[17][8] + kernel[1][0] ~^ image[18][4] + kernel[1][1] ~^ image[18][5] + kernel[1][2] ~^ image[18][6] + kernel[1][3] ~^ image[18][7] + kernel[1][4] ~^ image[18][8] + kernel[2][0] ~^ image[19][4] + kernel[2][1] ~^ image[19][5] + kernel[2][2] ~^ image[19][6] + kernel[2][3] ~^ image[19][7] + kernel[2][4] ~^ image[19][8] + kernel[3][0] ~^ image[20][4] + kernel[3][1] ~^ image[20][5] + kernel[3][2] ~^ image[20][6] + kernel[3][3] ~^ image[20][7] + kernel[3][4] ~^ image[20][8] + kernel[4][0] ~^ image[21][4] + kernel[4][1] ~^ image[21][5] + kernel[4][2] ~^ image[21][6] + kernel[4][3] ~^ image[21][7] + kernel[4][4] ~^ image[21][8];
assign xor_sum[17][5] = kernel[0][0] ~^ image[17][5] + kernel[0][1] ~^ image[17][6] + kernel[0][2] ~^ image[17][7] + kernel[0][3] ~^ image[17][8] + kernel[0][4] ~^ image[17][9] + kernel[1][0] ~^ image[18][5] + kernel[1][1] ~^ image[18][6] + kernel[1][2] ~^ image[18][7] + kernel[1][3] ~^ image[18][8] + kernel[1][4] ~^ image[18][9] + kernel[2][0] ~^ image[19][5] + kernel[2][1] ~^ image[19][6] + kernel[2][2] ~^ image[19][7] + kernel[2][3] ~^ image[19][8] + kernel[2][4] ~^ image[19][9] + kernel[3][0] ~^ image[20][5] + kernel[3][1] ~^ image[20][6] + kernel[3][2] ~^ image[20][7] + kernel[3][3] ~^ image[20][8] + kernel[3][4] ~^ image[20][9] + kernel[4][0] ~^ image[21][5] + kernel[4][1] ~^ image[21][6] + kernel[4][2] ~^ image[21][7] + kernel[4][3] ~^ image[21][8] + kernel[4][4] ~^ image[21][9];
assign xor_sum[17][6] = kernel[0][0] ~^ image[17][6] + kernel[0][1] ~^ image[17][7] + kernel[0][2] ~^ image[17][8] + kernel[0][3] ~^ image[17][9] + kernel[0][4] ~^ image[17][10] + kernel[1][0] ~^ image[18][6] + kernel[1][1] ~^ image[18][7] + kernel[1][2] ~^ image[18][8] + kernel[1][3] ~^ image[18][9] + kernel[1][4] ~^ image[18][10] + kernel[2][0] ~^ image[19][6] + kernel[2][1] ~^ image[19][7] + kernel[2][2] ~^ image[19][8] + kernel[2][3] ~^ image[19][9] + kernel[2][4] ~^ image[19][10] + kernel[3][0] ~^ image[20][6] + kernel[3][1] ~^ image[20][7] + kernel[3][2] ~^ image[20][8] + kernel[3][3] ~^ image[20][9] + kernel[3][4] ~^ image[20][10] + kernel[4][0] ~^ image[21][6] + kernel[4][1] ~^ image[21][7] + kernel[4][2] ~^ image[21][8] + kernel[4][3] ~^ image[21][9] + kernel[4][4] ~^ image[21][10];
assign xor_sum[17][7] = kernel[0][0] ~^ image[17][7] + kernel[0][1] ~^ image[17][8] + kernel[0][2] ~^ image[17][9] + kernel[0][3] ~^ image[17][10] + kernel[0][4] ~^ image[17][11] + kernel[1][0] ~^ image[18][7] + kernel[1][1] ~^ image[18][8] + kernel[1][2] ~^ image[18][9] + kernel[1][3] ~^ image[18][10] + kernel[1][4] ~^ image[18][11] + kernel[2][0] ~^ image[19][7] + kernel[2][1] ~^ image[19][8] + kernel[2][2] ~^ image[19][9] + kernel[2][3] ~^ image[19][10] + kernel[2][4] ~^ image[19][11] + kernel[3][0] ~^ image[20][7] + kernel[3][1] ~^ image[20][8] + kernel[3][2] ~^ image[20][9] + kernel[3][3] ~^ image[20][10] + kernel[3][4] ~^ image[20][11] + kernel[4][0] ~^ image[21][7] + kernel[4][1] ~^ image[21][8] + kernel[4][2] ~^ image[21][9] + kernel[4][3] ~^ image[21][10] + kernel[4][4] ~^ image[21][11];
assign xor_sum[17][8] = kernel[0][0] ~^ image[17][8] + kernel[0][1] ~^ image[17][9] + kernel[0][2] ~^ image[17][10] + kernel[0][3] ~^ image[17][11] + kernel[0][4] ~^ image[17][12] + kernel[1][0] ~^ image[18][8] + kernel[1][1] ~^ image[18][9] + kernel[1][2] ~^ image[18][10] + kernel[1][3] ~^ image[18][11] + kernel[1][4] ~^ image[18][12] + kernel[2][0] ~^ image[19][8] + kernel[2][1] ~^ image[19][9] + kernel[2][2] ~^ image[19][10] + kernel[2][3] ~^ image[19][11] + kernel[2][4] ~^ image[19][12] + kernel[3][0] ~^ image[20][8] + kernel[3][1] ~^ image[20][9] + kernel[3][2] ~^ image[20][10] + kernel[3][3] ~^ image[20][11] + kernel[3][4] ~^ image[20][12] + kernel[4][0] ~^ image[21][8] + kernel[4][1] ~^ image[21][9] + kernel[4][2] ~^ image[21][10] + kernel[4][3] ~^ image[21][11] + kernel[4][4] ~^ image[21][12];
assign xor_sum[17][9] = kernel[0][0] ~^ image[17][9] + kernel[0][1] ~^ image[17][10] + kernel[0][2] ~^ image[17][11] + kernel[0][3] ~^ image[17][12] + kernel[0][4] ~^ image[17][13] + kernel[1][0] ~^ image[18][9] + kernel[1][1] ~^ image[18][10] + kernel[1][2] ~^ image[18][11] + kernel[1][3] ~^ image[18][12] + kernel[1][4] ~^ image[18][13] + kernel[2][0] ~^ image[19][9] + kernel[2][1] ~^ image[19][10] + kernel[2][2] ~^ image[19][11] + kernel[2][3] ~^ image[19][12] + kernel[2][4] ~^ image[19][13] + kernel[3][0] ~^ image[20][9] + kernel[3][1] ~^ image[20][10] + kernel[3][2] ~^ image[20][11] + kernel[3][3] ~^ image[20][12] + kernel[3][4] ~^ image[20][13] + kernel[4][0] ~^ image[21][9] + kernel[4][1] ~^ image[21][10] + kernel[4][2] ~^ image[21][11] + kernel[4][3] ~^ image[21][12] + kernel[4][4] ~^ image[21][13];
assign xor_sum[17][10] = kernel[0][0] ~^ image[17][10] + kernel[0][1] ~^ image[17][11] + kernel[0][2] ~^ image[17][12] + kernel[0][3] ~^ image[17][13] + kernel[0][4] ~^ image[17][14] + kernel[1][0] ~^ image[18][10] + kernel[1][1] ~^ image[18][11] + kernel[1][2] ~^ image[18][12] + kernel[1][3] ~^ image[18][13] + kernel[1][4] ~^ image[18][14] + kernel[2][0] ~^ image[19][10] + kernel[2][1] ~^ image[19][11] + kernel[2][2] ~^ image[19][12] + kernel[2][3] ~^ image[19][13] + kernel[2][4] ~^ image[19][14] + kernel[3][0] ~^ image[20][10] + kernel[3][1] ~^ image[20][11] + kernel[3][2] ~^ image[20][12] + kernel[3][3] ~^ image[20][13] + kernel[3][4] ~^ image[20][14] + kernel[4][0] ~^ image[21][10] + kernel[4][1] ~^ image[21][11] + kernel[4][2] ~^ image[21][12] + kernel[4][3] ~^ image[21][13] + kernel[4][4] ~^ image[21][14];
assign xor_sum[17][11] = kernel[0][0] ~^ image[17][11] + kernel[0][1] ~^ image[17][12] + kernel[0][2] ~^ image[17][13] + kernel[0][3] ~^ image[17][14] + kernel[0][4] ~^ image[17][15] + kernel[1][0] ~^ image[18][11] + kernel[1][1] ~^ image[18][12] + kernel[1][2] ~^ image[18][13] + kernel[1][3] ~^ image[18][14] + kernel[1][4] ~^ image[18][15] + kernel[2][0] ~^ image[19][11] + kernel[2][1] ~^ image[19][12] + kernel[2][2] ~^ image[19][13] + kernel[2][3] ~^ image[19][14] + kernel[2][4] ~^ image[19][15] + kernel[3][0] ~^ image[20][11] + kernel[3][1] ~^ image[20][12] + kernel[3][2] ~^ image[20][13] + kernel[3][3] ~^ image[20][14] + kernel[3][4] ~^ image[20][15] + kernel[4][0] ~^ image[21][11] + kernel[4][1] ~^ image[21][12] + kernel[4][2] ~^ image[21][13] + kernel[4][3] ~^ image[21][14] + kernel[4][4] ~^ image[21][15];
assign xor_sum[17][12] = kernel[0][0] ~^ image[17][12] + kernel[0][1] ~^ image[17][13] + kernel[0][2] ~^ image[17][14] + kernel[0][3] ~^ image[17][15] + kernel[0][4] ~^ image[17][16] + kernel[1][0] ~^ image[18][12] + kernel[1][1] ~^ image[18][13] + kernel[1][2] ~^ image[18][14] + kernel[1][3] ~^ image[18][15] + kernel[1][4] ~^ image[18][16] + kernel[2][0] ~^ image[19][12] + kernel[2][1] ~^ image[19][13] + kernel[2][2] ~^ image[19][14] + kernel[2][3] ~^ image[19][15] + kernel[2][4] ~^ image[19][16] + kernel[3][0] ~^ image[20][12] + kernel[3][1] ~^ image[20][13] + kernel[3][2] ~^ image[20][14] + kernel[3][3] ~^ image[20][15] + kernel[3][4] ~^ image[20][16] + kernel[4][0] ~^ image[21][12] + kernel[4][1] ~^ image[21][13] + kernel[4][2] ~^ image[21][14] + kernel[4][3] ~^ image[21][15] + kernel[4][4] ~^ image[21][16];
assign xor_sum[17][13] = kernel[0][0] ~^ image[17][13] + kernel[0][1] ~^ image[17][14] + kernel[0][2] ~^ image[17][15] + kernel[0][3] ~^ image[17][16] + kernel[0][4] ~^ image[17][17] + kernel[1][0] ~^ image[18][13] + kernel[1][1] ~^ image[18][14] + kernel[1][2] ~^ image[18][15] + kernel[1][3] ~^ image[18][16] + kernel[1][4] ~^ image[18][17] + kernel[2][0] ~^ image[19][13] + kernel[2][1] ~^ image[19][14] + kernel[2][2] ~^ image[19][15] + kernel[2][3] ~^ image[19][16] + kernel[2][4] ~^ image[19][17] + kernel[3][0] ~^ image[20][13] + kernel[3][1] ~^ image[20][14] + kernel[3][2] ~^ image[20][15] + kernel[3][3] ~^ image[20][16] + kernel[3][4] ~^ image[20][17] + kernel[4][0] ~^ image[21][13] + kernel[4][1] ~^ image[21][14] + kernel[4][2] ~^ image[21][15] + kernel[4][3] ~^ image[21][16] + kernel[4][4] ~^ image[21][17];
assign xor_sum[17][14] = kernel[0][0] ~^ image[17][14] + kernel[0][1] ~^ image[17][15] + kernel[0][2] ~^ image[17][16] + kernel[0][3] ~^ image[17][17] + kernel[0][4] ~^ image[17][18] + kernel[1][0] ~^ image[18][14] + kernel[1][1] ~^ image[18][15] + kernel[1][2] ~^ image[18][16] + kernel[1][3] ~^ image[18][17] + kernel[1][4] ~^ image[18][18] + kernel[2][0] ~^ image[19][14] + kernel[2][1] ~^ image[19][15] + kernel[2][2] ~^ image[19][16] + kernel[2][3] ~^ image[19][17] + kernel[2][4] ~^ image[19][18] + kernel[3][0] ~^ image[20][14] + kernel[3][1] ~^ image[20][15] + kernel[3][2] ~^ image[20][16] + kernel[3][3] ~^ image[20][17] + kernel[3][4] ~^ image[20][18] + kernel[4][0] ~^ image[21][14] + kernel[4][1] ~^ image[21][15] + kernel[4][2] ~^ image[21][16] + kernel[4][3] ~^ image[21][17] + kernel[4][4] ~^ image[21][18];
assign xor_sum[17][15] = kernel[0][0] ~^ image[17][15] + kernel[0][1] ~^ image[17][16] + kernel[0][2] ~^ image[17][17] + kernel[0][3] ~^ image[17][18] + kernel[0][4] ~^ image[17][19] + kernel[1][0] ~^ image[18][15] + kernel[1][1] ~^ image[18][16] + kernel[1][2] ~^ image[18][17] + kernel[1][3] ~^ image[18][18] + kernel[1][4] ~^ image[18][19] + kernel[2][0] ~^ image[19][15] + kernel[2][1] ~^ image[19][16] + kernel[2][2] ~^ image[19][17] + kernel[2][3] ~^ image[19][18] + kernel[2][4] ~^ image[19][19] + kernel[3][0] ~^ image[20][15] + kernel[3][1] ~^ image[20][16] + kernel[3][2] ~^ image[20][17] + kernel[3][3] ~^ image[20][18] + kernel[3][4] ~^ image[20][19] + kernel[4][0] ~^ image[21][15] + kernel[4][1] ~^ image[21][16] + kernel[4][2] ~^ image[21][17] + kernel[4][3] ~^ image[21][18] + kernel[4][4] ~^ image[21][19];
assign xor_sum[17][16] = kernel[0][0] ~^ image[17][16] + kernel[0][1] ~^ image[17][17] + kernel[0][2] ~^ image[17][18] + kernel[0][3] ~^ image[17][19] + kernel[0][4] ~^ image[17][20] + kernel[1][0] ~^ image[18][16] + kernel[1][1] ~^ image[18][17] + kernel[1][2] ~^ image[18][18] + kernel[1][3] ~^ image[18][19] + kernel[1][4] ~^ image[18][20] + kernel[2][0] ~^ image[19][16] + kernel[2][1] ~^ image[19][17] + kernel[2][2] ~^ image[19][18] + kernel[2][3] ~^ image[19][19] + kernel[2][4] ~^ image[19][20] + kernel[3][0] ~^ image[20][16] + kernel[3][1] ~^ image[20][17] + kernel[3][2] ~^ image[20][18] + kernel[3][3] ~^ image[20][19] + kernel[3][4] ~^ image[20][20] + kernel[4][0] ~^ image[21][16] + kernel[4][1] ~^ image[21][17] + kernel[4][2] ~^ image[21][18] + kernel[4][3] ~^ image[21][19] + kernel[4][4] ~^ image[21][20];
assign xor_sum[17][17] = kernel[0][0] ~^ image[17][17] + kernel[0][1] ~^ image[17][18] + kernel[0][2] ~^ image[17][19] + kernel[0][3] ~^ image[17][20] + kernel[0][4] ~^ image[17][21] + kernel[1][0] ~^ image[18][17] + kernel[1][1] ~^ image[18][18] + kernel[1][2] ~^ image[18][19] + kernel[1][3] ~^ image[18][20] + kernel[1][4] ~^ image[18][21] + kernel[2][0] ~^ image[19][17] + kernel[2][1] ~^ image[19][18] + kernel[2][2] ~^ image[19][19] + kernel[2][3] ~^ image[19][20] + kernel[2][4] ~^ image[19][21] + kernel[3][0] ~^ image[20][17] + kernel[3][1] ~^ image[20][18] + kernel[3][2] ~^ image[20][19] + kernel[3][3] ~^ image[20][20] + kernel[3][4] ~^ image[20][21] + kernel[4][0] ~^ image[21][17] + kernel[4][1] ~^ image[21][18] + kernel[4][2] ~^ image[21][19] + kernel[4][3] ~^ image[21][20] + kernel[4][4] ~^ image[21][21];
assign xor_sum[17][18] = kernel[0][0] ~^ image[17][18] + kernel[0][1] ~^ image[17][19] + kernel[0][2] ~^ image[17][20] + kernel[0][3] ~^ image[17][21] + kernel[0][4] ~^ image[17][22] + kernel[1][0] ~^ image[18][18] + kernel[1][1] ~^ image[18][19] + kernel[1][2] ~^ image[18][20] + kernel[1][3] ~^ image[18][21] + kernel[1][4] ~^ image[18][22] + kernel[2][0] ~^ image[19][18] + kernel[2][1] ~^ image[19][19] + kernel[2][2] ~^ image[19][20] + kernel[2][3] ~^ image[19][21] + kernel[2][4] ~^ image[19][22] + kernel[3][0] ~^ image[20][18] + kernel[3][1] ~^ image[20][19] + kernel[3][2] ~^ image[20][20] + kernel[3][3] ~^ image[20][21] + kernel[3][4] ~^ image[20][22] + kernel[4][0] ~^ image[21][18] + kernel[4][1] ~^ image[21][19] + kernel[4][2] ~^ image[21][20] + kernel[4][3] ~^ image[21][21] + kernel[4][4] ~^ image[21][22];
assign xor_sum[17][19] = kernel[0][0] ~^ image[17][19] + kernel[0][1] ~^ image[17][20] + kernel[0][2] ~^ image[17][21] + kernel[0][3] ~^ image[17][22] + kernel[0][4] ~^ image[17][23] + kernel[1][0] ~^ image[18][19] + kernel[1][1] ~^ image[18][20] + kernel[1][2] ~^ image[18][21] + kernel[1][3] ~^ image[18][22] + kernel[1][4] ~^ image[18][23] + kernel[2][0] ~^ image[19][19] + kernel[2][1] ~^ image[19][20] + kernel[2][2] ~^ image[19][21] + kernel[2][3] ~^ image[19][22] + kernel[2][4] ~^ image[19][23] + kernel[3][0] ~^ image[20][19] + kernel[3][1] ~^ image[20][20] + kernel[3][2] ~^ image[20][21] + kernel[3][3] ~^ image[20][22] + kernel[3][4] ~^ image[20][23] + kernel[4][0] ~^ image[21][19] + kernel[4][1] ~^ image[21][20] + kernel[4][2] ~^ image[21][21] + kernel[4][3] ~^ image[21][22] + kernel[4][4] ~^ image[21][23];
assign xor_sum[17][20] = kernel[0][0] ~^ image[17][20] + kernel[0][1] ~^ image[17][21] + kernel[0][2] ~^ image[17][22] + kernel[0][3] ~^ image[17][23] + kernel[0][4] ~^ image[17][24] + kernel[1][0] ~^ image[18][20] + kernel[1][1] ~^ image[18][21] + kernel[1][2] ~^ image[18][22] + kernel[1][3] ~^ image[18][23] + kernel[1][4] ~^ image[18][24] + kernel[2][0] ~^ image[19][20] + kernel[2][1] ~^ image[19][21] + kernel[2][2] ~^ image[19][22] + kernel[2][3] ~^ image[19][23] + kernel[2][4] ~^ image[19][24] + kernel[3][0] ~^ image[20][20] + kernel[3][1] ~^ image[20][21] + kernel[3][2] ~^ image[20][22] + kernel[3][3] ~^ image[20][23] + kernel[3][4] ~^ image[20][24] + kernel[4][0] ~^ image[21][20] + kernel[4][1] ~^ image[21][21] + kernel[4][2] ~^ image[21][22] + kernel[4][3] ~^ image[21][23] + kernel[4][4] ~^ image[21][24];
assign xor_sum[17][21] = kernel[0][0] ~^ image[17][21] + kernel[0][1] ~^ image[17][22] + kernel[0][2] ~^ image[17][23] + kernel[0][3] ~^ image[17][24] + kernel[0][4] ~^ image[17][25] + kernel[1][0] ~^ image[18][21] + kernel[1][1] ~^ image[18][22] + kernel[1][2] ~^ image[18][23] + kernel[1][3] ~^ image[18][24] + kernel[1][4] ~^ image[18][25] + kernel[2][0] ~^ image[19][21] + kernel[2][1] ~^ image[19][22] + kernel[2][2] ~^ image[19][23] + kernel[2][3] ~^ image[19][24] + kernel[2][4] ~^ image[19][25] + kernel[3][0] ~^ image[20][21] + kernel[3][1] ~^ image[20][22] + kernel[3][2] ~^ image[20][23] + kernel[3][3] ~^ image[20][24] + kernel[3][4] ~^ image[20][25] + kernel[4][0] ~^ image[21][21] + kernel[4][1] ~^ image[21][22] + kernel[4][2] ~^ image[21][23] + kernel[4][3] ~^ image[21][24] + kernel[4][4] ~^ image[21][25];
assign xor_sum[17][22] = kernel[0][0] ~^ image[17][22] + kernel[0][1] ~^ image[17][23] + kernel[0][2] ~^ image[17][24] + kernel[0][3] ~^ image[17][25] + kernel[0][4] ~^ image[17][26] + kernel[1][0] ~^ image[18][22] + kernel[1][1] ~^ image[18][23] + kernel[1][2] ~^ image[18][24] + kernel[1][3] ~^ image[18][25] + kernel[1][4] ~^ image[18][26] + kernel[2][0] ~^ image[19][22] + kernel[2][1] ~^ image[19][23] + kernel[2][2] ~^ image[19][24] + kernel[2][3] ~^ image[19][25] + kernel[2][4] ~^ image[19][26] + kernel[3][0] ~^ image[20][22] + kernel[3][1] ~^ image[20][23] + kernel[3][2] ~^ image[20][24] + kernel[3][3] ~^ image[20][25] + kernel[3][4] ~^ image[20][26] + kernel[4][0] ~^ image[21][22] + kernel[4][1] ~^ image[21][23] + kernel[4][2] ~^ image[21][24] + kernel[4][3] ~^ image[21][25] + kernel[4][4] ~^ image[21][26];
assign xor_sum[17][23] = kernel[0][0] ~^ image[17][23] + kernel[0][1] ~^ image[17][24] + kernel[0][2] ~^ image[17][25] + kernel[0][3] ~^ image[17][26] + kernel[0][4] ~^ image[17][27] + kernel[1][0] ~^ image[18][23] + kernel[1][1] ~^ image[18][24] + kernel[1][2] ~^ image[18][25] + kernel[1][3] ~^ image[18][26] + kernel[1][4] ~^ image[18][27] + kernel[2][0] ~^ image[19][23] + kernel[2][1] ~^ image[19][24] + kernel[2][2] ~^ image[19][25] + kernel[2][3] ~^ image[19][26] + kernel[2][4] ~^ image[19][27] + kernel[3][0] ~^ image[20][23] + kernel[3][1] ~^ image[20][24] + kernel[3][2] ~^ image[20][25] + kernel[3][3] ~^ image[20][26] + kernel[3][4] ~^ image[20][27] + kernel[4][0] ~^ image[21][23] + kernel[4][1] ~^ image[21][24] + kernel[4][2] ~^ image[21][25] + kernel[4][3] ~^ image[21][26] + kernel[4][4] ~^ image[21][27];
assign xor_sum[18][0] = kernel[0][0] ~^ image[18][0] + kernel[0][1] ~^ image[18][1] + kernel[0][2] ~^ image[18][2] + kernel[0][3] ~^ image[18][3] + kernel[0][4] ~^ image[18][4] + kernel[1][0] ~^ image[19][0] + kernel[1][1] ~^ image[19][1] + kernel[1][2] ~^ image[19][2] + kernel[1][3] ~^ image[19][3] + kernel[1][4] ~^ image[19][4] + kernel[2][0] ~^ image[20][0] + kernel[2][1] ~^ image[20][1] + kernel[2][2] ~^ image[20][2] + kernel[2][3] ~^ image[20][3] + kernel[2][4] ~^ image[20][4] + kernel[3][0] ~^ image[21][0] + kernel[3][1] ~^ image[21][1] + kernel[3][2] ~^ image[21][2] + kernel[3][3] ~^ image[21][3] + kernel[3][4] ~^ image[21][4] + kernel[4][0] ~^ image[22][0] + kernel[4][1] ~^ image[22][1] + kernel[4][2] ~^ image[22][2] + kernel[4][3] ~^ image[22][3] + kernel[4][4] ~^ image[22][4];
assign xor_sum[18][1] = kernel[0][0] ~^ image[18][1] + kernel[0][1] ~^ image[18][2] + kernel[0][2] ~^ image[18][3] + kernel[0][3] ~^ image[18][4] + kernel[0][4] ~^ image[18][5] + kernel[1][0] ~^ image[19][1] + kernel[1][1] ~^ image[19][2] + kernel[1][2] ~^ image[19][3] + kernel[1][3] ~^ image[19][4] + kernel[1][4] ~^ image[19][5] + kernel[2][0] ~^ image[20][1] + kernel[2][1] ~^ image[20][2] + kernel[2][2] ~^ image[20][3] + kernel[2][3] ~^ image[20][4] + kernel[2][4] ~^ image[20][5] + kernel[3][0] ~^ image[21][1] + kernel[3][1] ~^ image[21][2] + kernel[3][2] ~^ image[21][3] + kernel[3][3] ~^ image[21][4] + kernel[3][4] ~^ image[21][5] + kernel[4][0] ~^ image[22][1] + kernel[4][1] ~^ image[22][2] + kernel[4][2] ~^ image[22][3] + kernel[4][3] ~^ image[22][4] + kernel[4][4] ~^ image[22][5];
assign xor_sum[18][2] = kernel[0][0] ~^ image[18][2] + kernel[0][1] ~^ image[18][3] + kernel[0][2] ~^ image[18][4] + kernel[0][3] ~^ image[18][5] + kernel[0][4] ~^ image[18][6] + kernel[1][0] ~^ image[19][2] + kernel[1][1] ~^ image[19][3] + kernel[1][2] ~^ image[19][4] + kernel[1][3] ~^ image[19][5] + kernel[1][4] ~^ image[19][6] + kernel[2][0] ~^ image[20][2] + kernel[2][1] ~^ image[20][3] + kernel[2][2] ~^ image[20][4] + kernel[2][3] ~^ image[20][5] + kernel[2][4] ~^ image[20][6] + kernel[3][0] ~^ image[21][2] + kernel[3][1] ~^ image[21][3] + kernel[3][2] ~^ image[21][4] + kernel[3][3] ~^ image[21][5] + kernel[3][4] ~^ image[21][6] + kernel[4][0] ~^ image[22][2] + kernel[4][1] ~^ image[22][3] + kernel[4][2] ~^ image[22][4] + kernel[4][3] ~^ image[22][5] + kernel[4][4] ~^ image[22][6];
assign xor_sum[18][3] = kernel[0][0] ~^ image[18][3] + kernel[0][1] ~^ image[18][4] + kernel[0][2] ~^ image[18][5] + kernel[0][3] ~^ image[18][6] + kernel[0][4] ~^ image[18][7] + kernel[1][0] ~^ image[19][3] + kernel[1][1] ~^ image[19][4] + kernel[1][2] ~^ image[19][5] + kernel[1][3] ~^ image[19][6] + kernel[1][4] ~^ image[19][7] + kernel[2][0] ~^ image[20][3] + kernel[2][1] ~^ image[20][4] + kernel[2][2] ~^ image[20][5] + kernel[2][3] ~^ image[20][6] + kernel[2][4] ~^ image[20][7] + kernel[3][0] ~^ image[21][3] + kernel[3][1] ~^ image[21][4] + kernel[3][2] ~^ image[21][5] + kernel[3][3] ~^ image[21][6] + kernel[3][4] ~^ image[21][7] + kernel[4][0] ~^ image[22][3] + kernel[4][1] ~^ image[22][4] + kernel[4][2] ~^ image[22][5] + kernel[4][3] ~^ image[22][6] + kernel[4][4] ~^ image[22][7];
assign xor_sum[18][4] = kernel[0][0] ~^ image[18][4] + kernel[0][1] ~^ image[18][5] + kernel[0][2] ~^ image[18][6] + kernel[0][3] ~^ image[18][7] + kernel[0][4] ~^ image[18][8] + kernel[1][0] ~^ image[19][4] + kernel[1][1] ~^ image[19][5] + kernel[1][2] ~^ image[19][6] + kernel[1][3] ~^ image[19][7] + kernel[1][4] ~^ image[19][8] + kernel[2][0] ~^ image[20][4] + kernel[2][1] ~^ image[20][5] + kernel[2][2] ~^ image[20][6] + kernel[2][3] ~^ image[20][7] + kernel[2][4] ~^ image[20][8] + kernel[3][0] ~^ image[21][4] + kernel[3][1] ~^ image[21][5] + kernel[3][2] ~^ image[21][6] + kernel[3][3] ~^ image[21][7] + kernel[3][4] ~^ image[21][8] + kernel[4][0] ~^ image[22][4] + kernel[4][1] ~^ image[22][5] + kernel[4][2] ~^ image[22][6] + kernel[4][3] ~^ image[22][7] + kernel[4][4] ~^ image[22][8];
assign xor_sum[18][5] = kernel[0][0] ~^ image[18][5] + kernel[0][1] ~^ image[18][6] + kernel[0][2] ~^ image[18][7] + kernel[0][3] ~^ image[18][8] + kernel[0][4] ~^ image[18][9] + kernel[1][0] ~^ image[19][5] + kernel[1][1] ~^ image[19][6] + kernel[1][2] ~^ image[19][7] + kernel[1][3] ~^ image[19][8] + kernel[1][4] ~^ image[19][9] + kernel[2][0] ~^ image[20][5] + kernel[2][1] ~^ image[20][6] + kernel[2][2] ~^ image[20][7] + kernel[2][3] ~^ image[20][8] + kernel[2][4] ~^ image[20][9] + kernel[3][0] ~^ image[21][5] + kernel[3][1] ~^ image[21][6] + kernel[3][2] ~^ image[21][7] + kernel[3][3] ~^ image[21][8] + kernel[3][4] ~^ image[21][9] + kernel[4][0] ~^ image[22][5] + kernel[4][1] ~^ image[22][6] + kernel[4][2] ~^ image[22][7] + kernel[4][3] ~^ image[22][8] + kernel[4][4] ~^ image[22][9];
assign xor_sum[18][6] = kernel[0][0] ~^ image[18][6] + kernel[0][1] ~^ image[18][7] + kernel[0][2] ~^ image[18][8] + kernel[0][3] ~^ image[18][9] + kernel[0][4] ~^ image[18][10] + kernel[1][0] ~^ image[19][6] + kernel[1][1] ~^ image[19][7] + kernel[1][2] ~^ image[19][8] + kernel[1][3] ~^ image[19][9] + kernel[1][4] ~^ image[19][10] + kernel[2][0] ~^ image[20][6] + kernel[2][1] ~^ image[20][7] + kernel[2][2] ~^ image[20][8] + kernel[2][3] ~^ image[20][9] + kernel[2][4] ~^ image[20][10] + kernel[3][0] ~^ image[21][6] + kernel[3][1] ~^ image[21][7] + kernel[3][2] ~^ image[21][8] + kernel[3][3] ~^ image[21][9] + kernel[3][4] ~^ image[21][10] + kernel[4][0] ~^ image[22][6] + kernel[4][1] ~^ image[22][7] + kernel[4][2] ~^ image[22][8] + kernel[4][3] ~^ image[22][9] + kernel[4][4] ~^ image[22][10];
assign xor_sum[18][7] = kernel[0][0] ~^ image[18][7] + kernel[0][1] ~^ image[18][8] + kernel[0][2] ~^ image[18][9] + kernel[0][3] ~^ image[18][10] + kernel[0][4] ~^ image[18][11] + kernel[1][0] ~^ image[19][7] + kernel[1][1] ~^ image[19][8] + kernel[1][2] ~^ image[19][9] + kernel[1][3] ~^ image[19][10] + kernel[1][4] ~^ image[19][11] + kernel[2][0] ~^ image[20][7] + kernel[2][1] ~^ image[20][8] + kernel[2][2] ~^ image[20][9] + kernel[2][3] ~^ image[20][10] + kernel[2][4] ~^ image[20][11] + kernel[3][0] ~^ image[21][7] + kernel[3][1] ~^ image[21][8] + kernel[3][2] ~^ image[21][9] + kernel[3][3] ~^ image[21][10] + kernel[3][4] ~^ image[21][11] + kernel[4][0] ~^ image[22][7] + kernel[4][1] ~^ image[22][8] + kernel[4][2] ~^ image[22][9] + kernel[4][3] ~^ image[22][10] + kernel[4][4] ~^ image[22][11];
assign xor_sum[18][8] = kernel[0][0] ~^ image[18][8] + kernel[0][1] ~^ image[18][9] + kernel[0][2] ~^ image[18][10] + kernel[0][3] ~^ image[18][11] + kernel[0][4] ~^ image[18][12] + kernel[1][0] ~^ image[19][8] + kernel[1][1] ~^ image[19][9] + kernel[1][2] ~^ image[19][10] + kernel[1][3] ~^ image[19][11] + kernel[1][4] ~^ image[19][12] + kernel[2][0] ~^ image[20][8] + kernel[2][1] ~^ image[20][9] + kernel[2][2] ~^ image[20][10] + kernel[2][3] ~^ image[20][11] + kernel[2][4] ~^ image[20][12] + kernel[3][0] ~^ image[21][8] + kernel[3][1] ~^ image[21][9] + kernel[3][2] ~^ image[21][10] + kernel[3][3] ~^ image[21][11] + kernel[3][4] ~^ image[21][12] + kernel[4][0] ~^ image[22][8] + kernel[4][1] ~^ image[22][9] + kernel[4][2] ~^ image[22][10] + kernel[4][3] ~^ image[22][11] + kernel[4][4] ~^ image[22][12];
assign xor_sum[18][9] = kernel[0][0] ~^ image[18][9] + kernel[0][1] ~^ image[18][10] + kernel[0][2] ~^ image[18][11] + kernel[0][3] ~^ image[18][12] + kernel[0][4] ~^ image[18][13] + kernel[1][0] ~^ image[19][9] + kernel[1][1] ~^ image[19][10] + kernel[1][2] ~^ image[19][11] + kernel[1][3] ~^ image[19][12] + kernel[1][4] ~^ image[19][13] + kernel[2][0] ~^ image[20][9] + kernel[2][1] ~^ image[20][10] + kernel[2][2] ~^ image[20][11] + kernel[2][3] ~^ image[20][12] + kernel[2][4] ~^ image[20][13] + kernel[3][0] ~^ image[21][9] + kernel[3][1] ~^ image[21][10] + kernel[3][2] ~^ image[21][11] + kernel[3][3] ~^ image[21][12] + kernel[3][4] ~^ image[21][13] + kernel[4][0] ~^ image[22][9] + kernel[4][1] ~^ image[22][10] + kernel[4][2] ~^ image[22][11] + kernel[4][3] ~^ image[22][12] + kernel[4][4] ~^ image[22][13];
assign xor_sum[18][10] = kernel[0][0] ~^ image[18][10] + kernel[0][1] ~^ image[18][11] + kernel[0][2] ~^ image[18][12] + kernel[0][3] ~^ image[18][13] + kernel[0][4] ~^ image[18][14] + kernel[1][0] ~^ image[19][10] + kernel[1][1] ~^ image[19][11] + kernel[1][2] ~^ image[19][12] + kernel[1][3] ~^ image[19][13] + kernel[1][4] ~^ image[19][14] + kernel[2][0] ~^ image[20][10] + kernel[2][1] ~^ image[20][11] + kernel[2][2] ~^ image[20][12] + kernel[2][3] ~^ image[20][13] + kernel[2][4] ~^ image[20][14] + kernel[3][0] ~^ image[21][10] + kernel[3][1] ~^ image[21][11] + kernel[3][2] ~^ image[21][12] + kernel[3][3] ~^ image[21][13] + kernel[3][4] ~^ image[21][14] + kernel[4][0] ~^ image[22][10] + kernel[4][1] ~^ image[22][11] + kernel[4][2] ~^ image[22][12] + kernel[4][3] ~^ image[22][13] + kernel[4][4] ~^ image[22][14];
assign xor_sum[18][11] = kernel[0][0] ~^ image[18][11] + kernel[0][1] ~^ image[18][12] + kernel[0][2] ~^ image[18][13] + kernel[0][3] ~^ image[18][14] + kernel[0][4] ~^ image[18][15] + kernel[1][0] ~^ image[19][11] + kernel[1][1] ~^ image[19][12] + kernel[1][2] ~^ image[19][13] + kernel[1][3] ~^ image[19][14] + kernel[1][4] ~^ image[19][15] + kernel[2][0] ~^ image[20][11] + kernel[2][1] ~^ image[20][12] + kernel[2][2] ~^ image[20][13] + kernel[2][3] ~^ image[20][14] + kernel[2][4] ~^ image[20][15] + kernel[3][0] ~^ image[21][11] + kernel[3][1] ~^ image[21][12] + kernel[3][2] ~^ image[21][13] + kernel[3][3] ~^ image[21][14] + kernel[3][4] ~^ image[21][15] + kernel[4][0] ~^ image[22][11] + kernel[4][1] ~^ image[22][12] + kernel[4][2] ~^ image[22][13] + kernel[4][3] ~^ image[22][14] + kernel[4][4] ~^ image[22][15];
assign xor_sum[18][12] = kernel[0][0] ~^ image[18][12] + kernel[0][1] ~^ image[18][13] + kernel[0][2] ~^ image[18][14] + kernel[0][3] ~^ image[18][15] + kernel[0][4] ~^ image[18][16] + kernel[1][0] ~^ image[19][12] + kernel[1][1] ~^ image[19][13] + kernel[1][2] ~^ image[19][14] + kernel[1][3] ~^ image[19][15] + kernel[1][4] ~^ image[19][16] + kernel[2][0] ~^ image[20][12] + kernel[2][1] ~^ image[20][13] + kernel[2][2] ~^ image[20][14] + kernel[2][3] ~^ image[20][15] + kernel[2][4] ~^ image[20][16] + kernel[3][0] ~^ image[21][12] + kernel[3][1] ~^ image[21][13] + kernel[3][2] ~^ image[21][14] + kernel[3][3] ~^ image[21][15] + kernel[3][4] ~^ image[21][16] + kernel[4][0] ~^ image[22][12] + kernel[4][1] ~^ image[22][13] + kernel[4][2] ~^ image[22][14] + kernel[4][3] ~^ image[22][15] + kernel[4][4] ~^ image[22][16];
assign xor_sum[18][13] = kernel[0][0] ~^ image[18][13] + kernel[0][1] ~^ image[18][14] + kernel[0][2] ~^ image[18][15] + kernel[0][3] ~^ image[18][16] + kernel[0][4] ~^ image[18][17] + kernel[1][0] ~^ image[19][13] + kernel[1][1] ~^ image[19][14] + kernel[1][2] ~^ image[19][15] + kernel[1][3] ~^ image[19][16] + kernel[1][4] ~^ image[19][17] + kernel[2][0] ~^ image[20][13] + kernel[2][1] ~^ image[20][14] + kernel[2][2] ~^ image[20][15] + kernel[2][3] ~^ image[20][16] + kernel[2][4] ~^ image[20][17] + kernel[3][0] ~^ image[21][13] + kernel[3][1] ~^ image[21][14] + kernel[3][2] ~^ image[21][15] + kernel[3][3] ~^ image[21][16] + kernel[3][4] ~^ image[21][17] + kernel[4][0] ~^ image[22][13] + kernel[4][1] ~^ image[22][14] + kernel[4][2] ~^ image[22][15] + kernel[4][3] ~^ image[22][16] + kernel[4][4] ~^ image[22][17];
assign xor_sum[18][14] = kernel[0][0] ~^ image[18][14] + kernel[0][1] ~^ image[18][15] + kernel[0][2] ~^ image[18][16] + kernel[0][3] ~^ image[18][17] + kernel[0][4] ~^ image[18][18] + kernel[1][0] ~^ image[19][14] + kernel[1][1] ~^ image[19][15] + kernel[1][2] ~^ image[19][16] + kernel[1][3] ~^ image[19][17] + kernel[1][4] ~^ image[19][18] + kernel[2][0] ~^ image[20][14] + kernel[2][1] ~^ image[20][15] + kernel[2][2] ~^ image[20][16] + kernel[2][3] ~^ image[20][17] + kernel[2][4] ~^ image[20][18] + kernel[3][0] ~^ image[21][14] + kernel[3][1] ~^ image[21][15] + kernel[3][2] ~^ image[21][16] + kernel[3][3] ~^ image[21][17] + kernel[3][4] ~^ image[21][18] + kernel[4][0] ~^ image[22][14] + kernel[4][1] ~^ image[22][15] + kernel[4][2] ~^ image[22][16] + kernel[4][3] ~^ image[22][17] + kernel[4][4] ~^ image[22][18];
assign xor_sum[18][15] = kernel[0][0] ~^ image[18][15] + kernel[0][1] ~^ image[18][16] + kernel[0][2] ~^ image[18][17] + kernel[0][3] ~^ image[18][18] + kernel[0][4] ~^ image[18][19] + kernel[1][0] ~^ image[19][15] + kernel[1][1] ~^ image[19][16] + kernel[1][2] ~^ image[19][17] + kernel[1][3] ~^ image[19][18] + kernel[1][4] ~^ image[19][19] + kernel[2][0] ~^ image[20][15] + kernel[2][1] ~^ image[20][16] + kernel[2][2] ~^ image[20][17] + kernel[2][3] ~^ image[20][18] + kernel[2][4] ~^ image[20][19] + kernel[3][0] ~^ image[21][15] + kernel[3][1] ~^ image[21][16] + kernel[3][2] ~^ image[21][17] + kernel[3][3] ~^ image[21][18] + kernel[3][4] ~^ image[21][19] + kernel[4][0] ~^ image[22][15] + kernel[4][1] ~^ image[22][16] + kernel[4][2] ~^ image[22][17] + kernel[4][3] ~^ image[22][18] + kernel[4][4] ~^ image[22][19];
assign xor_sum[18][16] = kernel[0][0] ~^ image[18][16] + kernel[0][1] ~^ image[18][17] + kernel[0][2] ~^ image[18][18] + kernel[0][3] ~^ image[18][19] + kernel[0][4] ~^ image[18][20] + kernel[1][0] ~^ image[19][16] + kernel[1][1] ~^ image[19][17] + kernel[1][2] ~^ image[19][18] + kernel[1][3] ~^ image[19][19] + kernel[1][4] ~^ image[19][20] + kernel[2][0] ~^ image[20][16] + kernel[2][1] ~^ image[20][17] + kernel[2][2] ~^ image[20][18] + kernel[2][3] ~^ image[20][19] + kernel[2][4] ~^ image[20][20] + kernel[3][0] ~^ image[21][16] + kernel[3][1] ~^ image[21][17] + kernel[3][2] ~^ image[21][18] + kernel[3][3] ~^ image[21][19] + kernel[3][4] ~^ image[21][20] + kernel[4][0] ~^ image[22][16] + kernel[4][1] ~^ image[22][17] + kernel[4][2] ~^ image[22][18] + kernel[4][3] ~^ image[22][19] + kernel[4][4] ~^ image[22][20];
assign xor_sum[18][17] = kernel[0][0] ~^ image[18][17] + kernel[0][1] ~^ image[18][18] + kernel[0][2] ~^ image[18][19] + kernel[0][3] ~^ image[18][20] + kernel[0][4] ~^ image[18][21] + kernel[1][0] ~^ image[19][17] + kernel[1][1] ~^ image[19][18] + kernel[1][2] ~^ image[19][19] + kernel[1][3] ~^ image[19][20] + kernel[1][4] ~^ image[19][21] + kernel[2][0] ~^ image[20][17] + kernel[2][1] ~^ image[20][18] + kernel[2][2] ~^ image[20][19] + kernel[2][3] ~^ image[20][20] + kernel[2][4] ~^ image[20][21] + kernel[3][0] ~^ image[21][17] + kernel[3][1] ~^ image[21][18] + kernel[3][2] ~^ image[21][19] + kernel[3][3] ~^ image[21][20] + kernel[3][4] ~^ image[21][21] + kernel[4][0] ~^ image[22][17] + kernel[4][1] ~^ image[22][18] + kernel[4][2] ~^ image[22][19] + kernel[4][3] ~^ image[22][20] + kernel[4][4] ~^ image[22][21];
assign xor_sum[18][18] = kernel[0][0] ~^ image[18][18] + kernel[0][1] ~^ image[18][19] + kernel[0][2] ~^ image[18][20] + kernel[0][3] ~^ image[18][21] + kernel[0][4] ~^ image[18][22] + kernel[1][0] ~^ image[19][18] + kernel[1][1] ~^ image[19][19] + kernel[1][2] ~^ image[19][20] + kernel[1][3] ~^ image[19][21] + kernel[1][4] ~^ image[19][22] + kernel[2][0] ~^ image[20][18] + kernel[2][1] ~^ image[20][19] + kernel[2][2] ~^ image[20][20] + kernel[2][3] ~^ image[20][21] + kernel[2][4] ~^ image[20][22] + kernel[3][0] ~^ image[21][18] + kernel[3][1] ~^ image[21][19] + kernel[3][2] ~^ image[21][20] + kernel[3][3] ~^ image[21][21] + kernel[3][4] ~^ image[21][22] + kernel[4][0] ~^ image[22][18] + kernel[4][1] ~^ image[22][19] + kernel[4][2] ~^ image[22][20] + kernel[4][3] ~^ image[22][21] + kernel[4][4] ~^ image[22][22];
assign xor_sum[18][19] = kernel[0][0] ~^ image[18][19] + kernel[0][1] ~^ image[18][20] + kernel[0][2] ~^ image[18][21] + kernel[0][3] ~^ image[18][22] + kernel[0][4] ~^ image[18][23] + kernel[1][0] ~^ image[19][19] + kernel[1][1] ~^ image[19][20] + kernel[1][2] ~^ image[19][21] + kernel[1][3] ~^ image[19][22] + kernel[1][4] ~^ image[19][23] + kernel[2][0] ~^ image[20][19] + kernel[2][1] ~^ image[20][20] + kernel[2][2] ~^ image[20][21] + kernel[2][3] ~^ image[20][22] + kernel[2][4] ~^ image[20][23] + kernel[3][0] ~^ image[21][19] + kernel[3][1] ~^ image[21][20] + kernel[3][2] ~^ image[21][21] + kernel[3][3] ~^ image[21][22] + kernel[3][4] ~^ image[21][23] + kernel[4][0] ~^ image[22][19] + kernel[4][1] ~^ image[22][20] + kernel[4][2] ~^ image[22][21] + kernel[4][3] ~^ image[22][22] + kernel[4][4] ~^ image[22][23];
assign xor_sum[18][20] = kernel[0][0] ~^ image[18][20] + kernel[0][1] ~^ image[18][21] + kernel[0][2] ~^ image[18][22] + kernel[0][3] ~^ image[18][23] + kernel[0][4] ~^ image[18][24] + kernel[1][0] ~^ image[19][20] + kernel[1][1] ~^ image[19][21] + kernel[1][2] ~^ image[19][22] + kernel[1][3] ~^ image[19][23] + kernel[1][4] ~^ image[19][24] + kernel[2][0] ~^ image[20][20] + kernel[2][1] ~^ image[20][21] + kernel[2][2] ~^ image[20][22] + kernel[2][3] ~^ image[20][23] + kernel[2][4] ~^ image[20][24] + kernel[3][0] ~^ image[21][20] + kernel[3][1] ~^ image[21][21] + kernel[3][2] ~^ image[21][22] + kernel[3][3] ~^ image[21][23] + kernel[3][4] ~^ image[21][24] + kernel[4][0] ~^ image[22][20] + kernel[4][1] ~^ image[22][21] + kernel[4][2] ~^ image[22][22] + kernel[4][3] ~^ image[22][23] + kernel[4][4] ~^ image[22][24];
assign xor_sum[18][21] = kernel[0][0] ~^ image[18][21] + kernel[0][1] ~^ image[18][22] + kernel[0][2] ~^ image[18][23] + kernel[0][3] ~^ image[18][24] + kernel[0][4] ~^ image[18][25] + kernel[1][0] ~^ image[19][21] + kernel[1][1] ~^ image[19][22] + kernel[1][2] ~^ image[19][23] + kernel[1][3] ~^ image[19][24] + kernel[1][4] ~^ image[19][25] + kernel[2][0] ~^ image[20][21] + kernel[2][1] ~^ image[20][22] + kernel[2][2] ~^ image[20][23] + kernel[2][3] ~^ image[20][24] + kernel[2][4] ~^ image[20][25] + kernel[3][0] ~^ image[21][21] + kernel[3][1] ~^ image[21][22] + kernel[3][2] ~^ image[21][23] + kernel[3][3] ~^ image[21][24] + kernel[3][4] ~^ image[21][25] + kernel[4][0] ~^ image[22][21] + kernel[4][1] ~^ image[22][22] + kernel[4][2] ~^ image[22][23] + kernel[4][3] ~^ image[22][24] + kernel[4][4] ~^ image[22][25];
assign xor_sum[18][22] = kernel[0][0] ~^ image[18][22] + kernel[0][1] ~^ image[18][23] + kernel[0][2] ~^ image[18][24] + kernel[0][3] ~^ image[18][25] + kernel[0][4] ~^ image[18][26] + kernel[1][0] ~^ image[19][22] + kernel[1][1] ~^ image[19][23] + kernel[1][2] ~^ image[19][24] + kernel[1][3] ~^ image[19][25] + kernel[1][4] ~^ image[19][26] + kernel[2][0] ~^ image[20][22] + kernel[2][1] ~^ image[20][23] + kernel[2][2] ~^ image[20][24] + kernel[2][3] ~^ image[20][25] + kernel[2][4] ~^ image[20][26] + kernel[3][0] ~^ image[21][22] + kernel[3][1] ~^ image[21][23] + kernel[3][2] ~^ image[21][24] + kernel[3][3] ~^ image[21][25] + kernel[3][4] ~^ image[21][26] + kernel[4][0] ~^ image[22][22] + kernel[4][1] ~^ image[22][23] + kernel[4][2] ~^ image[22][24] + kernel[4][3] ~^ image[22][25] + kernel[4][4] ~^ image[22][26];
assign xor_sum[18][23] = kernel[0][0] ~^ image[18][23] + kernel[0][1] ~^ image[18][24] + kernel[0][2] ~^ image[18][25] + kernel[0][3] ~^ image[18][26] + kernel[0][4] ~^ image[18][27] + kernel[1][0] ~^ image[19][23] + kernel[1][1] ~^ image[19][24] + kernel[1][2] ~^ image[19][25] + kernel[1][3] ~^ image[19][26] + kernel[1][4] ~^ image[19][27] + kernel[2][0] ~^ image[20][23] + kernel[2][1] ~^ image[20][24] + kernel[2][2] ~^ image[20][25] + kernel[2][3] ~^ image[20][26] + kernel[2][4] ~^ image[20][27] + kernel[3][0] ~^ image[21][23] + kernel[3][1] ~^ image[21][24] + kernel[3][2] ~^ image[21][25] + kernel[3][3] ~^ image[21][26] + kernel[3][4] ~^ image[21][27] + kernel[4][0] ~^ image[22][23] + kernel[4][1] ~^ image[22][24] + kernel[4][2] ~^ image[22][25] + kernel[4][3] ~^ image[22][26] + kernel[4][4] ~^ image[22][27];
assign xor_sum[19][0] = kernel[0][0] ~^ image[19][0] + kernel[0][1] ~^ image[19][1] + kernel[0][2] ~^ image[19][2] + kernel[0][3] ~^ image[19][3] + kernel[0][4] ~^ image[19][4] + kernel[1][0] ~^ image[20][0] + kernel[1][1] ~^ image[20][1] + kernel[1][2] ~^ image[20][2] + kernel[1][3] ~^ image[20][3] + kernel[1][4] ~^ image[20][4] + kernel[2][0] ~^ image[21][0] + kernel[2][1] ~^ image[21][1] + kernel[2][2] ~^ image[21][2] + kernel[2][3] ~^ image[21][3] + kernel[2][4] ~^ image[21][4] + kernel[3][0] ~^ image[22][0] + kernel[3][1] ~^ image[22][1] + kernel[3][2] ~^ image[22][2] + kernel[3][3] ~^ image[22][3] + kernel[3][4] ~^ image[22][4] + kernel[4][0] ~^ image[23][0] + kernel[4][1] ~^ image[23][1] + kernel[4][2] ~^ image[23][2] + kernel[4][3] ~^ image[23][3] + kernel[4][4] ~^ image[23][4];
assign xor_sum[19][1] = kernel[0][0] ~^ image[19][1] + kernel[0][1] ~^ image[19][2] + kernel[0][2] ~^ image[19][3] + kernel[0][3] ~^ image[19][4] + kernel[0][4] ~^ image[19][5] + kernel[1][0] ~^ image[20][1] + kernel[1][1] ~^ image[20][2] + kernel[1][2] ~^ image[20][3] + kernel[1][3] ~^ image[20][4] + kernel[1][4] ~^ image[20][5] + kernel[2][0] ~^ image[21][1] + kernel[2][1] ~^ image[21][2] + kernel[2][2] ~^ image[21][3] + kernel[2][3] ~^ image[21][4] + kernel[2][4] ~^ image[21][5] + kernel[3][0] ~^ image[22][1] + kernel[3][1] ~^ image[22][2] + kernel[3][2] ~^ image[22][3] + kernel[3][3] ~^ image[22][4] + kernel[3][4] ~^ image[22][5] + kernel[4][0] ~^ image[23][1] + kernel[4][1] ~^ image[23][2] + kernel[4][2] ~^ image[23][3] + kernel[4][3] ~^ image[23][4] + kernel[4][4] ~^ image[23][5];
assign xor_sum[19][2] = kernel[0][0] ~^ image[19][2] + kernel[0][1] ~^ image[19][3] + kernel[0][2] ~^ image[19][4] + kernel[0][3] ~^ image[19][5] + kernel[0][4] ~^ image[19][6] + kernel[1][0] ~^ image[20][2] + kernel[1][1] ~^ image[20][3] + kernel[1][2] ~^ image[20][4] + kernel[1][3] ~^ image[20][5] + kernel[1][4] ~^ image[20][6] + kernel[2][0] ~^ image[21][2] + kernel[2][1] ~^ image[21][3] + kernel[2][2] ~^ image[21][4] + kernel[2][3] ~^ image[21][5] + kernel[2][4] ~^ image[21][6] + kernel[3][0] ~^ image[22][2] + kernel[3][1] ~^ image[22][3] + kernel[3][2] ~^ image[22][4] + kernel[3][3] ~^ image[22][5] + kernel[3][4] ~^ image[22][6] + kernel[4][0] ~^ image[23][2] + kernel[4][1] ~^ image[23][3] + kernel[4][2] ~^ image[23][4] + kernel[4][3] ~^ image[23][5] + kernel[4][4] ~^ image[23][6];
assign xor_sum[19][3] = kernel[0][0] ~^ image[19][3] + kernel[0][1] ~^ image[19][4] + kernel[0][2] ~^ image[19][5] + kernel[0][3] ~^ image[19][6] + kernel[0][4] ~^ image[19][7] + kernel[1][0] ~^ image[20][3] + kernel[1][1] ~^ image[20][4] + kernel[1][2] ~^ image[20][5] + kernel[1][3] ~^ image[20][6] + kernel[1][4] ~^ image[20][7] + kernel[2][0] ~^ image[21][3] + kernel[2][1] ~^ image[21][4] + kernel[2][2] ~^ image[21][5] + kernel[2][3] ~^ image[21][6] + kernel[2][4] ~^ image[21][7] + kernel[3][0] ~^ image[22][3] + kernel[3][1] ~^ image[22][4] + kernel[3][2] ~^ image[22][5] + kernel[3][3] ~^ image[22][6] + kernel[3][4] ~^ image[22][7] + kernel[4][0] ~^ image[23][3] + kernel[4][1] ~^ image[23][4] + kernel[4][2] ~^ image[23][5] + kernel[4][3] ~^ image[23][6] + kernel[4][4] ~^ image[23][7];
assign xor_sum[19][4] = kernel[0][0] ~^ image[19][4] + kernel[0][1] ~^ image[19][5] + kernel[0][2] ~^ image[19][6] + kernel[0][3] ~^ image[19][7] + kernel[0][4] ~^ image[19][8] + kernel[1][0] ~^ image[20][4] + kernel[1][1] ~^ image[20][5] + kernel[1][2] ~^ image[20][6] + kernel[1][3] ~^ image[20][7] + kernel[1][4] ~^ image[20][8] + kernel[2][0] ~^ image[21][4] + kernel[2][1] ~^ image[21][5] + kernel[2][2] ~^ image[21][6] + kernel[2][3] ~^ image[21][7] + kernel[2][4] ~^ image[21][8] + kernel[3][0] ~^ image[22][4] + kernel[3][1] ~^ image[22][5] + kernel[3][2] ~^ image[22][6] + kernel[3][3] ~^ image[22][7] + kernel[3][4] ~^ image[22][8] + kernel[4][0] ~^ image[23][4] + kernel[4][1] ~^ image[23][5] + kernel[4][2] ~^ image[23][6] + kernel[4][3] ~^ image[23][7] + kernel[4][4] ~^ image[23][8];
assign xor_sum[19][5] = kernel[0][0] ~^ image[19][5] + kernel[0][1] ~^ image[19][6] + kernel[0][2] ~^ image[19][7] + kernel[0][3] ~^ image[19][8] + kernel[0][4] ~^ image[19][9] + kernel[1][0] ~^ image[20][5] + kernel[1][1] ~^ image[20][6] + kernel[1][2] ~^ image[20][7] + kernel[1][3] ~^ image[20][8] + kernel[1][4] ~^ image[20][9] + kernel[2][0] ~^ image[21][5] + kernel[2][1] ~^ image[21][6] + kernel[2][2] ~^ image[21][7] + kernel[2][3] ~^ image[21][8] + kernel[2][4] ~^ image[21][9] + kernel[3][0] ~^ image[22][5] + kernel[3][1] ~^ image[22][6] + kernel[3][2] ~^ image[22][7] + kernel[3][3] ~^ image[22][8] + kernel[3][4] ~^ image[22][9] + kernel[4][0] ~^ image[23][5] + kernel[4][1] ~^ image[23][6] + kernel[4][2] ~^ image[23][7] + kernel[4][3] ~^ image[23][8] + kernel[4][4] ~^ image[23][9];
assign xor_sum[19][6] = kernel[0][0] ~^ image[19][6] + kernel[0][1] ~^ image[19][7] + kernel[0][2] ~^ image[19][8] + kernel[0][3] ~^ image[19][9] + kernel[0][4] ~^ image[19][10] + kernel[1][0] ~^ image[20][6] + kernel[1][1] ~^ image[20][7] + kernel[1][2] ~^ image[20][8] + kernel[1][3] ~^ image[20][9] + kernel[1][4] ~^ image[20][10] + kernel[2][0] ~^ image[21][6] + kernel[2][1] ~^ image[21][7] + kernel[2][2] ~^ image[21][8] + kernel[2][3] ~^ image[21][9] + kernel[2][4] ~^ image[21][10] + kernel[3][0] ~^ image[22][6] + kernel[3][1] ~^ image[22][7] + kernel[3][2] ~^ image[22][8] + kernel[3][3] ~^ image[22][9] + kernel[3][4] ~^ image[22][10] + kernel[4][0] ~^ image[23][6] + kernel[4][1] ~^ image[23][7] + kernel[4][2] ~^ image[23][8] + kernel[4][3] ~^ image[23][9] + kernel[4][4] ~^ image[23][10];
assign xor_sum[19][7] = kernel[0][0] ~^ image[19][7] + kernel[0][1] ~^ image[19][8] + kernel[0][2] ~^ image[19][9] + kernel[0][3] ~^ image[19][10] + kernel[0][4] ~^ image[19][11] + kernel[1][0] ~^ image[20][7] + kernel[1][1] ~^ image[20][8] + kernel[1][2] ~^ image[20][9] + kernel[1][3] ~^ image[20][10] + kernel[1][4] ~^ image[20][11] + kernel[2][0] ~^ image[21][7] + kernel[2][1] ~^ image[21][8] + kernel[2][2] ~^ image[21][9] + kernel[2][3] ~^ image[21][10] + kernel[2][4] ~^ image[21][11] + kernel[3][0] ~^ image[22][7] + kernel[3][1] ~^ image[22][8] + kernel[3][2] ~^ image[22][9] + kernel[3][3] ~^ image[22][10] + kernel[3][4] ~^ image[22][11] + kernel[4][0] ~^ image[23][7] + kernel[4][1] ~^ image[23][8] + kernel[4][2] ~^ image[23][9] + kernel[4][3] ~^ image[23][10] + kernel[4][4] ~^ image[23][11];
assign xor_sum[19][8] = kernel[0][0] ~^ image[19][8] + kernel[0][1] ~^ image[19][9] + kernel[0][2] ~^ image[19][10] + kernel[0][3] ~^ image[19][11] + kernel[0][4] ~^ image[19][12] + kernel[1][0] ~^ image[20][8] + kernel[1][1] ~^ image[20][9] + kernel[1][2] ~^ image[20][10] + kernel[1][3] ~^ image[20][11] + kernel[1][4] ~^ image[20][12] + kernel[2][0] ~^ image[21][8] + kernel[2][1] ~^ image[21][9] + kernel[2][2] ~^ image[21][10] + kernel[2][3] ~^ image[21][11] + kernel[2][4] ~^ image[21][12] + kernel[3][0] ~^ image[22][8] + kernel[3][1] ~^ image[22][9] + kernel[3][2] ~^ image[22][10] + kernel[3][3] ~^ image[22][11] + kernel[3][4] ~^ image[22][12] + kernel[4][0] ~^ image[23][8] + kernel[4][1] ~^ image[23][9] + kernel[4][2] ~^ image[23][10] + kernel[4][3] ~^ image[23][11] + kernel[4][4] ~^ image[23][12];
assign xor_sum[19][9] = kernel[0][0] ~^ image[19][9] + kernel[0][1] ~^ image[19][10] + kernel[0][2] ~^ image[19][11] + kernel[0][3] ~^ image[19][12] + kernel[0][4] ~^ image[19][13] + kernel[1][0] ~^ image[20][9] + kernel[1][1] ~^ image[20][10] + kernel[1][2] ~^ image[20][11] + kernel[1][3] ~^ image[20][12] + kernel[1][4] ~^ image[20][13] + kernel[2][0] ~^ image[21][9] + kernel[2][1] ~^ image[21][10] + kernel[2][2] ~^ image[21][11] + kernel[2][3] ~^ image[21][12] + kernel[2][4] ~^ image[21][13] + kernel[3][0] ~^ image[22][9] + kernel[3][1] ~^ image[22][10] + kernel[3][2] ~^ image[22][11] + kernel[3][3] ~^ image[22][12] + kernel[3][4] ~^ image[22][13] + kernel[4][0] ~^ image[23][9] + kernel[4][1] ~^ image[23][10] + kernel[4][2] ~^ image[23][11] + kernel[4][3] ~^ image[23][12] + kernel[4][4] ~^ image[23][13];
assign xor_sum[19][10] = kernel[0][0] ~^ image[19][10] + kernel[0][1] ~^ image[19][11] + kernel[0][2] ~^ image[19][12] + kernel[0][3] ~^ image[19][13] + kernel[0][4] ~^ image[19][14] + kernel[1][0] ~^ image[20][10] + kernel[1][1] ~^ image[20][11] + kernel[1][2] ~^ image[20][12] + kernel[1][3] ~^ image[20][13] + kernel[1][4] ~^ image[20][14] + kernel[2][0] ~^ image[21][10] + kernel[2][1] ~^ image[21][11] + kernel[2][2] ~^ image[21][12] + kernel[2][3] ~^ image[21][13] + kernel[2][4] ~^ image[21][14] + kernel[3][0] ~^ image[22][10] + kernel[3][1] ~^ image[22][11] + kernel[3][2] ~^ image[22][12] + kernel[3][3] ~^ image[22][13] + kernel[3][4] ~^ image[22][14] + kernel[4][0] ~^ image[23][10] + kernel[4][1] ~^ image[23][11] + kernel[4][2] ~^ image[23][12] + kernel[4][3] ~^ image[23][13] + kernel[4][4] ~^ image[23][14];
assign xor_sum[19][11] = kernel[0][0] ~^ image[19][11] + kernel[0][1] ~^ image[19][12] + kernel[0][2] ~^ image[19][13] + kernel[0][3] ~^ image[19][14] + kernel[0][4] ~^ image[19][15] + kernel[1][0] ~^ image[20][11] + kernel[1][1] ~^ image[20][12] + kernel[1][2] ~^ image[20][13] + kernel[1][3] ~^ image[20][14] + kernel[1][4] ~^ image[20][15] + kernel[2][0] ~^ image[21][11] + kernel[2][1] ~^ image[21][12] + kernel[2][2] ~^ image[21][13] + kernel[2][3] ~^ image[21][14] + kernel[2][4] ~^ image[21][15] + kernel[3][0] ~^ image[22][11] + kernel[3][1] ~^ image[22][12] + kernel[3][2] ~^ image[22][13] + kernel[3][3] ~^ image[22][14] + kernel[3][4] ~^ image[22][15] + kernel[4][0] ~^ image[23][11] + kernel[4][1] ~^ image[23][12] + kernel[4][2] ~^ image[23][13] + kernel[4][3] ~^ image[23][14] + kernel[4][4] ~^ image[23][15];
assign xor_sum[19][12] = kernel[0][0] ~^ image[19][12] + kernel[0][1] ~^ image[19][13] + kernel[0][2] ~^ image[19][14] + kernel[0][3] ~^ image[19][15] + kernel[0][4] ~^ image[19][16] + kernel[1][0] ~^ image[20][12] + kernel[1][1] ~^ image[20][13] + kernel[1][2] ~^ image[20][14] + kernel[1][3] ~^ image[20][15] + kernel[1][4] ~^ image[20][16] + kernel[2][0] ~^ image[21][12] + kernel[2][1] ~^ image[21][13] + kernel[2][2] ~^ image[21][14] + kernel[2][3] ~^ image[21][15] + kernel[2][4] ~^ image[21][16] + kernel[3][0] ~^ image[22][12] + kernel[3][1] ~^ image[22][13] + kernel[3][2] ~^ image[22][14] + kernel[3][3] ~^ image[22][15] + kernel[3][4] ~^ image[22][16] + kernel[4][0] ~^ image[23][12] + kernel[4][1] ~^ image[23][13] + kernel[4][2] ~^ image[23][14] + kernel[4][3] ~^ image[23][15] + kernel[4][4] ~^ image[23][16];
assign xor_sum[19][13] = kernel[0][0] ~^ image[19][13] + kernel[0][1] ~^ image[19][14] + kernel[0][2] ~^ image[19][15] + kernel[0][3] ~^ image[19][16] + kernel[0][4] ~^ image[19][17] + kernel[1][0] ~^ image[20][13] + kernel[1][1] ~^ image[20][14] + kernel[1][2] ~^ image[20][15] + kernel[1][3] ~^ image[20][16] + kernel[1][4] ~^ image[20][17] + kernel[2][0] ~^ image[21][13] + kernel[2][1] ~^ image[21][14] + kernel[2][2] ~^ image[21][15] + kernel[2][3] ~^ image[21][16] + kernel[2][4] ~^ image[21][17] + kernel[3][0] ~^ image[22][13] + kernel[3][1] ~^ image[22][14] + kernel[3][2] ~^ image[22][15] + kernel[3][3] ~^ image[22][16] + kernel[3][4] ~^ image[22][17] + kernel[4][0] ~^ image[23][13] + kernel[4][1] ~^ image[23][14] + kernel[4][2] ~^ image[23][15] + kernel[4][3] ~^ image[23][16] + kernel[4][4] ~^ image[23][17];
assign xor_sum[19][14] = kernel[0][0] ~^ image[19][14] + kernel[0][1] ~^ image[19][15] + kernel[0][2] ~^ image[19][16] + kernel[0][3] ~^ image[19][17] + kernel[0][4] ~^ image[19][18] + kernel[1][0] ~^ image[20][14] + kernel[1][1] ~^ image[20][15] + kernel[1][2] ~^ image[20][16] + kernel[1][3] ~^ image[20][17] + kernel[1][4] ~^ image[20][18] + kernel[2][0] ~^ image[21][14] + kernel[2][1] ~^ image[21][15] + kernel[2][2] ~^ image[21][16] + kernel[2][3] ~^ image[21][17] + kernel[2][4] ~^ image[21][18] + kernel[3][0] ~^ image[22][14] + kernel[3][1] ~^ image[22][15] + kernel[3][2] ~^ image[22][16] + kernel[3][3] ~^ image[22][17] + kernel[3][4] ~^ image[22][18] + kernel[4][0] ~^ image[23][14] + kernel[4][1] ~^ image[23][15] + kernel[4][2] ~^ image[23][16] + kernel[4][3] ~^ image[23][17] + kernel[4][4] ~^ image[23][18];
assign xor_sum[19][15] = kernel[0][0] ~^ image[19][15] + kernel[0][1] ~^ image[19][16] + kernel[0][2] ~^ image[19][17] + kernel[0][3] ~^ image[19][18] + kernel[0][4] ~^ image[19][19] + kernel[1][0] ~^ image[20][15] + kernel[1][1] ~^ image[20][16] + kernel[1][2] ~^ image[20][17] + kernel[1][3] ~^ image[20][18] + kernel[1][4] ~^ image[20][19] + kernel[2][0] ~^ image[21][15] + kernel[2][1] ~^ image[21][16] + kernel[2][2] ~^ image[21][17] + kernel[2][3] ~^ image[21][18] + kernel[2][4] ~^ image[21][19] + kernel[3][0] ~^ image[22][15] + kernel[3][1] ~^ image[22][16] + kernel[3][2] ~^ image[22][17] + kernel[3][3] ~^ image[22][18] + kernel[3][4] ~^ image[22][19] + kernel[4][0] ~^ image[23][15] + kernel[4][1] ~^ image[23][16] + kernel[4][2] ~^ image[23][17] + kernel[4][3] ~^ image[23][18] + kernel[4][4] ~^ image[23][19];
assign xor_sum[19][16] = kernel[0][0] ~^ image[19][16] + kernel[0][1] ~^ image[19][17] + kernel[0][2] ~^ image[19][18] + kernel[0][3] ~^ image[19][19] + kernel[0][4] ~^ image[19][20] + kernel[1][0] ~^ image[20][16] + kernel[1][1] ~^ image[20][17] + kernel[1][2] ~^ image[20][18] + kernel[1][3] ~^ image[20][19] + kernel[1][4] ~^ image[20][20] + kernel[2][0] ~^ image[21][16] + kernel[2][1] ~^ image[21][17] + kernel[2][2] ~^ image[21][18] + kernel[2][3] ~^ image[21][19] + kernel[2][4] ~^ image[21][20] + kernel[3][0] ~^ image[22][16] + kernel[3][1] ~^ image[22][17] + kernel[3][2] ~^ image[22][18] + kernel[3][3] ~^ image[22][19] + kernel[3][4] ~^ image[22][20] + kernel[4][0] ~^ image[23][16] + kernel[4][1] ~^ image[23][17] + kernel[4][2] ~^ image[23][18] + kernel[4][3] ~^ image[23][19] + kernel[4][4] ~^ image[23][20];
assign xor_sum[19][17] = kernel[0][0] ~^ image[19][17] + kernel[0][1] ~^ image[19][18] + kernel[0][2] ~^ image[19][19] + kernel[0][3] ~^ image[19][20] + kernel[0][4] ~^ image[19][21] + kernel[1][0] ~^ image[20][17] + kernel[1][1] ~^ image[20][18] + kernel[1][2] ~^ image[20][19] + kernel[1][3] ~^ image[20][20] + kernel[1][4] ~^ image[20][21] + kernel[2][0] ~^ image[21][17] + kernel[2][1] ~^ image[21][18] + kernel[2][2] ~^ image[21][19] + kernel[2][3] ~^ image[21][20] + kernel[2][4] ~^ image[21][21] + kernel[3][0] ~^ image[22][17] + kernel[3][1] ~^ image[22][18] + kernel[3][2] ~^ image[22][19] + kernel[3][3] ~^ image[22][20] + kernel[3][4] ~^ image[22][21] + kernel[4][0] ~^ image[23][17] + kernel[4][1] ~^ image[23][18] + kernel[4][2] ~^ image[23][19] + kernel[4][3] ~^ image[23][20] + kernel[4][4] ~^ image[23][21];
assign xor_sum[19][18] = kernel[0][0] ~^ image[19][18] + kernel[0][1] ~^ image[19][19] + kernel[0][2] ~^ image[19][20] + kernel[0][3] ~^ image[19][21] + kernel[0][4] ~^ image[19][22] + kernel[1][0] ~^ image[20][18] + kernel[1][1] ~^ image[20][19] + kernel[1][2] ~^ image[20][20] + kernel[1][3] ~^ image[20][21] + kernel[1][4] ~^ image[20][22] + kernel[2][0] ~^ image[21][18] + kernel[2][1] ~^ image[21][19] + kernel[2][2] ~^ image[21][20] + kernel[2][3] ~^ image[21][21] + kernel[2][4] ~^ image[21][22] + kernel[3][0] ~^ image[22][18] + kernel[3][1] ~^ image[22][19] + kernel[3][2] ~^ image[22][20] + kernel[3][3] ~^ image[22][21] + kernel[3][4] ~^ image[22][22] + kernel[4][0] ~^ image[23][18] + kernel[4][1] ~^ image[23][19] + kernel[4][2] ~^ image[23][20] + kernel[4][3] ~^ image[23][21] + kernel[4][4] ~^ image[23][22];
assign xor_sum[19][19] = kernel[0][0] ~^ image[19][19] + kernel[0][1] ~^ image[19][20] + kernel[0][2] ~^ image[19][21] + kernel[0][3] ~^ image[19][22] + kernel[0][4] ~^ image[19][23] + kernel[1][0] ~^ image[20][19] + kernel[1][1] ~^ image[20][20] + kernel[1][2] ~^ image[20][21] + kernel[1][3] ~^ image[20][22] + kernel[1][4] ~^ image[20][23] + kernel[2][0] ~^ image[21][19] + kernel[2][1] ~^ image[21][20] + kernel[2][2] ~^ image[21][21] + kernel[2][3] ~^ image[21][22] + kernel[2][4] ~^ image[21][23] + kernel[3][0] ~^ image[22][19] + kernel[3][1] ~^ image[22][20] + kernel[3][2] ~^ image[22][21] + kernel[3][3] ~^ image[22][22] + kernel[3][4] ~^ image[22][23] + kernel[4][0] ~^ image[23][19] + kernel[4][1] ~^ image[23][20] + kernel[4][2] ~^ image[23][21] + kernel[4][3] ~^ image[23][22] + kernel[4][4] ~^ image[23][23];
assign xor_sum[19][20] = kernel[0][0] ~^ image[19][20] + kernel[0][1] ~^ image[19][21] + kernel[0][2] ~^ image[19][22] + kernel[0][3] ~^ image[19][23] + kernel[0][4] ~^ image[19][24] + kernel[1][0] ~^ image[20][20] + kernel[1][1] ~^ image[20][21] + kernel[1][2] ~^ image[20][22] + kernel[1][3] ~^ image[20][23] + kernel[1][4] ~^ image[20][24] + kernel[2][0] ~^ image[21][20] + kernel[2][1] ~^ image[21][21] + kernel[2][2] ~^ image[21][22] + kernel[2][3] ~^ image[21][23] + kernel[2][4] ~^ image[21][24] + kernel[3][0] ~^ image[22][20] + kernel[3][1] ~^ image[22][21] + kernel[3][2] ~^ image[22][22] + kernel[3][3] ~^ image[22][23] + kernel[3][4] ~^ image[22][24] + kernel[4][0] ~^ image[23][20] + kernel[4][1] ~^ image[23][21] + kernel[4][2] ~^ image[23][22] + kernel[4][3] ~^ image[23][23] + kernel[4][4] ~^ image[23][24];
assign xor_sum[19][21] = kernel[0][0] ~^ image[19][21] + kernel[0][1] ~^ image[19][22] + kernel[0][2] ~^ image[19][23] + kernel[0][3] ~^ image[19][24] + kernel[0][4] ~^ image[19][25] + kernel[1][0] ~^ image[20][21] + kernel[1][1] ~^ image[20][22] + kernel[1][2] ~^ image[20][23] + kernel[1][3] ~^ image[20][24] + kernel[1][4] ~^ image[20][25] + kernel[2][0] ~^ image[21][21] + kernel[2][1] ~^ image[21][22] + kernel[2][2] ~^ image[21][23] + kernel[2][3] ~^ image[21][24] + kernel[2][4] ~^ image[21][25] + kernel[3][0] ~^ image[22][21] + kernel[3][1] ~^ image[22][22] + kernel[3][2] ~^ image[22][23] + kernel[3][3] ~^ image[22][24] + kernel[3][4] ~^ image[22][25] + kernel[4][0] ~^ image[23][21] + kernel[4][1] ~^ image[23][22] + kernel[4][2] ~^ image[23][23] + kernel[4][3] ~^ image[23][24] + kernel[4][4] ~^ image[23][25];
assign xor_sum[19][22] = kernel[0][0] ~^ image[19][22] + kernel[0][1] ~^ image[19][23] + kernel[0][2] ~^ image[19][24] + kernel[0][3] ~^ image[19][25] + kernel[0][4] ~^ image[19][26] + kernel[1][0] ~^ image[20][22] + kernel[1][1] ~^ image[20][23] + kernel[1][2] ~^ image[20][24] + kernel[1][3] ~^ image[20][25] + kernel[1][4] ~^ image[20][26] + kernel[2][0] ~^ image[21][22] + kernel[2][1] ~^ image[21][23] + kernel[2][2] ~^ image[21][24] + kernel[2][3] ~^ image[21][25] + kernel[2][4] ~^ image[21][26] + kernel[3][0] ~^ image[22][22] + kernel[3][1] ~^ image[22][23] + kernel[3][2] ~^ image[22][24] + kernel[3][3] ~^ image[22][25] + kernel[3][4] ~^ image[22][26] + kernel[4][0] ~^ image[23][22] + kernel[4][1] ~^ image[23][23] + kernel[4][2] ~^ image[23][24] + kernel[4][3] ~^ image[23][25] + kernel[4][4] ~^ image[23][26];
assign xor_sum[19][23] = kernel[0][0] ~^ image[19][23] + kernel[0][1] ~^ image[19][24] + kernel[0][2] ~^ image[19][25] + kernel[0][3] ~^ image[19][26] + kernel[0][4] ~^ image[19][27] + kernel[1][0] ~^ image[20][23] + kernel[1][1] ~^ image[20][24] + kernel[1][2] ~^ image[20][25] + kernel[1][3] ~^ image[20][26] + kernel[1][4] ~^ image[20][27] + kernel[2][0] ~^ image[21][23] + kernel[2][1] ~^ image[21][24] + kernel[2][2] ~^ image[21][25] + kernel[2][3] ~^ image[21][26] + kernel[2][4] ~^ image[21][27] + kernel[3][0] ~^ image[22][23] + kernel[3][1] ~^ image[22][24] + kernel[3][2] ~^ image[22][25] + kernel[3][3] ~^ image[22][26] + kernel[3][4] ~^ image[22][27] + kernel[4][0] ~^ image[23][23] + kernel[4][1] ~^ image[23][24] + kernel[4][2] ~^ image[23][25] + kernel[4][3] ~^ image[23][26] + kernel[4][4] ~^ image[23][27];
assign xor_sum[20][0] = kernel[0][0] ~^ image[20][0] + kernel[0][1] ~^ image[20][1] + kernel[0][2] ~^ image[20][2] + kernel[0][3] ~^ image[20][3] + kernel[0][4] ~^ image[20][4] + kernel[1][0] ~^ image[21][0] + kernel[1][1] ~^ image[21][1] + kernel[1][2] ~^ image[21][2] + kernel[1][3] ~^ image[21][3] + kernel[1][4] ~^ image[21][4] + kernel[2][0] ~^ image[22][0] + kernel[2][1] ~^ image[22][1] + kernel[2][2] ~^ image[22][2] + kernel[2][3] ~^ image[22][3] + kernel[2][4] ~^ image[22][4] + kernel[3][0] ~^ image[23][0] + kernel[3][1] ~^ image[23][1] + kernel[3][2] ~^ image[23][2] + kernel[3][3] ~^ image[23][3] + kernel[3][4] ~^ image[23][4] + kernel[4][0] ~^ image[24][0] + kernel[4][1] ~^ image[24][1] + kernel[4][2] ~^ image[24][2] + kernel[4][3] ~^ image[24][3] + kernel[4][4] ~^ image[24][4];
assign xor_sum[20][1] = kernel[0][0] ~^ image[20][1] + kernel[0][1] ~^ image[20][2] + kernel[0][2] ~^ image[20][3] + kernel[0][3] ~^ image[20][4] + kernel[0][4] ~^ image[20][5] + kernel[1][0] ~^ image[21][1] + kernel[1][1] ~^ image[21][2] + kernel[1][2] ~^ image[21][3] + kernel[1][3] ~^ image[21][4] + kernel[1][4] ~^ image[21][5] + kernel[2][0] ~^ image[22][1] + kernel[2][1] ~^ image[22][2] + kernel[2][2] ~^ image[22][3] + kernel[2][3] ~^ image[22][4] + kernel[2][4] ~^ image[22][5] + kernel[3][0] ~^ image[23][1] + kernel[3][1] ~^ image[23][2] + kernel[3][2] ~^ image[23][3] + kernel[3][3] ~^ image[23][4] + kernel[3][4] ~^ image[23][5] + kernel[4][0] ~^ image[24][1] + kernel[4][1] ~^ image[24][2] + kernel[4][2] ~^ image[24][3] + kernel[4][3] ~^ image[24][4] + kernel[4][4] ~^ image[24][5];
assign xor_sum[20][2] = kernel[0][0] ~^ image[20][2] + kernel[0][1] ~^ image[20][3] + kernel[0][2] ~^ image[20][4] + kernel[0][3] ~^ image[20][5] + kernel[0][4] ~^ image[20][6] + kernel[1][0] ~^ image[21][2] + kernel[1][1] ~^ image[21][3] + kernel[1][2] ~^ image[21][4] + kernel[1][3] ~^ image[21][5] + kernel[1][4] ~^ image[21][6] + kernel[2][0] ~^ image[22][2] + kernel[2][1] ~^ image[22][3] + kernel[2][2] ~^ image[22][4] + kernel[2][3] ~^ image[22][5] + kernel[2][4] ~^ image[22][6] + kernel[3][0] ~^ image[23][2] + kernel[3][1] ~^ image[23][3] + kernel[3][2] ~^ image[23][4] + kernel[3][3] ~^ image[23][5] + kernel[3][4] ~^ image[23][6] + kernel[4][0] ~^ image[24][2] + kernel[4][1] ~^ image[24][3] + kernel[4][2] ~^ image[24][4] + kernel[4][3] ~^ image[24][5] + kernel[4][4] ~^ image[24][6];
assign xor_sum[20][3] = kernel[0][0] ~^ image[20][3] + kernel[0][1] ~^ image[20][4] + kernel[0][2] ~^ image[20][5] + kernel[0][3] ~^ image[20][6] + kernel[0][4] ~^ image[20][7] + kernel[1][0] ~^ image[21][3] + kernel[1][1] ~^ image[21][4] + kernel[1][2] ~^ image[21][5] + kernel[1][3] ~^ image[21][6] + kernel[1][4] ~^ image[21][7] + kernel[2][0] ~^ image[22][3] + kernel[2][1] ~^ image[22][4] + kernel[2][2] ~^ image[22][5] + kernel[2][3] ~^ image[22][6] + kernel[2][4] ~^ image[22][7] + kernel[3][0] ~^ image[23][3] + kernel[3][1] ~^ image[23][4] + kernel[3][2] ~^ image[23][5] + kernel[3][3] ~^ image[23][6] + kernel[3][4] ~^ image[23][7] + kernel[4][0] ~^ image[24][3] + kernel[4][1] ~^ image[24][4] + kernel[4][2] ~^ image[24][5] + kernel[4][3] ~^ image[24][6] + kernel[4][4] ~^ image[24][7];
assign xor_sum[20][4] = kernel[0][0] ~^ image[20][4] + kernel[0][1] ~^ image[20][5] + kernel[0][2] ~^ image[20][6] + kernel[0][3] ~^ image[20][7] + kernel[0][4] ~^ image[20][8] + kernel[1][0] ~^ image[21][4] + kernel[1][1] ~^ image[21][5] + kernel[1][2] ~^ image[21][6] + kernel[1][3] ~^ image[21][7] + kernel[1][4] ~^ image[21][8] + kernel[2][0] ~^ image[22][4] + kernel[2][1] ~^ image[22][5] + kernel[2][2] ~^ image[22][6] + kernel[2][3] ~^ image[22][7] + kernel[2][4] ~^ image[22][8] + kernel[3][0] ~^ image[23][4] + kernel[3][1] ~^ image[23][5] + kernel[3][2] ~^ image[23][6] + kernel[3][3] ~^ image[23][7] + kernel[3][4] ~^ image[23][8] + kernel[4][0] ~^ image[24][4] + kernel[4][1] ~^ image[24][5] + kernel[4][2] ~^ image[24][6] + kernel[4][3] ~^ image[24][7] + kernel[4][4] ~^ image[24][8];
assign xor_sum[20][5] = kernel[0][0] ~^ image[20][5] + kernel[0][1] ~^ image[20][6] + kernel[0][2] ~^ image[20][7] + kernel[0][3] ~^ image[20][8] + kernel[0][4] ~^ image[20][9] + kernel[1][0] ~^ image[21][5] + kernel[1][1] ~^ image[21][6] + kernel[1][2] ~^ image[21][7] + kernel[1][3] ~^ image[21][8] + kernel[1][4] ~^ image[21][9] + kernel[2][0] ~^ image[22][5] + kernel[2][1] ~^ image[22][6] + kernel[2][2] ~^ image[22][7] + kernel[2][3] ~^ image[22][8] + kernel[2][4] ~^ image[22][9] + kernel[3][0] ~^ image[23][5] + kernel[3][1] ~^ image[23][6] + kernel[3][2] ~^ image[23][7] + kernel[3][3] ~^ image[23][8] + kernel[3][4] ~^ image[23][9] + kernel[4][0] ~^ image[24][5] + kernel[4][1] ~^ image[24][6] + kernel[4][2] ~^ image[24][7] + kernel[4][3] ~^ image[24][8] + kernel[4][4] ~^ image[24][9];
assign xor_sum[20][6] = kernel[0][0] ~^ image[20][6] + kernel[0][1] ~^ image[20][7] + kernel[0][2] ~^ image[20][8] + kernel[0][3] ~^ image[20][9] + kernel[0][4] ~^ image[20][10] + kernel[1][0] ~^ image[21][6] + kernel[1][1] ~^ image[21][7] + kernel[1][2] ~^ image[21][8] + kernel[1][3] ~^ image[21][9] + kernel[1][4] ~^ image[21][10] + kernel[2][0] ~^ image[22][6] + kernel[2][1] ~^ image[22][7] + kernel[2][2] ~^ image[22][8] + kernel[2][3] ~^ image[22][9] + kernel[2][4] ~^ image[22][10] + kernel[3][0] ~^ image[23][6] + kernel[3][1] ~^ image[23][7] + kernel[3][2] ~^ image[23][8] + kernel[3][3] ~^ image[23][9] + kernel[3][4] ~^ image[23][10] + kernel[4][0] ~^ image[24][6] + kernel[4][1] ~^ image[24][7] + kernel[4][2] ~^ image[24][8] + kernel[4][3] ~^ image[24][9] + kernel[4][4] ~^ image[24][10];
assign xor_sum[20][7] = kernel[0][0] ~^ image[20][7] + kernel[0][1] ~^ image[20][8] + kernel[0][2] ~^ image[20][9] + kernel[0][3] ~^ image[20][10] + kernel[0][4] ~^ image[20][11] + kernel[1][0] ~^ image[21][7] + kernel[1][1] ~^ image[21][8] + kernel[1][2] ~^ image[21][9] + kernel[1][3] ~^ image[21][10] + kernel[1][4] ~^ image[21][11] + kernel[2][0] ~^ image[22][7] + kernel[2][1] ~^ image[22][8] + kernel[2][2] ~^ image[22][9] + kernel[2][3] ~^ image[22][10] + kernel[2][4] ~^ image[22][11] + kernel[3][0] ~^ image[23][7] + kernel[3][1] ~^ image[23][8] + kernel[3][2] ~^ image[23][9] + kernel[3][3] ~^ image[23][10] + kernel[3][4] ~^ image[23][11] + kernel[4][0] ~^ image[24][7] + kernel[4][1] ~^ image[24][8] + kernel[4][2] ~^ image[24][9] + kernel[4][3] ~^ image[24][10] + kernel[4][4] ~^ image[24][11];
assign xor_sum[20][8] = kernel[0][0] ~^ image[20][8] + kernel[0][1] ~^ image[20][9] + kernel[0][2] ~^ image[20][10] + kernel[0][3] ~^ image[20][11] + kernel[0][4] ~^ image[20][12] + kernel[1][0] ~^ image[21][8] + kernel[1][1] ~^ image[21][9] + kernel[1][2] ~^ image[21][10] + kernel[1][3] ~^ image[21][11] + kernel[1][4] ~^ image[21][12] + kernel[2][0] ~^ image[22][8] + kernel[2][1] ~^ image[22][9] + kernel[2][2] ~^ image[22][10] + kernel[2][3] ~^ image[22][11] + kernel[2][4] ~^ image[22][12] + kernel[3][0] ~^ image[23][8] + kernel[3][1] ~^ image[23][9] + kernel[3][2] ~^ image[23][10] + kernel[3][3] ~^ image[23][11] + kernel[3][4] ~^ image[23][12] + kernel[4][0] ~^ image[24][8] + kernel[4][1] ~^ image[24][9] + kernel[4][2] ~^ image[24][10] + kernel[4][3] ~^ image[24][11] + kernel[4][4] ~^ image[24][12];
assign xor_sum[20][9] = kernel[0][0] ~^ image[20][9] + kernel[0][1] ~^ image[20][10] + kernel[0][2] ~^ image[20][11] + kernel[0][3] ~^ image[20][12] + kernel[0][4] ~^ image[20][13] + kernel[1][0] ~^ image[21][9] + kernel[1][1] ~^ image[21][10] + kernel[1][2] ~^ image[21][11] + kernel[1][3] ~^ image[21][12] + kernel[1][4] ~^ image[21][13] + kernel[2][0] ~^ image[22][9] + kernel[2][1] ~^ image[22][10] + kernel[2][2] ~^ image[22][11] + kernel[2][3] ~^ image[22][12] + kernel[2][4] ~^ image[22][13] + kernel[3][0] ~^ image[23][9] + kernel[3][1] ~^ image[23][10] + kernel[3][2] ~^ image[23][11] + kernel[3][3] ~^ image[23][12] + kernel[3][4] ~^ image[23][13] + kernel[4][0] ~^ image[24][9] + kernel[4][1] ~^ image[24][10] + kernel[4][2] ~^ image[24][11] + kernel[4][3] ~^ image[24][12] + kernel[4][4] ~^ image[24][13];
assign xor_sum[20][10] = kernel[0][0] ~^ image[20][10] + kernel[0][1] ~^ image[20][11] + kernel[0][2] ~^ image[20][12] + kernel[0][3] ~^ image[20][13] + kernel[0][4] ~^ image[20][14] + kernel[1][0] ~^ image[21][10] + kernel[1][1] ~^ image[21][11] + kernel[1][2] ~^ image[21][12] + kernel[1][3] ~^ image[21][13] + kernel[1][4] ~^ image[21][14] + kernel[2][0] ~^ image[22][10] + kernel[2][1] ~^ image[22][11] + kernel[2][2] ~^ image[22][12] + kernel[2][3] ~^ image[22][13] + kernel[2][4] ~^ image[22][14] + kernel[3][0] ~^ image[23][10] + kernel[3][1] ~^ image[23][11] + kernel[3][2] ~^ image[23][12] + kernel[3][3] ~^ image[23][13] + kernel[3][4] ~^ image[23][14] + kernel[4][0] ~^ image[24][10] + kernel[4][1] ~^ image[24][11] + kernel[4][2] ~^ image[24][12] + kernel[4][3] ~^ image[24][13] + kernel[4][4] ~^ image[24][14];
assign xor_sum[20][11] = kernel[0][0] ~^ image[20][11] + kernel[0][1] ~^ image[20][12] + kernel[0][2] ~^ image[20][13] + kernel[0][3] ~^ image[20][14] + kernel[0][4] ~^ image[20][15] + kernel[1][0] ~^ image[21][11] + kernel[1][1] ~^ image[21][12] + kernel[1][2] ~^ image[21][13] + kernel[1][3] ~^ image[21][14] + kernel[1][4] ~^ image[21][15] + kernel[2][0] ~^ image[22][11] + kernel[2][1] ~^ image[22][12] + kernel[2][2] ~^ image[22][13] + kernel[2][3] ~^ image[22][14] + kernel[2][4] ~^ image[22][15] + kernel[3][0] ~^ image[23][11] + kernel[3][1] ~^ image[23][12] + kernel[3][2] ~^ image[23][13] + kernel[3][3] ~^ image[23][14] + kernel[3][4] ~^ image[23][15] + kernel[4][0] ~^ image[24][11] + kernel[4][1] ~^ image[24][12] + kernel[4][2] ~^ image[24][13] + kernel[4][3] ~^ image[24][14] + kernel[4][4] ~^ image[24][15];
assign xor_sum[20][12] = kernel[0][0] ~^ image[20][12] + kernel[0][1] ~^ image[20][13] + kernel[0][2] ~^ image[20][14] + kernel[0][3] ~^ image[20][15] + kernel[0][4] ~^ image[20][16] + kernel[1][0] ~^ image[21][12] + kernel[1][1] ~^ image[21][13] + kernel[1][2] ~^ image[21][14] + kernel[1][3] ~^ image[21][15] + kernel[1][4] ~^ image[21][16] + kernel[2][0] ~^ image[22][12] + kernel[2][1] ~^ image[22][13] + kernel[2][2] ~^ image[22][14] + kernel[2][3] ~^ image[22][15] + kernel[2][4] ~^ image[22][16] + kernel[3][0] ~^ image[23][12] + kernel[3][1] ~^ image[23][13] + kernel[3][2] ~^ image[23][14] + kernel[3][3] ~^ image[23][15] + kernel[3][4] ~^ image[23][16] + kernel[4][0] ~^ image[24][12] + kernel[4][1] ~^ image[24][13] + kernel[4][2] ~^ image[24][14] + kernel[4][3] ~^ image[24][15] + kernel[4][4] ~^ image[24][16];
assign xor_sum[20][13] = kernel[0][0] ~^ image[20][13] + kernel[0][1] ~^ image[20][14] + kernel[0][2] ~^ image[20][15] + kernel[0][3] ~^ image[20][16] + kernel[0][4] ~^ image[20][17] + kernel[1][0] ~^ image[21][13] + kernel[1][1] ~^ image[21][14] + kernel[1][2] ~^ image[21][15] + kernel[1][3] ~^ image[21][16] + kernel[1][4] ~^ image[21][17] + kernel[2][0] ~^ image[22][13] + kernel[2][1] ~^ image[22][14] + kernel[2][2] ~^ image[22][15] + kernel[2][3] ~^ image[22][16] + kernel[2][4] ~^ image[22][17] + kernel[3][0] ~^ image[23][13] + kernel[3][1] ~^ image[23][14] + kernel[3][2] ~^ image[23][15] + kernel[3][3] ~^ image[23][16] + kernel[3][4] ~^ image[23][17] + kernel[4][0] ~^ image[24][13] + kernel[4][1] ~^ image[24][14] + kernel[4][2] ~^ image[24][15] + kernel[4][3] ~^ image[24][16] + kernel[4][4] ~^ image[24][17];
assign xor_sum[20][14] = kernel[0][0] ~^ image[20][14] + kernel[0][1] ~^ image[20][15] + kernel[0][2] ~^ image[20][16] + kernel[0][3] ~^ image[20][17] + kernel[0][4] ~^ image[20][18] + kernel[1][0] ~^ image[21][14] + kernel[1][1] ~^ image[21][15] + kernel[1][2] ~^ image[21][16] + kernel[1][3] ~^ image[21][17] + kernel[1][4] ~^ image[21][18] + kernel[2][0] ~^ image[22][14] + kernel[2][1] ~^ image[22][15] + kernel[2][2] ~^ image[22][16] + kernel[2][3] ~^ image[22][17] + kernel[2][4] ~^ image[22][18] + kernel[3][0] ~^ image[23][14] + kernel[3][1] ~^ image[23][15] + kernel[3][2] ~^ image[23][16] + kernel[3][3] ~^ image[23][17] + kernel[3][4] ~^ image[23][18] + kernel[4][0] ~^ image[24][14] + kernel[4][1] ~^ image[24][15] + kernel[4][2] ~^ image[24][16] + kernel[4][3] ~^ image[24][17] + kernel[4][4] ~^ image[24][18];
assign xor_sum[20][15] = kernel[0][0] ~^ image[20][15] + kernel[0][1] ~^ image[20][16] + kernel[0][2] ~^ image[20][17] + kernel[0][3] ~^ image[20][18] + kernel[0][4] ~^ image[20][19] + kernel[1][0] ~^ image[21][15] + kernel[1][1] ~^ image[21][16] + kernel[1][2] ~^ image[21][17] + kernel[1][3] ~^ image[21][18] + kernel[1][4] ~^ image[21][19] + kernel[2][0] ~^ image[22][15] + kernel[2][1] ~^ image[22][16] + kernel[2][2] ~^ image[22][17] + kernel[2][3] ~^ image[22][18] + kernel[2][4] ~^ image[22][19] + kernel[3][0] ~^ image[23][15] + kernel[3][1] ~^ image[23][16] + kernel[3][2] ~^ image[23][17] + kernel[3][3] ~^ image[23][18] + kernel[3][4] ~^ image[23][19] + kernel[4][0] ~^ image[24][15] + kernel[4][1] ~^ image[24][16] + kernel[4][2] ~^ image[24][17] + kernel[4][3] ~^ image[24][18] + kernel[4][4] ~^ image[24][19];
assign xor_sum[20][16] = kernel[0][0] ~^ image[20][16] + kernel[0][1] ~^ image[20][17] + kernel[0][2] ~^ image[20][18] + kernel[0][3] ~^ image[20][19] + kernel[0][4] ~^ image[20][20] + kernel[1][0] ~^ image[21][16] + kernel[1][1] ~^ image[21][17] + kernel[1][2] ~^ image[21][18] + kernel[1][3] ~^ image[21][19] + kernel[1][4] ~^ image[21][20] + kernel[2][0] ~^ image[22][16] + kernel[2][1] ~^ image[22][17] + kernel[2][2] ~^ image[22][18] + kernel[2][3] ~^ image[22][19] + kernel[2][4] ~^ image[22][20] + kernel[3][0] ~^ image[23][16] + kernel[3][1] ~^ image[23][17] + kernel[3][2] ~^ image[23][18] + kernel[3][3] ~^ image[23][19] + kernel[3][4] ~^ image[23][20] + kernel[4][0] ~^ image[24][16] + kernel[4][1] ~^ image[24][17] + kernel[4][2] ~^ image[24][18] + kernel[4][3] ~^ image[24][19] + kernel[4][4] ~^ image[24][20];
assign xor_sum[20][17] = kernel[0][0] ~^ image[20][17] + kernel[0][1] ~^ image[20][18] + kernel[0][2] ~^ image[20][19] + kernel[0][3] ~^ image[20][20] + kernel[0][4] ~^ image[20][21] + kernel[1][0] ~^ image[21][17] + kernel[1][1] ~^ image[21][18] + kernel[1][2] ~^ image[21][19] + kernel[1][3] ~^ image[21][20] + kernel[1][4] ~^ image[21][21] + kernel[2][0] ~^ image[22][17] + kernel[2][1] ~^ image[22][18] + kernel[2][2] ~^ image[22][19] + kernel[2][3] ~^ image[22][20] + kernel[2][4] ~^ image[22][21] + kernel[3][0] ~^ image[23][17] + kernel[3][1] ~^ image[23][18] + kernel[3][2] ~^ image[23][19] + kernel[3][3] ~^ image[23][20] + kernel[3][4] ~^ image[23][21] + kernel[4][0] ~^ image[24][17] + kernel[4][1] ~^ image[24][18] + kernel[4][2] ~^ image[24][19] + kernel[4][3] ~^ image[24][20] + kernel[4][4] ~^ image[24][21];
assign xor_sum[20][18] = kernel[0][0] ~^ image[20][18] + kernel[0][1] ~^ image[20][19] + kernel[0][2] ~^ image[20][20] + kernel[0][3] ~^ image[20][21] + kernel[0][4] ~^ image[20][22] + kernel[1][0] ~^ image[21][18] + kernel[1][1] ~^ image[21][19] + kernel[1][2] ~^ image[21][20] + kernel[1][3] ~^ image[21][21] + kernel[1][4] ~^ image[21][22] + kernel[2][0] ~^ image[22][18] + kernel[2][1] ~^ image[22][19] + kernel[2][2] ~^ image[22][20] + kernel[2][3] ~^ image[22][21] + kernel[2][4] ~^ image[22][22] + kernel[3][0] ~^ image[23][18] + kernel[3][1] ~^ image[23][19] + kernel[3][2] ~^ image[23][20] + kernel[3][3] ~^ image[23][21] + kernel[3][4] ~^ image[23][22] + kernel[4][0] ~^ image[24][18] + kernel[4][1] ~^ image[24][19] + kernel[4][2] ~^ image[24][20] + kernel[4][3] ~^ image[24][21] + kernel[4][4] ~^ image[24][22];
assign xor_sum[20][19] = kernel[0][0] ~^ image[20][19] + kernel[0][1] ~^ image[20][20] + kernel[0][2] ~^ image[20][21] + kernel[0][3] ~^ image[20][22] + kernel[0][4] ~^ image[20][23] + kernel[1][0] ~^ image[21][19] + kernel[1][1] ~^ image[21][20] + kernel[1][2] ~^ image[21][21] + kernel[1][3] ~^ image[21][22] + kernel[1][4] ~^ image[21][23] + kernel[2][0] ~^ image[22][19] + kernel[2][1] ~^ image[22][20] + kernel[2][2] ~^ image[22][21] + kernel[2][3] ~^ image[22][22] + kernel[2][4] ~^ image[22][23] + kernel[3][0] ~^ image[23][19] + kernel[3][1] ~^ image[23][20] + kernel[3][2] ~^ image[23][21] + kernel[3][3] ~^ image[23][22] + kernel[3][4] ~^ image[23][23] + kernel[4][0] ~^ image[24][19] + kernel[4][1] ~^ image[24][20] + kernel[4][2] ~^ image[24][21] + kernel[4][3] ~^ image[24][22] + kernel[4][4] ~^ image[24][23];
assign xor_sum[20][20] = kernel[0][0] ~^ image[20][20] + kernel[0][1] ~^ image[20][21] + kernel[0][2] ~^ image[20][22] + kernel[0][3] ~^ image[20][23] + kernel[0][4] ~^ image[20][24] + kernel[1][0] ~^ image[21][20] + kernel[1][1] ~^ image[21][21] + kernel[1][2] ~^ image[21][22] + kernel[1][3] ~^ image[21][23] + kernel[1][4] ~^ image[21][24] + kernel[2][0] ~^ image[22][20] + kernel[2][1] ~^ image[22][21] + kernel[2][2] ~^ image[22][22] + kernel[2][3] ~^ image[22][23] + kernel[2][4] ~^ image[22][24] + kernel[3][0] ~^ image[23][20] + kernel[3][1] ~^ image[23][21] + kernel[3][2] ~^ image[23][22] + kernel[3][3] ~^ image[23][23] + kernel[3][4] ~^ image[23][24] + kernel[4][0] ~^ image[24][20] + kernel[4][1] ~^ image[24][21] + kernel[4][2] ~^ image[24][22] + kernel[4][3] ~^ image[24][23] + kernel[4][4] ~^ image[24][24];
assign xor_sum[20][21] = kernel[0][0] ~^ image[20][21] + kernel[0][1] ~^ image[20][22] + kernel[0][2] ~^ image[20][23] + kernel[0][3] ~^ image[20][24] + kernel[0][4] ~^ image[20][25] + kernel[1][0] ~^ image[21][21] + kernel[1][1] ~^ image[21][22] + kernel[1][2] ~^ image[21][23] + kernel[1][3] ~^ image[21][24] + kernel[1][4] ~^ image[21][25] + kernel[2][0] ~^ image[22][21] + kernel[2][1] ~^ image[22][22] + kernel[2][2] ~^ image[22][23] + kernel[2][3] ~^ image[22][24] + kernel[2][4] ~^ image[22][25] + kernel[3][0] ~^ image[23][21] + kernel[3][1] ~^ image[23][22] + kernel[3][2] ~^ image[23][23] + kernel[3][3] ~^ image[23][24] + kernel[3][4] ~^ image[23][25] + kernel[4][0] ~^ image[24][21] + kernel[4][1] ~^ image[24][22] + kernel[4][2] ~^ image[24][23] + kernel[4][3] ~^ image[24][24] + kernel[4][4] ~^ image[24][25];
assign xor_sum[20][22] = kernel[0][0] ~^ image[20][22] + kernel[0][1] ~^ image[20][23] + kernel[0][2] ~^ image[20][24] + kernel[0][3] ~^ image[20][25] + kernel[0][4] ~^ image[20][26] + kernel[1][0] ~^ image[21][22] + kernel[1][1] ~^ image[21][23] + kernel[1][2] ~^ image[21][24] + kernel[1][3] ~^ image[21][25] + kernel[1][4] ~^ image[21][26] + kernel[2][0] ~^ image[22][22] + kernel[2][1] ~^ image[22][23] + kernel[2][2] ~^ image[22][24] + kernel[2][3] ~^ image[22][25] + kernel[2][4] ~^ image[22][26] + kernel[3][0] ~^ image[23][22] + kernel[3][1] ~^ image[23][23] + kernel[3][2] ~^ image[23][24] + kernel[3][3] ~^ image[23][25] + kernel[3][4] ~^ image[23][26] + kernel[4][0] ~^ image[24][22] + kernel[4][1] ~^ image[24][23] + kernel[4][2] ~^ image[24][24] + kernel[4][3] ~^ image[24][25] + kernel[4][4] ~^ image[24][26];
assign xor_sum[20][23] = kernel[0][0] ~^ image[20][23] + kernel[0][1] ~^ image[20][24] + kernel[0][2] ~^ image[20][25] + kernel[0][3] ~^ image[20][26] + kernel[0][4] ~^ image[20][27] + kernel[1][0] ~^ image[21][23] + kernel[1][1] ~^ image[21][24] + kernel[1][2] ~^ image[21][25] + kernel[1][3] ~^ image[21][26] + kernel[1][4] ~^ image[21][27] + kernel[2][0] ~^ image[22][23] + kernel[2][1] ~^ image[22][24] + kernel[2][2] ~^ image[22][25] + kernel[2][3] ~^ image[22][26] + kernel[2][4] ~^ image[22][27] + kernel[3][0] ~^ image[23][23] + kernel[3][1] ~^ image[23][24] + kernel[3][2] ~^ image[23][25] + kernel[3][3] ~^ image[23][26] + kernel[3][4] ~^ image[23][27] + kernel[4][0] ~^ image[24][23] + kernel[4][1] ~^ image[24][24] + kernel[4][2] ~^ image[24][25] + kernel[4][3] ~^ image[24][26] + kernel[4][4] ~^ image[24][27];
assign xor_sum[21][0] = kernel[0][0] ~^ image[21][0] + kernel[0][1] ~^ image[21][1] + kernel[0][2] ~^ image[21][2] + kernel[0][3] ~^ image[21][3] + kernel[0][4] ~^ image[21][4] + kernel[1][0] ~^ image[22][0] + kernel[1][1] ~^ image[22][1] + kernel[1][2] ~^ image[22][2] + kernel[1][3] ~^ image[22][3] + kernel[1][4] ~^ image[22][4] + kernel[2][0] ~^ image[23][0] + kernel[2][1] ~^ image[23][1] + kernel[2][2] ~^ image[23][2] + kernel[2][3] ~^ image[23][3] + kernel[2][4] ~^ image[23][4] + kernel[3][0] ~^ image[24][0] + kernel[3][1] ~^ image[24][1] + kernel[3][2] ~^ image[24][2] + kernel[3][3] ~^ image[24][3] + kernel[3][4] ~^ image[24][4] + kernel[4][0] ~^ image[25][0] + kernel[4][1] ~^ image[25][1] + kernel[4][2] ~^ image[25][2] + kernel[4][3] ~^ image[25][3] + kernel[4][4] ~^ image[25][4];
assign xor_sum[21][1] = kernel[0][0] ~^ image[21][1] + kernel[0][1] ~^ image[21][2] + kernel[0][2] ~^ image[21][3] + kernel[0][3] ~^ image[21][4] + kernel[0][4] ~^ image[21][5] + kernel[1][0] ~^ image[22][1] + kernel[1][1] ~^ image[22][2] + kernel[1][2] ~^ image[22][3] + kernel[1][3] ~^ image[22][4] + kernel[1][4] ~^ image[22][5] + kernel[2][0] ~^ image[23][1] + kernel[2][1] ~^ image[23][2] + kernel[2][2] ~^ image[23][3] + kernel[2][3] ~^ image[23][4] + kernel[2][4] ~^ image[23][5] + kernel[3][0] ~^ image[24][1] + kernel[3][1] ~^ image[24][2] + kernel[3][2] ~^ image[24][3] + kernel[3][3] ~^ image[24][4] + kernel[3][4] ~^ image[24][5] + kernel[4][0] ~^ image[25][1] + kernel[4][1] ~^ image[25][2] + kernel[4][2] ~^ image[25][3] + kernel[4][3] ~^ image[25][4] + kernel[4][4] ~^ image[25][5];
assign xor_sum[21][2] = kernel[0][0] ~^ image[21][2] + kernel[0][1] ~^ image[21][3] + kernel[0][2] ~^ image[21][4] + kernel[0][3] ~^ image[21][5] + kernel[0][4] ~^ image[21][6] + kernel[1][0] ~^ image[22][2] + kernel[1][1] ~^ image[22][3] + kernel[1][2] ~^ image[22][4] + kernel[1][3] ~^ image[22][5] + kernel[1][4] ~^ image[22][6] + kernel[2][0] ~^ image[23][2] + kernel[2][1] ~^ image[23][3] + kernel[2][2] ~^ image[23][4] + kernel[2][3] ~^ image[23][5] + kernel[2][4] ~^ image[23][6] + kernel[3][0] ~^ image[24][2] + kernel[3][1] ~^ image[24][3] + kernel[3][2] ~^ image[24][4] + kernel[3][3] ~^ image[24][5] + kernel[3][4] ~^ image[24][6] + kernel[4][0] ~^ image[25][2] + kernel[4][1] ~^ image[25][3] + kernel[4][2] ~^ image[25][4] + kernel[4][3] ~^ image[25][5] + kernel[4][4] ~^ image[25][6];
assign xor_sum[21][3] = kernel[0][0] ~^ image[21][3] + kernel[0][1] ~^ image[21][4] + kernel[0][2] ~^ image[21][5] + kernel[0][3] ~^ image[21][6] + kernel[0][4] ~^ image[21][7] + kernel[1][0] ~^ image[22][3] + kernel[1][1] ~^ image[22][4] + kernel[1][2] ~^ image[22][5] + kernel[1][3] ~^ image[22][6] + kernel[1][4] ~^ image[22][7] + kernel[2][0] ~^ image[23][3] + kernel[2][1] ~^ image[23][4] + kernel[2][2] ~^ image[23][5] + kernel[2][3] ~^ image[23][6] + kernel[2][4] ~^ image[23][7] + kernel[3][0] ~^ image[24][3] + kernel[3][1] ~^ image[24][4] + kernel[3][2] ~^ image[24][5] + kernel[3][3] ~^ image[24][6] + kernel[3][4] ~^ image[24][7] + kernel[4][0] ~^ image[25][3] + kernel[4][1] ~^ image[25][4] + kernel[4][2] ~^ image[25][5] + kernel[4][3] ~^ image[25][6] + kernel[4][4] ~^ image[25][7];
assign xor_sum[21][4] = kernel[0][0] ~^ image[21][4] + kernel[0][1] ~^ image[21][5] + kernel[0][2] ~^ image[21][6] + kernel[0][3] ~^ image[21][7] + kernel[0][4] ~^ image[21][8] + kernel[1][0] ~^ image[22][4] + kernel[1][1] ~^ image[22][5] + kernel[1][2] ~^ image[22][6] + kernel[1][3] ~^ image[22][7] + kernel[1][4] ~^ image[22][8] + kernel[2][0] ~^ image[23][4] + kernel[2][1] ~^ image[23][5] + kernel[2][2] ~^ image[23][6] + kernel[2][3] ~^ image[23][7] + kernel[2][4] ~^ image[23][8] + kernel[3][0] ~^ image[24][4] + kernel[3][1] ~^ image[24][5] + kernel[3][2] ~^ image[24][6] + kernel[3][3] ~^ image[24][7] + kernel[3][4] ~^ image[24][8] + kernel[4][0] ~^ image[25][4] + kernel[4][1] ~^ image[25][5] + kernel[4][2] ~^ image[25][6] + kernel[4][3] ~^ image[25][7] + kernel[4][4] ~^ image[25][8];
assign xor_sum[21][5] = kernel[0][0] ~^ image[21][5] + kernel[0][1] ~^ image[21][6] + kernel[0][2] ~^ image[21][7] + kernel[0][3] ~^ image[21][8] + kernel[0][4] ~^ image[21][9] + kernel[1][0] ~^ image[22][5] + kernel[1][1] ~^ image[22][6] + kernel[1][2] ~^ image[22][7] + kernel[1][3] ~^ image[22][8] + kernel[1][4] ~^ image[22][9] + kernel[2][0] ~^ image[23][5] + kernel[2][1] ~^ image[23][6] + kernel[2][2] ~^ image[23][7] + kernel[2][3] ~^ image[23][8] + kernel[2][4] ~^ image[23][9] + kernel[3][0] ~^ image[24][5] + kernel[3][1] ~^ image[24][6] + kernel[3][2] ~^ image[24][7] + kernel[3][3] ~^ image[24][8] + kernel[3][4] ~^ image[24][9] + kernel[4][0] ~^ image[25][5] + kernel[4][1] ~^ image[25][6] + kernel[4][2] ~^ image[25][7] + kernel[4][3] ~^ image[25][8] + kernel[4][4] ~^ image[25][9];
assign xor_sum[21][6] = kernel[0][0] ~^ image[21][6] + kernel[0][1] ~^ image[21][7] + kernel[0][2] ~^ image[21][8] + kernel[0][3] ~^ image[21][9] + kernel[0][4] ~^ image[21][10] + kernel[1][0] ~^ image[22][6] + kernel[1][1] ~^ image[22][7] + kernel[1][2] ~^ image[22][8] + kernel[1][3] ~^ image[22][9] + kernel[1][4] ~^ image[22][10] + kernel[2][0] ~^ image[23][6] + kernel[2][1] ~^ image[23][7] + kernel[2][2] ~^ image[23][8] + kernel[2][3] ~^ image[23][9] + kernel[2][4] ~^ image[23][10] + kernel[3][0] ~^ image[24][6] + kernel[3][1] ~^ image[24][7] + kernel[3][2] ~^ image[24][8] + kernel[3][3] ~^ image[24][9] + kernel[3][4] ~^ image[24][10] + kernel[4][0] ~^ image[25][6] + kernel[4][1] ~^ image[25][7] + kernel[4][2] ~^ image[25][8] + kernel[4][3] ~^ image[25][9] + kernel[4][4] ~^ image[25][10];
assign xor_sum[21][7] = kernel[0][0] ~^ image[21][7] + kernel[0][1] ~^ image[21][8] + kernel[0][2] ~^ image[21][9] + kernel[0][3] ~^ image[21][10] + kernel[0][4] ~^ image[21][11] + kernel[1][0] ~^ image[22][7] + kernel[1][1] ~^ image[22][8] + kernel[1][2] ~^ image[22][9] + kernel[1][3] ~^ image[22][10] + kernel[1][4] ~^ image[22][11] + kernel[2][0] ~^ image[23][7] + kernel[2][1] ~^ image[23][8] + kernel[2][2] ~^ image[23][9] + kernel[2][3] ~^ image[23][10] + kernel[2][4] ~^ image[23][11] + kernel[3][0] ~^ image[24][7] + kernel[3][1] ~^ image[24][8] + kernel[3][2] ~^ image[24][9] + kernel[3][3] ~^ image[24][10] + kernel[3][4] ~^ image[24][11] + kernel[4][0] ~^ image[25][7] + kernel[4][1] ~^ image[25][8] + kernel[4][2] ~^ image[25][9] + kernel[4][3] ~^ image[25][10] + kernel[4][4] ~^ image[25][11];
assign xor_sum[21][8] = kernel[0][0] ~^ image[21][8] + kernel[0][1] ~^ image[21][9] + kernel[0][2] ~^ image[21][10] + kernel[0][3] ~^ image[21][11] + kernel[0][4] ~^ image[21][12] + kernel[1][0] ~^ image[22][8] + kernel[1][1] ~^ image[22][9] + kernel[1][2] ~^ image[22][10] + kernel[1][3] ~^ image[22][11] + kernel[1][4] ~^ image[22][12] + kernel[2][0] ~^ image[23][8] + kernel[2][1] ~^ image[23][9] + kernel[2][2] ~^ image[23][10] + kernel[2][3] ~^ image[23][11] + kernel[2][4] ~^ image[23][12] + kernel[3][0] ~^ image[24][8] + kernel[3][1] ~^ image[24][9] + kernel[3][2] ~^ image[24][10] + kernel[3][3] ~^ image[24][11] + kernel[3][4] ~^ image[24][12] + kernel[4][0] ~^ image[25][8] + kernel[4][1] ~^ image[25][9] + kernel[4][2] ~^ image[25][10] + kernel[4][3] ~^ image[25][11] + kernel[4][4] ~^ image[25][12];
assign xor_sum[21][9] = kernel[0][0] ~^ image[21][9] + kernel[0][1] ~^ image[21][10] + kernel[0][2] ~^ image[21][11] + kernel[0][3] ~^ image[21][12] + kernel[0][4] ~^ image[21][13] + kernel[1][0] ~^ image[22][9] + kernel[1][1] ~^ image[22][10] + kernel[1][2] ~^ image[22][11] + kernel[1][3] ~^ image[22][12] + kernel[1][4] ~^ image[22][13] + kernel[2][0] ~^ image[23][9] + kernel[2][1] ~^ image[23][10] + kernel[2][2] ~^ image[23][11] + kernel[2][3] ~^ image[23][12] + kernel[2][4] ~^ image[23][13] + kernel[3][0] ~^ image[24][9] + kernel[3][1] ~^ image[24][10] + kernel[3][2] ~^ image[24][11] + kernel[3][3] ~^ image[24][12] + kernel[3][4] ~^ image[24][13] + kernel[4][0] ~^ image[25][9] + kernel[4][1] ~^ image[25][10] + kernel[4][2] ~^ image[25][11] + kernel[4][3] ~^ image[25][12] + kernel[4][4] ~^ image[25][13];
assign xor_sum[21][10] = kernel[0][0] ~^ image[21][10] + kernel[0][1] ~^ image[21][11] + kernel[0][2] ~^ image[21][12] + kernel[0][3] ~^ image[21][13] + kernel[0][4] ~^ image[21][14] + kernel[1][0] ~^ image[22][10] + kernel[1][1] ~^ image[22][11] + kernel[1][2] ~^ image[22][12] + kernel[1][3] ~^ image[22][13] + kernel[1][4] ~^ image[22][14] + kernel[2][0] ~^ image[23][10] + kernel[2][1] ~^ image[23][11] + kernel[2][2] ~^ image[23][12] + kernel[2][3] ~^ image[23][13] + kernel[2][4] ~^ image[23][14] + kernel[3][0] ~^ image[24][10] + kernel[3][1] ~^ image[24][11] + kernel[3][2] ~^ image[24][12] + kernel[3][3] ~^ image[24][13] + kernel[3][4] ~^ image[24][14] + kernel[4][0] ~^ image[25][10] + kernel[4][1] ~^ image[25][11] + kernel[4][2] ~^ image[25][12] + kernel[4][3] ~^ image[25][13] + kernel[4][4] ~^ image[25][14];
assign xor_sum[21][11] = kernel[0][0] ~^ image[21][11] + kernel[0][1] ~^ image[21][12] + kernel[0][2] ~^ image[21][13] + kernel[0][3] ~^ image[21][14] + kernel[0][4] ~^ image[21][15] + kernel[1][0] ~^ image[22][11] + kernel[1][1] ~^ image[22][12] + kernel[1][2] ~^ image[22][13] + kernel[1][3] ~^ image[22][14] + kernel[1][4] ~^ image[22][15] + kernel[2][0] ~^ image[23][11] + kernel[2][1] ~^ image[23][12] + kernel[2][2] ~^ image[23][13] + kernel[2][3] ~^ image[23][14] + kernel[2][4] ~^ image[23][15] + kernel[3][0] ~^ image[24][11] + kernel[3][1] ~^ image[24][12] + kernel[3][2] ~^ image[24][13] + kernel[3][3] ~^ image[24][14] + kernel[3][4] ~^ image[24][15] + kernel[4][0] ~^ image[25][11] + kernel[4][1] ~^ image[25][12] + kernel[4][2] ~^ image[25][13] + kernel[4][3] ~^ image[25][14] + kernel[4][4] ~^ image[25][15];
assign xor_sum[21][12] = kernel[0][0] ~^ image[21][12] + kernel[0][1] ~^ image[21][13] + kernel[0][2] ~^ image[21][14] + kernel[0][3] ~^ image[21][15] + kernel[0][4] ~^ image[21][16] + kernel[1][0] ~^ image[22][12] + kernel[1][1] ~^ image[22][13] + kernel[1][2] ~^ image[22][14] + kernel[1][3] ~^ image[22][15] + kernel[1][4] ~^ image[22][16] + kernel[2][0] ~^ image[23][12] + kernel[2][1] ~^ image[23][13] + kernel[2][2] ~^ image[23][14] + kernel[2][3] ~^ image[23][15] + kernel[2][4] ~^ image[23][16] + kernel[3][0] ~^ image[24][12] + kernel[3][1] ~^ image[24][13] + kernel[3][2] ~^ image[24][14] + kernel[3][3] ~^ image[24][15] + kernel[3][4] ~^ image[24][16] + kernel[4][0] ~^ image[25][12] + kernel[4][1] ~^ image[25][13] + kernel[4][2] ~^ image[25][14] + kernel[4][3] ~^ image[25][15] + kernel[4][4] ~^ image[25][16];
assign xor_sum[21][13] = kernel[0][0] ~^ image[21][13] + kernel[0][1] ~^ image[21][14] + kernel[0][2] ~^ image[21][15] + kernel[0][3] ~^ image[21][16] + kernel[0][4] ~^ image[21][17] + kernel[1][0] ~^ image[22][13] + kernel[1][1] ~^ image[22][14] + kernel[1][2] ~^ image[22][15] + kernel[1][3] ~^ image[22][16] + kernel[1][4] ~^ image[22][17] + kernel[2][0] ~^ image[23][13] + kernel[2][1] ~^ image[23][14] + kernel[2][2] ~^ image[23][15] + kernel[2][3] ~^ image[23][16] + kernel[2][4] ~^ image[23][17] + kernel[3][0] ~^ image[24][13] + kernel[3][1] ~^ image[24][14] + kernel[3][2] ~^ image[24][15] + kernel[3][3] ~^ image[24][16] + kernel[3][4] ~^ image[24][17] + kernel[4][0] ~^ image[25][13] + kernel[4][1] ~^ image[25][14] + kernel[4][2] ~^ image[25][15] + kernel[4][3] ~^ image[25][16] + kernel[4][4] ~^ image[25][17];
assign xor_sum[21][14] = kernel[0][0] ~^ image[21][14] + kernel[0][1] ~^ image[21][15] + kernel[0][2] ~^ image[21][16] + kernel[0][3] ~^ image[21][17] + kernel[0][4] ~^ image[21][18] + kernel[1][0] ~^ image[22][14] + kernel[1][1] ~^ image[22][15] + kernel[1][2] ~^ image[22][16] + kernel[1][3] ~^ image[22][17] + kernel[1][4] ~^ image[22][18] + kernel[2][0] ~^ image[23][14] + kernel[2][1] ~^ image[23][15] + kernel[2][2] ~^ image[23][16] + kernel[2][3] ~^ image[23][17] + kernel[2][4] ~^ image[23][18] + kernel[3][0] ~^ image[24][14] + kernel[3][1] ~^ image[24][15] + kernel[3][2] ~^ image[24][16] + kernel[3][3] ~^ image[24][17] + kernel[3][4] ~^ image[24][18] + kernel[4][0] ~^ image[25][14] + kernel[4][1] ~^ image[25][15] + kernel[4][2] ~^ image[25][16] + kernel[4][3] ~^ image[25][17] + kernel[4][4] ~^ image[25][18];
assign xor_sum[21][15] = kernel[0][0] ~^ image[21][15] + kernel[0][1] ~^ image[21][16] + kernel[0][2] ~^ image[21][17] + kernel[0][3] ~^ image[21][18] + kernel[0][4] ~^ image[21][19] + kernel[1][0] ~^ image[22][15] + kernel[1][1] ~^ image[22][16] + kernel[1][2] ~^ image[22][17] + kernel[1][3] ~^ image[22][18] + kernel[1][4] ~^ image[22][19] + kernel[2][0] ~^ image[23][15] + kernel[2][1] ~^ image[23][16] + kernel[2][2] ~^ image[23][17] + kernel[2][3] ~^ image[23][18] + kernel[2][4] ~^ image[23][19] + kernel[3][0] ~^ image[24][15] + kernel[3][1] ~^ image[24][16] + kernel[3][2] ~^ image[24][17] + kernel[3][3] ~^ image[24][18] + kernel[3][4] ~^ image[24][19] + kernel[4][0] ~^ image[25][15] + kernel[4][1] ~^ image[25][16] + kernel[4][2] ~^ image[25][17] + kernel[4][3] ~^ image[25][18] + kernel[4][4] ~^ image[25][19];
assign xor_sum[21][16] = kernel[0][0] ~^ image[21][16] + kernel[0][1] ~^ image[21][17] + kernel[0][2] ~^ image[21][18] + kernel[0][3] ~^ image[21][19] + kernel[0][4] ~^ image[21][20] + kernel[1][0] ~^ image[22][16] + kernel[1][1] ~^ image[22][17] + kernel[1][2] ~^ image[22][18] + kernel[1][3] ~^ image[22][19] + kernel[1][4] ~^ image[22][20] + kernel[2][0] ~^ image[23][16] + kernel[2][1] ~^ image[23][17] + kernel[2][2] ~^ image[23][18] + kernel[2][3] ~^ image[23][19] + kernel[2][4] ~^ image[23][20] + kernel[3][0] ~^ image[24][16] + kernel[3][1] ~^ image[24][17] + kernel[3][2] ~^ image[24][18] + kernel[3][3] ~^ image[24][19] + kernel[3][4] ~^ image[24][20] + kernel[4][0] ~^ image[25][16] + kernel[4][1] ~^ image[25][17] + kernel[4][2] ~^ image[25][18] + kernel[4][3] ~^ image[25][19] + kernel[4][4] ~^ image[25][20];
assign xor_sum[21][17] = kernel[0][0] ~^ image[21][17] + kernel[0][1] ~^ image[21][18] + kernel[0][2] ~^ image[21][19] + kernel[0][3] ~^ image[21][20] + kernel[0][4] ~^ image[21][21] + kernel[1][0] ~^ image[22][17] + kernel[1][1] ~^ image[22][18] + kernel[1][2] ~^ image[22][19] + kernel[1][3] ~^ image[22][20] + kernel[1][4] ~^ image[22][21] + kernel[2][0] ~^ image[23][17] + kernel[2][1] ~^ image[23][18] + kernel[2][2] ~^ image[23][19] + kernel[2][3] ~^ image[23][20] + kernel[2][4] ~^ image[23][21] + kernel[3][0] ~^ image[24][17] + kernel[3][1] ~^ image[24][18] + kernel[3][2] ~^ image[24][19] + kernel[3][3] ~^ image[24][20] + kernel[3][4] ~^ image[24][21] + kernel[4][0] ~^ image[25][17] + kernel[4][1] ~^ image[25][18] + kernel[4][2] ~^ image[25][19] + kernel[4][3] ~^ image[25][20] + kernel[4][4] ~^ image[25][21];
assign xor_sum[21][18] = kernel[0][0] ~^ image[21][18] + kernel[0][1] ~^ image[21][19] + kernel[0][2] ~^ image[21][20] + kernel[0][3] ~^ image[21][21] + kernel[0][4] ~^ image[21][22] + kernel[1][0] ~^ image[22][18] + kernel[1][1] ~^ image[22][19] + kernel[1][2] ~^ image[22][20] + kernel[1][3] ~^ image[22][21] + kernel[1][4] ~^ image[22][22] + kernel[2][0] ~^ image[23][18] + kernel[2][1] ~^ image[23][19] + kernel[2][2] ~^ image[23][20] + kernel[2][3] ~^ image[23][21] + kernel[2][4] ~^ image[23][22] + kernel[3][0] ~^ image[24][18] + kernel[3][1] ~^ image[24][19] + kernel[3][2] ~^ image[24][20] + kernel[3][3] ~^ image[24][21] + kernel[3][4] ~^ image[24][22] + kernel[4][0] ~^ image[25][18] + kernel[4][1] ~^ image[25][19] + kernel[4][2] ~^ image[25][20] + kernel[4][3] ~^ image[25][21] + kernel[4][4] ~^ image[25][22];
assign xor_sum[21][19] = kernel[0][0] ~^ image[21][19] + kernel[0][1] ~^ image[21][20] + kernel[0][2] ~^ image[21][21] + kernel[0][3] ~^ image[21][22] + kernel[0][4] ~^ image[21][23] + kernel[1][0] ~^ image[22][19] + kernel[1][1] ~^ image[22][20] + kernel[1][2] ~^ image[22][21] + kernel[1][3] ~^ image[22][22] + kernel[1][4] ~^ image[22][23] + kernel[2][0] ~^ image[23][19] + kernel[2][1] ~^ image[23][20] + kernel[2][2] ~^ image[23][21] + kernel[2][3] ~^ image[23][22] + kernel[2][4] ~^ image[23][23] + kernel[3][0] ~^ image[24][19] + kernel[3][1] ~^ image[24][20] + kernel[3][2] ~^ image[24][21] + kernel[3][3] ~^ image[24][22] + kernel[3][4] ~^ image[24][23] + kernel[4][0] ~^ image[25][19] + kernel[4][1] ~^ image[25][20] + kernel[4][2] ~^ image[25][21] + kernel[4][3] ~^ image[25][22] + kernel[4][4] ~^ image[25][23];
assign xor_sum[21][20] = kernel[0][0] ~^ image[21][20] + kernel[0][1] ~^ image[21][21] + kernel[0][2] ~^ image[21][22] + kernel[0][3] ~^ image[21][23] + kernel[0][4] ~^ image[21][24] + kernel[1][0] ~^ image[22][20] + kernel[1][1] ~^ image[22][21] + kernel[1][2] ~^ image[22][22] + kernel[1][3] ~^ image[22][23] + kernel[1][4] ~^ image[22][24] + kernel[2][0] ~^ image[23][20] + kernel[2][1] ~^ image[23][21] + kernel[2][2] ~^ image[23][22] + kernel[2][3] ~^ image[23][23] + kernel[2][4] ~^ image[23][24] + kernel[3][0] ~^ image[24][20] + kernel[3][1] ~^ image[24][21] + kernel[3][2] ~^ image[24][22] + kernel[3][3] ~^ image[24][23] + kernel[3][4] ~^ image[24][24] + kernel[4][0] ~^ image[25][20] + kernel[4][1] ~^ image[25][21] + kernel[4][2] ~^ image[25][22] + kernel[4][3] ~^ image[25][23] + kernel[4][4] ~^ image[25][24];
assign xor_sum[21][21] = kernel[0][0] ~^ image[21][21] + kernel[0][1] ~^ image[21][22] + kernel[0][2] ~^ image[21][23] + kernel[0][3] ~^ image[21][24] + kernel[0][4] ~^ image[21][25] + kernel[1][0] ~^ image[22][21] + kernel[1][1] ~^ image[22][22] + kernel[1][2] ~^ image[22][23] + kernel[1][3] ~^ image[22][24] + kernel[1][4] ~^ image[22][25] + kernel[2][0] ~^ image[23][21] + kernel[2][1] ~^ image[23][22] + kernel[2][2] ~^ image[23][23] + kernel[2][3] ~^ image[23][24] + kernel[2][4] ~^ image[23][25] + kernel[3][0] ~^ image[24][21] + kernel[3][1] ~^ image[24][22] + kernel[3][2] ~^ image[24][23] + kernel[3][3] ~^ image[24][24] + kernel[3][4] ~^ image[24][25] + kernel[4][0] ~^ image[25][21] + kernel[4][1] ~^ image[25][22] + kernel[4][2] ~^ image[25][23] + kernel[4][3] ~^ image[25][24] + kernel[4][4] ~^ image[25][25];
assign xor_sum[21][22] = kernel[0][0] ~^ image[21][22] + kernel[0][1] ~^ image[21][23] + kernel[0][2] ~^ image[21][24] + kernel[0][3] ~^ image[21][25] + kernel[0][4] ~^ image[21][26] + kernel[1][0] ~^ image[22][22] + kernel[1][1] ~^ image[22][23] + kernel[1][2] ~^ image[22][24] + kernel[1][3] ~^ image[22][25] + kernel[1][4] ~^ image[22][26] + kernel[2][0] ~^ image[23][22] + kernel[2][1] ~^ image[23][23] + kernel[2][2] ~^ image[23][24] + kernel[2][3] ~^ image[23][25] + kernel[2][4] ~^ image[23][26] + kernel[3][0] ~^ image[24][22] + kernel[3][1] ~^ image[24][23] + kernel[3][2] ~^ image[24][24] + kernel[3][3] ~^ image[24][25] + kernel[3][4] ~^ image[24][26] + kernel[4][0] ~^ image[25][22] + kernel[4][1] ~^ image[25][23] + kernel[4][2] ~^ image[25][24] + kernel[4][3] ~^ image[25][25] + kernel[4][4] ~^ image[25][26];
assign xor_sum[21][23] = kernel[0][0] ~^ image[21][23] + kernel[0][1] ~^ image[21][24] + kernel[0][2] ~^ image[21][25] + kernel[0][3] ~^ image[21][26] + kernel[0][4] ~^ image[21][27] + kernel[1][0] ~^ image[22][23] + kernel[1][1] ~^ image[22][24] + kernel[1][2] ~^ image[22][25] + kernel[1][3] ~^ image[22][26] + kernel[1][4] ~^ image[22][27] + kernel[2][0] ~^ image[23][23] + kernel[2][1] ~^ image[23][24] + kernel[2][2] ~^ image[23][25] + kernel[2][3] ~^ image[23][26] + kernel[2][4] ~^ image[23][27] + kernel[3][0] ~^ image[24][23] + kernel[3][1] ~^ image[24][24] + kernel[3][2] ~^ image[24][25] + kernel[3][3] ~^ image[24][26] + kernel[3][4] ~^ image[24][27] + kernel[4][0] ~^ image[25][23] + kernel[4][1] ~^ image[25][24] + kernel[4][2] ~^ image[25][25] + kernel[4][3] ~^ image[25][26] + kernel[4][4] ~^ image[25][27];
assign xor_sum[22][0] = kernel[0][0] ~^ image[22][0] + kernel[0][1] ~^ image[22][1] + kernel[0][2] ~^ image[22][2] + kernel[0][3] ~^ image[22][3] + kernel[0][4] ~^ image[22][4] + kernel[1][0] ~^ image[23][0] + kernel[1][1] ~^ image[23][1] + kernel[1][2] ~^ image[23][2] + kernel[1][3] ~^ image[23][3] + kernel[1][4] ~^ image[23][4] + kernel[2][0] ~^ image[24][0] + kernel[2][1] ~^ image[24][1] + kernel[2][2] ~^ image[24][2] + kernel[2][3] ~^ image[24][3] + kernel[2][4] ~^ image[24][4] + kernel[3][0] ~^ image[25][0] + kernel[3][1] ~^ image[25][1] + kernel[3][2] ~^ image[25][2] + kernel[3][3] ~^ image[25][3] + kernel[3][4] ~^ image[25][4] + kernel[4][0] ~^ image[26][0] + kernel[4][1] ~^ image[26][1] + kernel[4][2] ~^ image[26][2] + kernel[4][3] ~^ image[26][3] + kernel[4][4] ~^ image[26][4];
assign xor_sum[22][1] = kernel[0][0] ~^ image[22][1] + kernel[0][1] ~^ image[22][2] + kernel[0][2] ~^ image[22][3] + kernel[0][3] ~^ image[22][4] + kernel[0][4] ~^ image[22][5] + kernel[1][0] ~^ image[23][1] + kernel[1][1] ~^ image[23][2] + kernel[1][2] ~^ image[23][3] + kernel[1][3] ~^ image[23][4] + kernel[1][4] ~^ image[23][5] + kernel[2][0] ~^ image[24][1] + kernel[2][1] ~^ image[24][2] + kernel[2][2] ~^ image[24][3] + kernel[2][3] ~^ image[24][4] + kernel[2][4] ~^ image[24][5] + kernel[3][0] ~^ image[25][1] + kernel[3][1] ~^ image[25][2] + kernel[3][2] ~^ image[25][3] + kernel[3][3] ~^ image[25][4] + kernel[3][4] ~^ image[25][5] + kernel[4][0] ~^ image[26][1] + kernel[4][1] ~^ image[26][2] + kernel[4][2] ~^ image[26][3] + kernel[4][3] ~^ image[26][4] + kernel[4][4] ~^ image[26][5];
assign xor_sum[22][2] = kernel[0][0] ~^ image[22][2] + kernel[0][1] ~^ image[22][3] + kernel[0][2] ~^ image[22][4] + kernel[0][3] ~^ image[22][5] + kernel[0][4] ~^ image[22][6] + kernel[1][0] ~^ image[23][2] + kernel[1][1] ~^ image[23][3] + kernel[1][2] ~^ image[23][4] + kernel[1][3] ~^ image[23][5] + kernel[1][4] ~^ image[23][6] + kernel[2][0] ~^ image[24][2] + kernel[2][1] ~^ image[24][3] + kernel[2][2] ~^ image[24][4] + kernel[2][3] ~^ image[24][5] + kernel[2][4] ~^ image[24][6] + kernel[3][0] ~^ image[25][2] + kernel[3][1] ~^ image[25][3] + kernel[3][2] ~^ image[25][4] + kernel[3][3] ~^ image[25][5] + kernel[3][4] ~^ image[25][6] + kernel[4][0] ~^ image[26][2] + kernel[4][1] ~^ image[26][3] + kernel[4][2] ~^ image[26][4] + kernel[4][3] ~^ image[26][5] + kernel[4][4] ~^ image[26][6];
assign xor_sum[22][3] = kernel[0][0] ~^ image[22][3] + kernel[0][1] ~^ image[22][4] + kernel[0][2] ~^ image[22][5] + kernel[0][3] ~^ image[22][6] + kernel[0][4] ~^ image[22][7] + kernel[1][0] ~^ image[23][3] + kernel[1][1] ~^ image[23][4] + kernel[1][2] ~^ image[23][5] + kernel[1][3] ~^ image[23][6] + kernel[1][4] ~^ image[23][7] + kernel[2][0] ~^ image[24][3] + kernel[2][1] ~^ image[24][4] + kernel[2][2] ~^ image[24][5] + kernel[2][3] ~^ image[24][6] + kernel[2][4] ~^ image[24][7] + kernel[3][0] ~^ image[25][3] + kernel[3][1] ~^ image[25][4] + kernel[3][2] ~^ image[25][5] + kernel[3][3] ~^ image[25][6] + kernel[3][4] ~^ image[25][7] + kernel[4][0] ~^ image[26][3] + kernel[4][1] ~^ image[26][4] + kernel[4][2] ~^ image[26][5] + kernel[4][3] ~^ image[26][6] + kernel[4][4] ~^ image[26][7];
assign xor_sum[22][4] = kernel[0][0] ~^ image[22][4] + kernel[0][1] ~^ image[22][5] + kernel[0][2] ~^ image[22][6] + kernel[0][3] ~^ image[22][7] + kernel[0][4] ~^ image[22][8] + kernel[1][0] ~^ image[23][4] + kernel[1][1] ~^ image[23][5] + kernel[1][2] ~^ image[23][6] + kernel[1][3] ~^ image[23][7] + kernel[1][4] ~^ image[23][8] + kernel[2][0] ~^ image[24][4] + kernel[2][1] ~^ image[24][5] + kernel[2][2] ~^ image[24][6] + kernel[2][3] ~^ image[24][7] + kernel[2][4] ~^ image[24][8] + kernel[3][0] ~^ image[25][4] + kernel[3][1] ~^ image[25][5] + kernel[3][2] ~^ image[25][6] + kernel[3][3] ~^ image[25][7] + kernel[3][4] ~^ image[25][8] + kernel[4][0] ~^ image[26][4] + kernel[4][1] ~^ image[26][5] + kernel[4][2] ~^ image[26][6] + kernel[4][3] ~^ image[26][7] + kernel[4][4] ~^ image[26][8];
assign xor_sum[22][5] = kernel[0][0] ~^ image[22][5] + kernel[0][1] ~^ image[22][6] + kernel[0][2] ~^ image[22][7] + kernel[0][3] ~^ image[22][8] + kernel[0][4] ~^ image[22][9] + kernel[1][0] ~^ image[23][5] + kernel[1][1] ~^ image[23][6] + kernel[1][2] ~^ image[23][7] + kernel[1][3] ~^ image[23][8] + kernel[1][4] ~^ image[23][9] + kernel[2][0] ~^ image[24][5] + kernel[2][1] ~^ image[24][6] + kernel[2][2] ~^ image[24][7] + kernel[2][3] ~^ image[24][8] + kernel[2][4] ~^ image[24][9] + kernel[3][0] ~^ image[25][5] + kernel[3][1] ~^ image[25][6] + kernel[3][2] ~^ image[25][7] + kernel[3][3] ~^ image[25][8] + kernel[3][4] ~^ image[25][9] + kernel[4][0] ~^ image[26][5] + kernel[4][1] ~^ image[26][6] + kernel[4][2] ~^ image[26][7] + kernel[4][3] ~^ image[26][8] + kernel[4][4] ~^ image[26][9];
assign xor_sum[22][6] = kernel[0][0] ~^ image[22][6] + kernel[0][1] ~^ image[22][7] + kernel[0][2] ~^ image[22][8] + kernel[0][3] ~^ image[22][9] + kernel[0][4] ~^ image[22][10] + kernel[1][0] ~^ image[23][6] + kernel[1][1] ~^ image[23][7] + kernel[1][2] ~^ image[23][8] + kernel[1][3] ~^ image[23][9] + kernel[1][4] ~^ image[23][10] + kernel[2][0] ~^ image[24][6] + kernel[2][1] ~^ image[24][7] + kernel[2][2] ~^ image[24][8] + kernel[2][3] ~^ image[24][9] + kernel[2][4] ~^ image[24][10] + kernel[3][0] ~^ image[25][6] + kernel[3][1] ~^ image[25][7] + kernel[3][2] ~^ image[25][8] + kernel[3][3] ~^ image[25][9] + kernel[3][4] ~^ image[25][10] + kernel[4][0] ~^ image[26][6] + kernel[4][1] ~^ image[26][7] + kernel[4][2] ~^ image[26][8] + kernel[4][3] ~^ image[26][9] + kernel[4][4] ~^ image[26][10];
assign xor_sum[22][7] = kernel[0][0] ~^ image[22][7] + kernel[0][1] ~^ image[22][8] + kernel[0][2] ~^ image[22][9] + kernel[0][3] ~^ image[22][10] + kernel[0][4] ~^ image[22][11] + kernel[1][0] ~^ image[23][7] + kernel[1][1] ~^ image[23][8] + kernel[1][2] ~^ image[23][9] + kernel[1][3] ~^ image[23][10] + kernel[1][4] ~^ image[23][11] + kernel[2][0] ~^ image[24][7] + kernel[2][1] ~^ image[24][8] + kernel[2][2] ~^ image[24][9] + kernel[2][3] ~^ image[24][10] + kernel[2][4] ~^ image[24][11] + kernel[3][0] ~^ image[25][7] + kernel[3][1] ~^ image[25][8] + kernel[3][2] ~^ image[25][9] + kernel[3][3] ~^ image[25][10] + kernel[3][4] ~^ image[25][11] + kernel[4][0] ~^ image[26][7] + kernel[4][1] ~^ image[26][8] + kernel[4][2] ~^ image[26][9] + kernel[4][3] ~^ image[26][10] + kernel[4][4] ~^ image[26][11];
assign xor_sum[22][8] = kernel[0][0] ~^ image[22][8] + kernel[0][1] ~^ image[22][9] + kernel[0][2] ~^ image[22][10] + kernel[0][3] ~^ image[22][11] + kernel[0][4] ~^ image[22][12] + kernel[1][0] ~^ image[23][8] + kernel[1][1] ~^ image[23][9] + kernel[1][2] ~^ image[23][10] + kernel[1][3] ~^ image[23][11] + kernel[1][4] ~^ image[23][12] + kernel[2][0] ~^ image[24][8] + kernel[2][1] ~^ image[24][9] + kernel[2][2] ~^ image[24][10] + kernel[2][3] ~^ image[24][11] + kernel[2][4] ~^ image[24][12] + kernel[3][0] ~^ image[25][8] + kernel[3][1] ~^ image[25][9] + kernel[3][2] ~^ image[25][10] + kernel[3][3] ~^ image[25][11] + kernel[3][4] ~^ image[25][12] + kernel[4][0] ~^ image[26][8] + kernel[4][1] ~^ image[26][9] + kernel[4][2] ~^ image[26][10] + kernel[4][3] ~^ image[26][11] + kernel[4][4] ~^ image[26][12];
assign xor_sum[22][9] = kernel[0][0] ~^ image[22][9] + kernel[0][1] ~^ image[22][10] + kernel[0][2] ~^ image[22][11] + kernel[0][3] ~^ image[22][12] + kernel[0][4] ~^ image[22][13] + kernel[1][0] ~^ image[23][9] + kernel[1][1] ~^ image[23][10] + kernel[1][2] ~^ image[23][11] + kernel[1][3] ~^ image[23][12] + kernel[1][4] ~^ image[23][13] + kernel[2][0] ~^ image[24][9] + kernel[2][1] ~^ image[24][10] + kernel[2][2] ~^ image[24][11] + kernel[2][3] ~^ image[24][12] + kernel[2][4] ~^ image[24][13] + kernel[3][0] ~^ image[25][9] + kernel[3][1] ~^ image[25][10] + kernel[3][2] ~^ image[25][11] + kernel[3][3] ~^ image[25][12] + kernel[3][4] ~^ image[25][13] + kernel[4][0] ~^ image[26][9] + kernel[4][1] ~^ image[26][10] + kernel[4][2] ~^ image[26][11] + kernel[4][3] ~^ image[26][12] + kernel[4][4] ~^ image[26][13];
assign xor_sum[22][10] = kernel[0][0] ~^ image[22][10] + kernel[0][1] ~^ image[22][11] + kernel[0][2] ~^ image[22][12] + kernel[0][3] ~^ image[22][13] + kernel[0][4] ~^ image[22][14] + kernel[1][0] ~^ image[23][10] + kernel[1][1] ~^ image[23][11] + kernel[1][2] ~^ image[23][12] + kernel[1][3] ~^ image[23][13] + kernel[1][4] ~^ image[23][14] + kernel[2][0] ~^ image[24][10] + kernel[2][1] ~^ image[24][11] + kernel[2][2] ~^ image[24][12] + kernel[2][3] ~^ image[24][13] + kernel[2][4] ~^ image[24][14] + kernel[3][0] ~^ image[25][10] + kernel[3][1] ~^ image[25][11] + kernel[3][2] ~^ image[25][12] + kernel[3][3] ~^ image[25][13] + kernel[3][4] ~^ image[25][14] + kernel[4][0] ~^ image[26][10] + kernel[4][1] ~^ image[26][11] + kernel[4][2] ~^ image[26][12] + kernel[4][3] ~^ image[26][13] + kernel[4][4] ~^ image[26][14];
assign xor_sum[22][11] = kernel[0][0] ~^ image[22][11] + kernel[0][1] ~^ image[22][12] + kernel[0][2] ~^ image[22][13] + kernel[0][3] ~^ image[22][14] + kernel[0][4] ~^ image[22][15] + kernel[1][0] ~^ image[23][11] + kernel[1][1] ~^ image[23][12] + kernel[1][2] ~^ image[23][13] + kernel[1][3] ~^ image[23][14] + kernel[1][4] ~^ image[23][15] + kernel[2][0] ~^ image[24][11] + kernel[2][1] ~^ image[24][12] + kernel[2][2] ~^ image[24][13] + kernel[2][3] ~^ image[24][14] + kernel[2][4] ~^ image[24][15] + kernel[3][0] ~^ image[25][11] + kernel[3][1] ~^ image[25][12] + kernel[3][2] ~^ image[25][13] + kernel[3][3] ~^ image[25][14] + kernel[3][4] ~^ image[25][15] + kernel[4][0] ~^ image[26][11] + kernel[4][1] ~^ image[26][12] + kernel[4][2] ~^ image[26][13] + kernel[4][3] ~^ image[26][14] + kernel[4][4] ~^ image[26][15];
assign xor_sum[22][12] = kernel[0][0] ~^ image[22][12] + kernel[0][1] ~^ image[22][13] + kernel[0][2] ~^ image[22][14] + kernel[0][3] ~^ image[22][15] + kernel[0][4] ~^ image[22][16] + kernel[1][0] ~^ image[23][12] + kernel[1][1] ~^ image[23][13] + kernel[1][2] ~^ image[23][14] + kernel[1][3] ~^ image[23][15] + kernel[1][4] ~^ image[23][16] + kernel[2][0] ~^ image[24][12] + kernel[2][1] ~^ image[24][13] + kernel[2][2] ~^ image[24][14] + kernel[2][3] ~^ image[24][15] + kernel[2][4] ~^ image[24][16] + kernel[3][0] ~^ image[25][12] + kernel[3][1] ~^ image[25][13] + kernel[3][2] ~^ image[25][14] + kernel[3][3] ~^ image[25][15] + kernel[3][4] ~^ image[25][16] + kernel[4][0] ~^ image[26][12] + kernel[4][1] ~^ image[26][13] + kernel[4][2] ~^ image[26][14] + kernel[4][3] ~^ image[26][15] + kernel[4][4] ~^ image[26][16];
assign xor_sum[22][13] = kernel[0][0] ~^ image[22][13] + kernel[0][1] ~^ image[22][14] + kernel[0][2] ~^ image[22][15] + kernel[0][3] ~^ image[22][16] + kernel[0][4] ~^ image[22][17] + kernel[1][0] ~^ image[23][13] + kernel[1][1] ~^ image[23][14] + kernel[1][2] ~^ image[23][15] + kernel[1][3] ~^ image[23][16] + kernel[1][4] ~^ image[23][17] + kernel[2][0] ~^ image[24][13] + kernel[2][1] ~^ image[24][14] + kernel[2][2] ~^ image[24][15] + kernel[2][3] ~^ image[24][16] + kernel[2][4] ~^ image[24][17] + kernel[3][0] ~^ image[25][13] + kernel[3][1] ~^ image[25][14] + kernel[3][2] ~^ image[25][15] + kernel[3][3] ~^ image[25][16] + kernel[3][4] ~^ image[25][17] + kernel[4][0] ~^ image[26][13] + kernel[4][1] ~^ image[26][14] + kernel[4][2] ~^ image[26][15] + kernel[4][3] ~^ image[26][16] + kernel[4][4] ~^ image[26][17];
assign xor_sum[22][14] = kernel[0][0] ~^ image[22][14] + kernel[0][1] ~^ image[22][15] + kernel[0][2] ~^ image[22][16] + kernel[0][3] ~^ image[22][17] + kernel[0][4] ~^ image[22][18] + kernel[1][0] ~^ image[23][14] + kernel[1][1] ~^ image[23][15] + kernel[1][2] ~^ image[23][16] + kernel[1][3] ~^ image[23][17] + kernel[1][4] ~^ image[23][18] + kernel[2][0] ~^ image[24][14] + kernel[2][1] ~^ image[24][15] + kernel[2][2] ~^ image[24][16] + kernel[2][3] ~^ image[24][17] + kernel[2][4] ~^ image[24][18] + kernel[3][0] ~^ image[25][14] + kernel[3][1] ~^ image[25][15] + kernel[3][2] ~^ image[25][16] + kernel[3][3] ~^ image[25][17] + kernel[3][4] ~^ image[25][18] + kernel[4][0] ~^ image[26][14] + kernel[4][1] ~^ image[26][15] + kernel[4][2] ~^ image[26][16] + kernel[4][3] ~^ image[26][17] + kernel[4][4] ~^ image[26][18];
assign xor_sum[22][15] = kernel[0][0] ~^ image[22][15] + kernel[0][1] ~^ image[22][16] + kernel[0][2] ~^ image[22][17] + kernel[0][3] ~^ image[22][18] + kernel[0][4] ~^ image[22][19] + kernel[1][0] ~^ image[23][15] + kernel[1][1] ~^ image[23][16] + kernel[1][2] ~^ image[23][17] + kernel[1][3] ~^ image[23][18] + kernel[1][4] ~^ image[23][19] + kernel[2][0] ~^ image[24][15] + kernel[2][1] ~^ image[24][16] + kernel[2][2] ~^ image[24][17] + kernel[2][3] ~^ image[24][18] + kernel[2][4] ~^ image[24][19] + kernel[3][0] ~^ image[25][15] + kernel[3][1] ~^ image[25][16] + kernel[3][2] ~^ image[25][17] + kernel[3][3] ~^ image[25][18] + kernel[3][4] ~^ image[25][19] + kernel[4][0] ~^ image[26][15] + kernel[4][1] ~^ image[26][16] + kernel[4][2] ~^ image[26][17] + kernel[4][3] ~^ image[26][18] + kernel[4][4] ~^ image[26][19];
assign xor_sum[22][16] = kernel[0][0] ~^ image[22][16] + kernel[0][1] ~^ image[22][17] + kernel[0][2] ~^ image[22][18] + kernel[0][3] ~^ image[22][19] + kernel[0][4] ~^ image[22][20] + kernel[1][0] ~^ image[23][16] + kernel[1][1] ~^ image[23][17] + kernel[1][2] ~^ image[23][18] + kernel[1][3] ~^ image[23][19] + kernel[1][4] ~^ image[23][20] + kernel[2][0] ~^ image[24][16] + kernel[2][1] ~^ image[24][17] + kernel[2][2] ~^ image[24][18] + kernel[2][3] ~^ image[24][19] + kernel[2][4] ~^ image[24][20] + kernel[3][0] ~^ image[25][16] + kernel[3][1] ~^ image[25][17] + kernel[3][2] ~^ image[25][18] + kernel[3][3] ~^ image[25][19] + kernel[3][4] ~^ image[25][20] + kernel[4][0] ~^ image[26][16] + kernel[4][1] ~^ image[26][17] + kernel[4][2] ~^ image[26][18] + kernel[4][3] ~^ image[26][19] + kernel[4][4] ~^ image[26][20];
assign xor_sum[22][17] = kernel[0][0] ~^ image[22][17] + kernel[0][1] ~^ image[22][18] + kernel[0][2] ~^ image[22][19] + kernel[0][3] ~^ image[22][20] + kernel[0][4] ~^ image[22][21] + kernel[1][0] ~^ image[23][17] + kernel[1][1] ~^ image[23][18] + kernel[1][2] ~^ image[23][19] + kernel[1][3] ~^ image[23][20] + kernel[1][4] ~^ image[23][21] + kernel[2][0] ~^ image[24][17] + kernel[2][1] ~^ image[24][18] + kernel[2][2] ~^ image[24][19] + kernel[2][3] ~^ image[24][20] + kernel[2][4] ~^ image[24][21] + kernel[3][0] ~^ image[25][17] + kernel[3][1] ~^ image[25][18] + kernel[3][2] ~^ image[25][19] + kernel[3][3] ~^ image[25][20] + kernel[3][4] ~^ image[25][21] + kernel[4][0] ~^ image[26][17] + kernel[4][1] ~^ image[26][18] + kernel[4][2] ~^ image[26][19] + kernel[4][3] ~^ image[26][20] + kernel[4][4] ~^ image[26][21];
assign xor_sum[22][18] = kernel[0][0] ~^ image[22][18] + kernel[0][1] ~^ image[22][19] + kernel[0][2] ~^ image[22][20] + kernel[0][3] ~^ image[22][21] + kernel[0][4] ~^ image[22][22] + kernel[1][0] ~^ image[23][18] + kernel[1][1] ~^ image[23][19] + kernel[1][2] ~^ image[23][20] + kernel[1][3] ~^ image[23][21] + kernel[1][4] ~^ image[23][22] + kernel[2][0] ~^ image[24][18] + kernel[2][1] ~^ image[24][19] + kernel[2][2] ~^ image[24][20] + kernel[2][3] ~^ image[24][21] + kernel[2][4] ~^ image[24][22] + kernel[3][0] ~^ image[25][18] + kernel[3][1] ~^ image[25][19] + kernel[3][2] ~^ image[25][20] + kernel[3][3] ~^ image[25][21] + kernel[3][4] ~^ image[25][22] + kernel[4][0] ~^ image[26][18] + kernel[4][1] ~^ image[26][19] + kernel[4][2] ~^ image[26][20] + kernel[4][3] ~^ image[26][21] + kernel[4][4] ~^ image[26][22];
assign xor_sum[22][19] = kernel[0][0] ~^ image[22][19] + kernel[0][1] ~^ image[22][20] + kernel[0][2] ~^ image[22][21] + kernel[0][3] ~^ image[22][22] + kernel[0][4] ~^ image[22][23] + kernel[1][0] ~^ image[23][19] + kernel[1][1] ~^ image[23][20] + kernel[1][2] ~^ image[23][21] + kernel[1][3] ~^ image[23][22] + kernel[1][4] ~^ image[23][23] + kernel[2][0] ~^ image[24][19] + kernel[2][1] ~^ image[24][20] + kernel[2][2] ~^ image[24][21] + kernel[2][3] ~^ image[24][22] + kernel[2][4] ~^ image[24][23] + kernel[3][0] ~^ image[25][19] + kernel[3][1] ~^ image[25][20] + kernel[3][2] ~^ image[25][21] + kernel[3][3] ~^ image[25][22] + kernel[3][4] ~^ image[25][23] + kernel[4][0] ~^ image[26][19] + kernel[4][1] ~^ image[26][20] + kernel[4][2] ~^ image[26][21] + kernel[4][3] ~^ image[26][22] + kernel[4][4] ~^ image[26][23];
assign xor_sum[22][20] = kernel[0][0] ~^ image[22][20] + kernel[0][1] ~^ image[22][21] + kernel[0][2] ~^ image[22][22] + kernel[0][3] ~^ image[22][23] + kernel[0][4] ~^ image[22][24] + kernel[1][0] ~^ image[23][20] + kernel[1][1] ~^ image[23][21] + kernel[1][2] ~^ image[23][22] + kernel[1][3] ~^ image[23][23] + kernel[1][4] ~^ image[23][24] + kernel[2][0] ~^ image[24][20] + kernel[2][1] ~^ image[24][21] + kernel[2][2] ~^ image[24][22] + kernel[2][3] ~^ image[24][23] + kernel[2][4] ~^ image[24][24] + kernel[3][0] ~^ image[25][20] + kernel[3][1] ~^ image[25][21] + kernel[3][2] ~^ image[25][22] + kernel[3][3] ~^ image[25][23] + kernel[3][4] ~^ image[25][24] + kernel[4][0] ~^ image[26][20] + kernel[4][1] ~^ image[26][21] + kernel[4][2] ~^ image[26][22] + kernel[4][3] ~^ image[26][23] + kernel[4][4] ~^ image[26][24];
assign xor_sum[22][21] = kernel[0][0] ~^ image[22][21] + kernel[0][1] ~^ image[22][22] + kernel[0][2] ~^ image[22][23] + kernel[0][3] ~^ image[22][24] + kernel[0][4] ~^ image[22][25] + kernel[1][0] ~^ image[23][21] + kernel[1][1] ~^ image[23][22] + kernel[1][2] ~^ image[23][23] + kernel[1][3] ~^ image[23][24] + kernel[1][4] ~^ image[23][25] + kernel[2][0] ~^ image[24][21] + kernel[2][1] ~^ image[24][22] + kernel[2][2] ~^ image[24][23] + kernel[2][3] ~^ image[24][24] + kernel[2][4] ~^ image[24][25] + kernel[3][0] ~^ image[25][21] + kernel[3][1] ~^ image[25][22] + kernel[3][2] ~^ image[25][23] + kernel[3][3] ~^ image[25][24] + kernel[3][4] ~^ image[25][25] + kernel[4][0] ~^ image[26][21] + kernel[4][1] ~^ image[26][22] + kernel[4][2] ~^ image[26][23] + kernel[4][3] ~^ image[26][24] + kernel[4][4] ~^ image[26][25];
assign xor_sum[22][22] = kernel[0][0] ~^ image[22][22] + kernel[0][1] ~^ image[22][23] + kernel[0][2] ~^ image[22][24] + kernel[0][3] ~^ image[22][25] + kernel[0][4] ~^ image[22][26] + kernel[1][0] ~^ image[23][22] + kernel[1][1] ~^ image[23][23] + kernel[1][2] ~^ image[23][24] + kernel[1][3] ~^ image[23][25] + kernel[1][4] ~^ image[23][26] + kernel[2][0] ~^ image[24][22] + kernel[2][1] ~^ image[24][23] + kernel[2][2] ~^ image[24][24] + kernel[2][3] ~^ image[24][25] + kernel[2][4] ~^ image[24][26] + kernel[3][0] ~^ image[25][22] + kernel[3][1] ~^ image[25][23] + kernel[3][2] ~^ image[25][24] + kernel[3][3] ~^ image[25][25] + kernel[3][4] ~^ image[25][26] + kernel[4][0] ~^ image[26][22] + kernel[4][1] ~^ image[26][23] + kernel[4][2] ~^ image[26][24] + kernel[4][3] ~^ image[26][25] + kernel[4][4] ~^ image[26][26];
assign xor_sum[22][23] = kernel[0][0] ~^ image[22][23] + kernel[0][1] ~^ image[22][24] + kernel[0][2] ~^ image[22][25] + kernel[0][3] ~^ image[22][26] + kernel[0][4] ~^ image[22][27] + kernel[1][0] ~^ image[23][23] + kernel[1][1] ~^ image[23][24] + kernel[1][2] ~^ image[23][25] + kernel[1][3] ~^ image[23][26] + kernel[1][4] ~^ image[23][27] + kernel[2][0] ~^ image[24][23] + kernel[2][1] ~^ image[24][24] + kernel[2][2] ~^ image[24][25] + kernel[2][3] ~^ image[24][26] + kernel[2][4] ~^ image[24][27] + kernel[3][0] ~^ image[25][23] + kernel[3][1] ~^ image[25][24] + kernel[3][2] ~^ image[25][25] + kernel[3][3] ~^ image[25][26] + kernel[3][4] ~^ image[25][27] + kernel[4][0] ~^ image[26][23] + kernel[4][1] ~^ image[26][24] + kernel[4][2] ~^ image[26][25] + kernel[4][3] ~^ image[26][26] + kernel[4][4] ~^ image[26][27];
assign xor_sum[23][0] = kernel[0][0] ~^ image[23][0] + kernel[0][1] ~^ image[23][1] + kernel[0][2] ~^ image[23][2] + kernel[0][3] ~^ image[23][3] + kernel[0][4] ~^ image[23][4] + kernel[1][0] ~^ image[24][0] + kernel[1][1] ~^ image[24][1] + kernel[1][2] ~^ image[24][2] + kernel[1][3] ~^ image[24][3] + kernel[1][4] ~^ image[24][4] + kernel[2][0] ~^ image[25][0] + kernel[2][1] ~^ image[25][1] + kernel[2][2] ~^ image[25][2] + kernel[2][3] ~^ image[25][3] + kernel[2][4] ~^ image[25][4] + kernel[3][0] ~^ image[26][0] + kernel[3][1] ~^ image[26][1] + kernel[3][2] ~^ image[26][2] + kernel[3][3] ~^ image[26][3] + kernel[3][4] ~^ image[26][4] + kernel[4][0] ~^ image[27][0] + kernel[4][1] ~^ image[27][1] + kernel[4][2] ~^ image[27][2] + kernel[4][3] ~^ image[27][3] + kernel[4][4] ~^ image[27][4];
assign xor_sum[23][1] = kernel[0][0] ~^ image[23][1] + kernel[0][1] ~^ image[23][2] + kernel[0][2] ~^ image[23][3] + kernel[0][3] ~^ image[23][4] + kernel[0][4] ~^ image[23][5] + kernel[1][0] ~^ image[24][1] + kernel[1][1] ~^ image[24][2] + kernel[1][2] ~^ image[24][3] + kernel[1][3] ~^ image[24][4] + kernel[1][4] ~^ image[24][5] + kernel[2][0] ~^ image[25][1] + kernel[2][1] ~^ image[25][2] + kernel[2][2] ~^ image[25][3] + kernel[2][3] ~^ image[25][4] + kernel[2][4] ~^ image[25][5] + kernel[3][0] ~^ image[26][1] + kernel[3][1] ~^ image[26][2] + kernel[3][2] ~^ image[26][3] + kernel[3][3] ~^ image[26][4] + kernel[3][4] ~^ image[26][5] + kernel[4][0] ~^ image[27][1] + kernel[4][1] ~^ image[27][2] + kernel[4][2] ~^ image[27][3] + kernel[4][3] ~^ image[27][4] + kernel[4][4] ~^ image[27][5];
assign xor_sum[23][2] = kernel[0][0] ~^ image[23][2] + kernel[0][1] ~^ image[23][3] + kernel[0][2] ~^ image[23][4] + kernel[0][3] ~^ image[23][5] + kernel[0][4] ~^ image[23][6] + kernel[1][0] ~^ image[24][2] + kernel[1][1] ~^ image[24][3] + kernel[1][2] ~^ image[24][4] + kernel[1][3] ~^ image[24][5] + kernel[1][4] ~^ image[24][6] + kernel[2][0] ~^ image[25][2] + kernel[2][1] ~^ image[25][3] + kernel[2][2] ~^ image[25][4] + kernel[2][3] ~^ image[25][5] + kernel[2][4] ~^ image[25][6] + kernel[3][0] ~^ image[26][2] + kernel[3][1] ~^ image[26][3] + kernel[3][2] ~^ image[26][4] + kernel[3][3] ~^ image[26][5] + kernel[3][4] ~^ image[26][6] + kernel[4][0] ~^ image[27][2] + kernel[4][1] ~^ image[27][3] + kernel[4][2] ~^ image[27][4] + kernel[4][3] ~^ image[27][5] + kernel[4][4] ~^ image[27][6];
assign xor_sum[23][3] = kernel[0][0] ~^ image[23][3] + kernel[0][1] ~^ image[23][4] + kernel[0][2] ~^ image[23][5] + kernel[0][3] ~^ image[23][6] + kernel[0][4] ~^ image[23][7] + kernel[1][0] ~^ image[24][3] + kernel[1][1] ~^ image[24][4] + kernel[1][2] ~^ image[24][5] + kernel[1][3] ~^ image[24][6] + kernel[1][4] ~^ image[24][7] + kernel[2][0] ~^ image[25][3] + kernel[2][1] ~^ image[25][4] + kernel[2][2] ~^ image[25][5] + kernel[2][3] ~^ image[25][6] + kernel[2][4] ~^ image[25][7] + kernel[3][0] ~^ image[26][3] + kernel[3][1] ~^ image[26][4] + kernel[3][2] ~^ image[26][5] + kernel[3][3] ~^ image[26][6] + kernel[3][4] ~^ image[26][7] + kernel[4][0] ~^ image[27][3] + kernel[4][1] ~^ image[27][4] + kernel[4][2] ~^ image[27][5] + kernel[4][3] ~^ image[27][6] + kernel[4][4] ~^ image[27][7];
assign xor_sum[23][4] = kernel[0][0] ~^ image[23][4] + kernel[0][1] ~^ image[23][5] + kernel[0][2] ~^ image[23][6] + kernel[0][3] ~^ image[23][7] + kernel[0][4] ~^ image[23][8] + kernel[1][0] ~^ image[24][4] + kernel[1][1] ~^ image[24][5] + kernel[1][2] ~^ image[24][6] + kernel[1][3] ~^ image[24][7] + kernel[1][4] ~^ image[24][8] + kernel[2][0] ~^ image[25][4] + kernel[2][1] ~^ image[25][5] + kernel[2][2] ~^ image[25][6] + kernel[2][3] ~^ image[25][7] + kernel[2][4] ~^ image[25][8] + kernel[3][0] ~^ image[26][4] + kernel[3][1] ~^ image[26][5] + kernel[3][2] ~^ image[26][6] + kernel[3][3] ~^ image[26][7] + kernel[3][4] ~^ image[26][8] + kernel[4][0] ~^ image[27][4] + kernel[4][1] ~^ image[27][5] + kernel[4][2] ~^ image[27][6] + kernel[4][3] ~^ image[27][7] + kernel[4][4] ~^ image[27][8];
assign xor_sum[23][5] = kernel[0][0] ~^ image[23][5] + kernel[0][1] ~^ image[23][6] + kernel[0][2] ~^ image[23][7] + kernel[0][3] ~^ image[23][8] + kernel[0][4] ~^ image[23][9] + kernel[1][0] ~^ image[24][5] + kernel[1][1] ~^ image[24][6] + kernel[1][2] ~^ image[24][7] + kernel[1][3] ~^ image[24][8] + kernel[1][4] ~^ image[24][9] + kernel[2][0] ~^ image[25][5] + kernel[2][1] ~^ image[25][6] + kernel[2][2] ~^ image[25][7] + kernel[2][3] ~^ image[25][8] + kernel[2][4] ~^ image[25][9] + kernel[3][0] ~^ image[26][5] + kernel[3][1] ~^ image[26][6] + kernel[3][2] ~^ image[26][7] + kernel[3][3] ~^ image[26][8] + kernel[3][4] ~^ image[26][9] + kernel[4][0] ~^ image[27][5] + kernel[4][1] ~^ image[27][6] + kernel[4][2] ~^ image[27][7] + kernel[4][3] ~^ image[27][8] + kernel[4][4] ~^ image[27][9];
assign xor_sum[23][6] = kernel[0][0] ~^ image[23][6] + kernel[0][1] ~^ image[23][7] + kernel[0][2] ~^ image[23][8] + kernel[0][3] ~^ image[23][9] + kernel[0][4] ~^ image[23][10] + kernel[1][0] ~^ image[24][6] + kernel[1][1] ~^ image[24][7] + kernel[1][2] ~^ image[24][8] + kernel[1][3] ~^ image[24][9] + kernel[1][4] ~^ image[24][10] + kernel[2][0] ~^ image[25][6] + kernel[2][1] ~^ image[25][7] + kernel[2][2] ~^ image[25][8] + kernel[2][3] ~^ image[25][9] + kernel[2][4] ~^ image[25][10] + kernel[3][0] ~^ image[26][6] + kernel[3][1] ~^ image[26][7] + kernel[3][2] ~^ image[26][8] + kernel[3][3] ~^ image[26][9] + kernel[3][4] ~^ image[26][10] + kernel[4][0] ~^ image[27][6] + kernel[4][1] ~^ image[27][7] + kernel[4][2] ~^ image[27][8] + kernel[4][3] ~^ image[27][9] + kernel[4][4] ~^ image[27][10];
assign xor_sum[23][7] = kernel[0][0] ~^ image[23][7] + kernel[0][1] ~^ image[23][8] + kernel[0][2] ~^ image[23][9] + kernel[0][3] ~^ image[23][10] + kernel[0][4] ~^ image[23][11] + kernel[1][0] ~^ image[24][7] + kernel[1][1] ~^ image[24][8] + kernel[1][2] ~^ image[24][9] + kernel[1][3] ~^ image[24][10] + kernel[1][4] ~^ image[24][11] + kernel[2][0] ~^ image[25][7] + kernel[2][1] ~^ image[25][8] + kernel[2][2] ~^ image[25][9] + kernel[2][3] ~^ image[25][10] + kernel[2][4] ~^ image[25][11] + kernel[3][0] ~^ image[26][7] + kernel[3][1] ~^ image[26][8] + kernel[3][2] ~^ image[26][9] + kernel[3][3] ~^ image[26][10] + kernel[3][4] ~^ image[26][11] + kernel[4][0] ~^ image[27][7] + kernel[4][1] ~^ image[27][8] + kernel[4][2] ~^ image[27][9] + kernel[4][3] ~^ image[27][10] + kernel[4][4] ~^ image[27][11];
assign xor_sum[23][8] = kernel[0][0] ~^ image[23][8] + kernel[0][1] ~^ image[23][9] + kernel[0][2] ~^ image[23][10] + kernel[0][3] ~^ image[23][11] + kernel[0][4] ~^ image[23][12] + kernel[1][0] ~^ image[24][8] + kernel[1][1] ~^ image[24][9] + kernel[1][2] ~^ image[24][10] + kernel[1][3] ~^ image[24][11] + kernel[1][4] ~^ image[24][12] + kernel[2][0] ~^ image[25][8] + kernel[2][1] ~^ image[25][9] + kernel[2][2] ~^ image[25][10] + kernel[2][3] ~^ image[25][11] + kernel[2][4] ~^ image[25][12] + kernel[3][0] ~^ image[26][8] + kernel[3][1] ~^ image[26][9] + kernel[3][2] ~^ image[26][10] + kernel[3][3] ~^ image[26][11] + kernel[3][4] ~^ image[26][12] + kernel[4][0] ~^ image[27][8] + kernel[4][1] ~^ image[27][9] + kernel[4][2] ~^ image[27][10] + kernel[4][3] ~^ image[27][11] + kernel[4][4] ~^ image[27][12];
assign xor_sum[23][9] = kernel[0][0] ~^ image[23][9] + kernel[0][1] ~^ image[23][10] + kernel[0][2] ~^ image[23][11] + kernel[0][3] ~^ image[23][12] + kernel[0][4] ~^ image[23][13] + kernel[1][0] ~^ image[24][9] + kernel[1][1] ~^ image[24][10] + kernel[1][2] ~^ image[24][11] + kernel[1][3] ~^ image[24][12] + kernel[1][4] ~^ image[24][13] + kernel[2][0] ~^ image[25][9] + kernel[2][1] ~^ image[25][10] + kernel[2][2] ~^ image[25][11] + kernel[2][3] ~^ image[25][12] + kernel[2][4] ~^ image[25][13] + kernel[3][0] ~^ image[26][9] + kernel[3][1] ~^ image[26][10] + kernel[3][2] ~^ image[26][11] + kernel[3][3] ~^ image[26][12] + kernel[3][4] ~^ image[26][13] + kernel[4][0] ~^ image[27][9] + kernel[4][1] ~^ image[27][10] + kernel[4][2] ~^ image[27][11] + kernel[4][3] ~^ image[27][12] + kernel[4][4] ~^ image[27][13];
assign xor_sum[23][10] = kernel[0][0] ~^ image[23][10] + kernel[0][1] ~^ image[23][11] + kernel[0][2] ~^ image[23][12] + kernel[0][3] ~^ image[23][13] + kernel[0][4] ~^ image[23][14] + kernel[1][0] ~^ image[24][10] + kernel[1][1] ~^ image[24][11] + kernel[1][2] ~^ image[24][12] + kernel[1][3] ~^ image[24][13] + kernel[1][4] ~^ image[24][14] + kernel[2][0] ~^ image[25][10] + kernel[2][1] ~^ image[25][11] + kernel[2][2] ~^ image[25][12] + kernel[2][3] ~^ image[25][13] + kernel[2][4] ~^ image[25][14] + kernel[3][0] ~^ image[26][10] + kernel[3][1] ~^ image[26][11] + kernel[3][2] ~^ image[26][12] + kernel[3][3] ~^ image[26][13] + kernel[3][4] ~^ image[26][14] + kernel[4][0] ~^ image[27][10] + kernel[4][1] ~^ image[27][11] + kernel[4][2] ~^ image[27][12] + kernel[4][3] ~^ image[27][13] + kernel[4][4] ~^ image[27][14];
assign xor_sum[23][11] = kernel[0][0] ~^ image[23][11] + kernel[0][1] ~^ image[23][12] + kernel[0][2] ~^ image[23][13] + kernel[0][3] ~^ image[23][14] + kernel[0][4] ~^ image[23][15] + kernel[1][0] ~^ image[24][11] + kernel[1][1] ~^ image[24][12] + kernel[1][2] ~^ image[24][13] + kernel[1][3] ~^ image[24][14] + kernel[1][4] ~^ image[24][15] + kernel[2][0] ~^ image[25][11] + kernel[2][1] ~^ image[25][12] + kernel[2][2] ~^ image[25][13] + kernel[2][3] ~^ image[25][14] + kernel[2][4] ~^ image[25][15] + kernel[3][0] ~^ image[26][11] + kernel[3][1] ~^ image[26][12] + kernel[3][2] ~^ image[26][13] + kernel[3][3] ~^ image[26][14] + kernel[3][4] ~^ image[26][15] + kernel[4][0] ~^ image[27][11] + kernel[4][1] ~^ image[27][12] + kernel[4][2] ~^ image[27][13] + kernel[4][3] ~^ image[27][14] + kernel[4][4] ~^ image[27][15];
assign xor_sum[23][12] = kernel[0][0] ~^ image[23][12] + kernel[0][1] ~^ image[23][13] + kernel[0][2] ~^ image[23][14] + kernel[0][3] ~^ image[23][15] + kernel[0][4] ~^ image[23][16] + kernel[1][0] ~^ image[24][12] + kernel[1][1] ~^ image[24][13] + kernel[1][2] ~^ image[24][14] + kernel[1][3] ~^ image[24][15] + kernel[1][4] ~^ image[24][16] + kernel[2][0] ~^ image[25][12] + kernel[2][1] ~^ image[25][13] + kernel[2][2] ~^ image[25][14] + kernel[2][3] ~^ image[25][15] + kernel[2][4] ~^ image[25][16] + kernel[3][0] ~^ image[26][12] + kernel[3][1] ~^ image[26][13] + kernel[3][2] ~^ image[26][14] + kernel[3][3] ~^ image[26][15] + kernel[3][4] ~^ image[26][16] + kernel[4][0] ~^ image[27][12] + kernel[4][1] ~^ image[27][13] + kernel[4][2] ~^ image[27][14] + kernel[4][3] ~^ image[27][15] + kernel[4][4] ~^ image[27][16];
assign xor_sum[23][13] = kernel[0][0] ~^ image[23][13] + kernel[0][1] ~^ image[23][14] + kernel[0][2] ~^ image[23][15] + kernel[0][3] ~^ image[23][16] + kernel[0][4] ~^ image[23][17] + kernel[1][0] ~^ image[24][13] + kernel[1][1] ~^ image[24][14] + kernel[1][2] ~^ image[24][15] + kernel[1][3] ~^ image[24][16] + kernel[1][4] ~^ image[24][17] + kernel[2][0] ~^ image[25][13] + kernel[2][1] ~^ image[25][14] + kernel[2][2] ~^ image[25][15] + kernel[2][3] ~^ image[25][16] + kernel[2][4] ~^ image[25][17] + kernel[3][0] ~^ image[26][13] + kernel[3][1] ~^ image[26][14] + kernel[3][2] ~^ image[26][15] + kernel[3][3] ~^ image[26][16] + kernel[3][4] ~^ image[26][17] + kernel[4][0] ~^ image[27][13] + kernel[4][1] ~^ image[27][14] + kernel[4][2] ~^ image[27][15] + kernel[4][3] ~^ image[27][16] + kernel[4][4] ~^ image[27][17];
assign xor_sum[23][14] = kernel[0][0] ~^ image[23][14] + kernel[0][1] ~^ image[23][15] + kernel[0][2] ~^ image[23][16] + kernel[0][3] ~^ image[23][17] + kernel[0][4] ~^ image[23][18] + kernel[1][0] ~^ image[24][14] + kernel[1][1] ~^ image[24][15] + kernel[1][2] ~^ image[24][16] + kernel[1][3] ~^ image[24][17] + kernel[1][4] ~^ image[24][18] + kernel[2][0] ~^ image[25][14] + kernel[2][1] ~^ image[25][15] + kernel[2][2] ~^ image[25][16] + kernel[2][3] ~^ image[25][17] + kernel[2][4] ~^ image[25][18] + kernel[3][0] ~^ image[26][14] + kernel[3][1] ~^ image[26][15] + kernel[3][2] ~^ image[26][16] + kernel[3][3] ~^ image[26][17] + kernel[3][4] ~^ image[26][18] + kernel[4][0] ~^ image[27][14] + kernel[4][1] ~^ image[27][15] + kernel[4][2] ~^ image[27][16] + kernel[4][3] ~^ image[27][17] + kernel[4][4] ~^ image[27][18];
assign xor_sum[23][15] = kernel[0][0] ~^ image[23][15] + kernel[0][1] ~^ image[23][16] + kernel[0][2] ~^ image[23][17] + kernel[0][3] ~^ image[23][18] + kernel[0][4] ~^ image[23][19] + kernel[1][0] ~^ image[24][15] + kernel[1][1] ~^ image[24][16] + kernel[1][2] ~^ image[24][17] + kernel[1][3] ~^ image[24][18] + kernel[1][4] ~^ image[24][19] + kernel[2][0] ~^ image[25][15] + kernel[2][1] ~^ image[25][16] + kernel[2][2] ~^ image[25][17] + kernel[2][3] ~^ image[25][18] + kernel[2][4] ~^ image[25][19] + kernel[3][0] ~^ image[26][15] + kernel[3][1] ~^ image[26][16] + kernel[3][2] ~^ image[26][17] + kernel[3][3] ~^ image[26][18] + kernel[3][4] ~^ image[26][19] + kernel[4][0] ~^ image[27][15] + kernel[4][1] ~^ image[27][16] + kernel[4][2] ~^ image[27][17] + kernel[4][3] ~^ image[27][18] + kernel[4][4] ~^ image[27][19];
assign xor_sum[23][16] = kernel[0][0] ~^ image[23][16] + kernel[0][1] ~^ image[23][17] + kernel[0][2] ~^ image[23][18] + kernel[0][3] ~^ image[23][19] + kernel[0][4] ~^ image[23][20] + kernel[1][0] ~^ image[24][16] + kernel[1][1] ~^ image[24][17] + kernel[1][2] ~^ image[24][18] + kernel[1][3] ~^ image[24][19] + kernel[1][4] ~^ image[24][20] + kernel[2][0] ~^ image[25][16] + kernel[2][1] ~^ image[25][17] + kernel[2][2] ~^ image[25][18] + kernel[2][3] ~^ image[25][19] + kernel[2][4] ~^ image[25][20] + kernel[3][0] ~^ image[26][16] + kernel[3][1] ~^ image[26][17] + kernel[3][2] ~^ image[26][18] + kernel[3][3] ~^ image[26][19] + kernel[3][4] ~^ image[26][20] + kernel[4][0] ~^ image[27][16] + kernel[4][1] ~^ image[27][17] + kernel[4][2] ~^ image[27][18] + kernel[4][3] ~^ image[27][19] + kernel[4][4] ~^ image[27][20];
assign xor_sum[23][17] = kernel[0][0] ~^ image[23][17] + kernel[0][1] ~^ image[23][18] + kernel[0][2] ~^ image[23][19] + kernel[0][3] ~^ image[23][20] + kernel[0][4] ~^ image[23][21] + kernel[1][0] ~^ image[24][17] + kernel[1][1] ~^ image[24][18] + kernel[1][2] ~^ image[24][19] + kernel[1][3] ~^ image[24][20] + kernel[1][4] ~^ image[24][21] + kernel[2][0] ~^ image[25][17] + kernel[2][1] ~^ image[25][18] + kernel[2][2] ~^ image[25][19] + kernel[2][3] ~^ image[25][20] + kernel[2][4] ~^ image[25][21] + kernel[3][0] ~^ image[26][17] + kernel[3][1] ~^ image[26][18] + kernel[3][2] ~^ image[26][19] + kernel[3][3] ~^ image[26][20] + kernel[3][4] ~^ image[26][21] + kernel[4][0] ~^ image[27][17] + kernel[4][1] ~^ image[27][18] + kernel[4][2] ~^ image[27][19] + kernel[4][3] ~^ image[27][20] + kernel[4][4] ~^ image[27][21];
assign xor_sum[23][18] = kernel[0][0] ~^ image[23][18] + kernel[0][1] ~^ image[23][19] + kernel[0][2] ~^ image[23][20] + kernel[0][3] ~^ image[23][21] + kernel[0][4] ~^ image[23][22] + kernel[1][0] ~^ image[24][18] + kernel[1][1] ~^ image[24][19] + kernel[1][2] ~^ image[24][20] + kernel[1][3] ~^ image[24][21] + kernel[1][4] ~^ image[24][22] + kernel[2][0] ~^ image[25][18] + kernel[2][1] ~^ image[25][19] + kernel[2][2] ~^ image[25][20] + kernel[2][3] ~^ image[25][21] + kernel[2][4] ~^ image[25][22] + kernel[3][0] ~^ image[26][18] + kernel[3][1] ~^ image[26][19] + kernel[3][2] ~^ image[26][20] + kernel[3][3] ~^ image[26][21] + kernel[3][4] ~^ image[26][22] + kernel[4][0] ~^ image[27][18] + kernel[4][1] ~^ image[27][19] + kernel[4][2] ~^ image[27][20] + kernel[4][3] ~^ image[27][21] + kernel[4][4] ~^ image[27][22];
assign xor_sum[23][19] = kernel[0][0] ~^ image[23][19] + kernel[0][1] ~^ image[23][20] + kernel[0][2] ~^ image[23][21] + kernel[0][3] ~^ image[23][22] + kernel[0][4] ~^ image[23][23] + kernel[1][0] ~^ image[24][19] + kernel[1][1] ~^ image[24][20] + kernel[1][2] ~^ image[24][21] + kernel[1][3] ~^ image[24][22] + kernel[1][4] ~^ image[24][23] + kernel[2][0] ~^ image[25][19] + kernel[2][1] ~^ image[25][20] + kernel[2][2] ~^ image[25][21] + kernel[2][3] ~^ image[25][22] + kernel[2][4] ~^ image[25][23] + kernel[3][0] ~^ image[26][19] + kernel[3][1] ~^ image[26][20] + kernel[3][2] ~^ image[26][21] + kernel[3][3] ~^ image[26][22] + kernel[3][4] ~^ image[26][23] + kernel[4][0] ~^ image[27][19] + kernel[4][1] ~^ image[27][20] + kernel[4][2] ~^ image[27][21] + kernel[4][3] ~^ image[27][22] + kernel[4][4] ~^ image[27][23];
assign xor_sum[23][20] = kernel[0][0] ~^ image[23][20] + kernel[0][1] ~^ image[23][21] + kernel[0][2] ~^ image[23][22] + kernel[0][3] ~^ image[23][23] + kernel[0][4] ~^ image[23][24] + kernel[1][0] ~^ image[24][20] + kernel[1][1] ~^ image[24][21] + kernel[1][2] ~^ image[24][22] + kernel[1][3] ~^ image[24][23] + kernel[1][4] ~^ image[24][24] + kernel[2][0] ~^ image[25][20] + kernel[2][1] ~^ image[25][21] + kernel[2][2] ~^ image[25][22] + kernel[2][3] ~^ image[25][23] + kernel[2][4] ~^ image[25][24] + kernel[3][0] ~^ image[26][20] + kernel[3][1] ~^ image[26][21] + kernel[3][2] ~^ image[26][22] + kernel[3][3] ~^ image[26][23] + kernel[3][4] ~^ image[26][24] + kernel[4][0] ~^ image[27][20] + kernel[4][1] ~^ image[27][21] + kernel[4][2] ~^ image[27][22] + kernel[4][3] ~^ image[27][23] + kernel[4][4] ~^ image[27][24];
assign xor_sum[23][21] = kernel[0][0] ~^ image[23][21] + kernel[0][1] ~^ image[23][22] + kernel[0][2] ~^ image[23][23] + kernel[0][3] ~^ image[23][24] + kernel[0][4] ~^ image[23][25] + kernel[1][0] ~^ image[24][21] + kernel[1][1] ~^ image[24][22] + kernel[1][2] ~^ image[24][23] + kernel[1][3] ~^ image[24][24] + kernel[1][4] ~^ image[24][25] + kernel[2][0] ~^ image[25][21] + kernel[2][1] ~^ image[25][22] + kernel[2][2] ~^ image[25][23] + kernel[2][3] ~^ image[25][24] + kernel[2][4] ~^ image[25][25] + kernel[3][0] ~^ image[26][21] + kernel[3][1] ~^ image[26][22] + kernel[3][2] ~^ image[26][23] + kernel[3][3] ~^ image[26][24] + kernel[3][4] ~^ image[26][25] + kernel[4][0] ~^ image[27][21] + kernel[4][1] ~^ image[27][22] + kernel[4][2] ~^ image[27][23] + kernel[4][3] ~^ image[27][24] + kernel[4][4] ~^ image[27][25];
assign xor_sum[23][22] = kernel[0][0] ~^ image[23][22] + kernel[0][1] ~^ image[23][23] + kernel[0][2] ~^ image[23][24] + kernel[0][3] ~^ image[23][25] + kernel[0][4] ~^ image[23][26] + kernel[1][0] ~^ image[24][22] + kernel[1][1] ~^ image[24][23] + kernel[1][2] ~^ image[24][24] + kernel[1][3] ~^ image[24][25] + kernel[1][4] ~^ image[24][26] + kernel[2][0] ~^ image[25][22] + kernel[2][1] ~^ image[25][23] + kernel[2][2] ~^ image[25][24] + kernel[2][3] ~^ image[25][25] + kernel[2][4] ~^ image[25][26] + kernel[3][0] ~^ image[26][22] + kernel[3][1] ~^ image[26][23] + kernel[3][2] ~^ image[26][24] + kernel[3][3] ~^ image[26][25] + kernel[3][4] ~^ image[26][26] + kernel[4][0] ~^ image[27][22] + kernel[4][1] ~^ image[27][23] + kernel[4][2] ~^ image[27][24] + kernel[4][3] ~^ image[27][25] + kernel[4][4] ~^ image[27][26];
assign xor_sum[23][23] = kernel[0][0] ~^ image[23][23] + kernel[0][1] ~^ image[23][24] + kernel[0][2] ~^ image[23][25] + kernel[0][3] ~^ image[23][26] + kernel[0][4] ~^ image[23][27] + kernel[1][0] ~^ image[24][23] + kernel[1][1] ~^ image[24][24] + kernel[1][2] ~^ image[24][25] + kernel[1][3] ~^ image[24][26] + kernel[1][4] ~^ image[24][27] + kernel[2][0] ~^ image[25][23] + kernel[2][1] ~^ image[25][24] + kernel[2][2] ~^ image[25][25] + kernel[2][3] ~^ image[25][26] + kernel[2][4] ~^ image[25][27] + kernel[3][0] ~^ image[26][23] + kernel[3][1] ~^ image[26][24] + kernel[3][2] ~^ image[26][25] + kernel[3][3] ~^ image[26][26] + kernel[3][4] ~^ image[26][27] + kernel[4][0] ~^ image[27][23] + kernel[4][1] ~^ image[27][24] + kernel[4][2] ~^ image[27][25] + kernel[4][3] ~^ image[27][26] + kernel[4][4] ~^ image[27][27];

endmodule