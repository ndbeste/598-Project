typedef logic          d_image_t    [0:11][0:11];
typedef logic          d_kernel_t   [0: 4][0: 4];
typedef logic [7:0]    d_fmap_out_t [0: 7][0: 7];

module convchan2 
    #( parameter bW = 8 )
    ( 
    input  logic [0:12*12 -1]   i_image    ,
    input  logic [0:5*5   -1]   i_kernel   ,
    output logic [0:8*8*bW-1]   o_out_fmap
    );

d_image_t    image    ;
d_kernel_t   kernel   ;
d_fmap_out_t out_fmap ;

genvar i,j,k;
for (i=0; i<12; i=i+1) begin
    for (j=0; j<12; j=j+1) begin
        assign image[i][j] = i_image[ 12*i + j ];
    end
end

for (i=0; i<5; i=i+1) begin
    for (j=0; j<5; j=j+1) begin
        assign kernel[i][j] = i_kernel[ 5*i + j ];
    end
end

for (i=0; i<8; i=i+1) begin
    for (j=0; j<8; j=j+1) begin
        for (k=0; k<bW; k=k+1) begin
            assign o_out_fmap[i][j][k] = out_fmap[ 8*bW*i + bW*j + k ];
        end
    end
end

assign out_fmap[0][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][0])} + {7'd0,(kernel[0][1] ~^ image[0][1])} + {7'd0,(kernel[0][2] ~^ image[0][2])} + {7'd0,(kernel[0][3] ~^ image[0][3])} + {7'd0,(kernel[0][4] ~^ image[0][4])} + {7'd0,(kernel[1][0] ~^ image[1][0])} + {7'd0,(kernel[1][1] ~^ image[1][1])} + {7'd0,(kernel[1][2] ~^ image[1][2])} + {7'd0,(kernel[1][3] ~^ image[1][3])} + {7'd0,(kernel[1][4] ~^ image[1][4])} + {7'd0,(kernel[2][0] ~^ image[2][0])} + {7'd0,(kernel[2][1] ~^ image[2][1])} + {7'd0,(kernel[2][2] ~^ image[2][2])} + {7'd0,(kernel[2][3] ~^ image[2][3])} + {7'd0,(kernel[2][4] ~^ image[2][4])} + {7'd0,(kernel[3][0] ~^ image[3][0])} + {7'd0,(kernel[3][1] ~^ image[3][1])} + {7'd0,(kernel[3][2] ~^ image[3][2])} + {7'd0,(kernel[3][3] ~^ image[3][3])} + {7'd0,(kernel[3][4] ~^ image[3][4])} + {7'd0,(kernel[4][0] ~^ image[4][0])} + {7'd0,(kernel[4][1] ~^ image[4][1])} + {7'd0,(kernel[4][2] ~^ image[4][2])} + {7'd0,(kernel[4][3] ~^ image[4][3])} + {7'd0,(kernel[4][4] ~^ image[4][4])};
assign out_fmap[0][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][1])} + {7'd0,(kernel[0][1] ~^ image[0][2])} + {7'd0,(kernel[0][2] ~^ image[0][3])} + {7'd0,(kernel[0][3] ~^ image[0][4])} + {7'd0,(kernel[0][4] ~^ image[0][5])} + {7'd0,(kernel[1][0] ~^ image[1][1])} + {7'd0,(kernel[1][1] ~^ image[1][2])} + {7'd0,(kernel[1][2] ~^ image[1][3])} + {7'd0,(kernel[1][3] ~^ image[1][4])} + {7'd0,(kernel[1][4] ~^ image[1][5])} + {7'd0,(kernel[2][0] ~^ image[2][1])} + {7'd0,(kernel[2][1] ~^ image[2][2])} + {7'd0,(kernel[2][2] ~^ image[2][3])} + {7'd0,(kernel[2][3] ~^ image[2][4])} + {7'd0,(kernel[2][4] ~^ image[2][5])} + {7'd0,(kernel[3][0] ~^ image[3][1])} + {7'd0,(kernel[3][1] ~^ image[3][2])} + {7'd0,(kernel[3][2] ~^ image[3][3])} + {7'd0,(kernel[3][3] ~^ image[3][4])} + {7'd0,(kernel[3][4] ~^ image[3][5])} + {7'd0,(kernel[4][0] ~^ image[4][1])} + {7'd0,(kernel[4][1] ~^ image[4][2])} + {7'd0,(kernel[4][2] ~^ image[4][3])} + {7'd0,(kernel[4][3] ~^ image[4][4])} + {7'd0,(kernel[4][4] ~^ image[4][5])};
assign out_fmap[0][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][2])} + {7'd0,(kernel[0][1] ~^ image[0][3])} + {7'd0,(kernel[0][2] ~^ image[0][4])} + {7'd0,(kernel[0][3] ~^ image[0][5])} + {7'd0,(kernel[0][4] ~^ image[0][6])} + {7'd0,(kernel[1][0] ~^ image[1][2])} + {7'd0,(kernel[1][1] ~^ image[1][3])} + {7'd0,(kernel[1][2] ~^ image[1][4])} + {7'd0,(kernel[1][3] ~^ image[1][5])} + {7'd0,(kernel[1][4] ~^ image[1][6])} + {7'd0,(kernel[2][0] ~^ image[2][2])} + {7'd0,(kernel[2][1] ~^ image[2][3])} + {7'd0,(kernel[2][2] ~^ image[2][4])} + {7'd0,(kernel[2][3] ~^ image[2][5])} + {7'd0,(kernel[2][4] ~^ image[2][6])} + {7'd0,(kernel[3][0] ~^ image[3][2])} + {7'd0,(kernel[3][1] ~^ image[3][3])} + {7'd0,(kernel[3][2] ~^ image[3][4])} + {7'd0,(kernel[3][3] ~^ image[3][5])} + {7'd0,(kernel[3][4] ~^ image[3][6])} + {7'd0,(kernel[4][0] ~^ image[4][2])} + {7'd0,(kernel[4][1] ~^ image[4][3])} + {7'd0,(kernel[4][2] ~^ image[4][4])} + {7'd0,(kernel[4][3] ~^ image[4][5])} + {7'd0,(kernel[4][4] ~^ image[4][6])};
assign out_fmap[0][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][3])} + {7'd0,(kernel[0][1] ~^ image[0][4])} + {7'd0,(kernel[0][2] ~^ image[0][5])} + {7'd0,(kernel[0][3] ~^ image[0][6])} + {7'd0,(kernel[0][4] ~^ image[0][7])} + {7'd0,(kernel[1][0] ~^ image[1][3])} + {7'd0,(kernel[1][1] ~^ image[1][4])} + {7'd0,(kernel[1][2] ~^ image[1][5])} + {7'd0,(kernel[1][3] ~^ image[1][6])} + {7'd0,(kernel[1][4] ~^ image[1][7])} + {7'd0,(kernel[2][0] ~^ image[2][3])} + {7'd0,(kernel[2][1] ~^ image[2][4])} + {7'd0,(kernel[2][2] ~^ image[2][5])} + {7'd0,(kernel[2][3] ~^ image[2][6])} + {7'd0,(kernel[2][4] ~^ image[2][7])} + {7'd0,(kernel[3][0] ~^ image[3][3])} + {7'd0,(kernel[3][1] ~^ image[3][4])} + {7'd0,(kernel[3][2] ~^ image[3][5])} + {7'd0,(kernel[3][3] ~^ image[3][6])} + {7'd0,(kernel[3][4] ~^ image[3][7])} + {7'd0,(kernel[4][0] ~^ image[4][3])} + {7'd0,(kernel[4][1] ~^ image[4][4])} + {7'd0,(kernel[4][2] ~^ image[4][5])} + {7'd0,(kernel[4][3] ~^ image[4][6])} + {7'd0,(kernel[4][4] ~^ image[4][7])};
assign out_fmap[0][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][4])} + {7'd0,(kernel[0][1] ~^ image[0][5])} + {7'd0,(kernel[0][2] ~^ image[0][6])} + {7'd0,(kernel[0][3] ~^ image[0][7])} + {7'd0,(kernel[0][4] ~^ image[0][8])} + {7'd0,(kernel[1][0] ~^ image[1][4])} + {7'd0,(kernel[1][1] ~^ image[1][5])} + {7'd0,(kernel[1][2] ~^ image[1][6])} + {7'd0,(kernel[1][3] ~^ image[1][7])} + {7'd0,(kernel[1][4] ~^ image[1][8])} + {7'd0,(kernel[2][0] ~^ image[2][4])} + {7'd0,(kernel[2][1] ~^ image[2][5])} + {7'd0,(kernel[2][2] ~^ image[2][6])} + {7'd0,(kernel[2][3] ~^ image[2][7])} + {7'd0,(kernel[2][4] ~^ image[2][8])} + {7'd0,(kernel[3][0] ~^ image[3][4])} + {7'd0,(kernel[3][1] ~^ image[3][5])} + {7'd0,(kernel[3][2] ~^ image[3][6])} + {7'd0,(kernel[3][3] ~^ image[3][7])} + {7'd0,(kernel[3][4] ~^ image[3][8])} + {7'd0,(kernel[4][0] ~^ image[4][4])} + {7'd0,(kernel[4][1] ~^ image[4][5])} + {7'd0,(kernel[4][2] ~^ image[4][6])} + {7'd0,(kernel[4][3] ~^ image[4][7])} + {7'd0,(kernel[4][4] ~^ image[4][8])};
assign out_fmap[0][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][5])} + {7'd0,(kernel[0][1] ~^ image[0][6])} + {7'd0,(kernel[0][2] ~^ image[0][7])} + {7'd0,(kernel[0][3] ~^ image[0][8])} + {7'd0,(kernel[0][4] ~^ image[0][9])} + {7'd0,(kernel[1][0] ~^ image[1][5])} + {7'd0,(kernel[1][1] ~^ image[1][6])} + {7'd0,(kernel[1][2] ~^ image[1][7])} + {7'd0,(kernel[1][3] ~^ image[1][8])} + {7'd0,(kernel[1][4] ~^ image[1][9])} + {7'd0,(kernel[2][0] ~^ image[2][5])} + {7'd0,(kernel[2][1] ~^ image[2][6])} + {7'd0,(kernel[2][2] ~^ image[2][7])} + {7'd0,(kernel[2][3] ~^ image[2][8])} + {7'd0,(kernel[2][4] ~^ image[2][9])} + {7'd0,(kernel[3][0] ~^ image[3][5])} + {7'd0,(kernel[3][1] ~^ image[3][6])} + {7'd0,(kernel[3][2] ~^ image[3][7])} + {7'd0,(kernel[3][3] ~^ image[3][8])} + {7'd0,(kernel[3][4] ~^ image[3][9])} + {7'd0,(kernel[4][0] ~^ image[4][5])} + {7'd0,(kernel[4][1] ~^ image[4][6])} + {7'd0,(kernel[4][2] ~^ image[4][7])} + {7'd0,(kernel[4][3] ~^ image[4][8])} + {7'd0,(kernel[4][4] ~^ image[4][9])};
assign out_fmap[0][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][6])} + {7'd0,(kernel[0][1] ~^ image[0][7])} + {7'd0,(kernel[0][2] ~^ image[0][8])} + {7'd0,(kernel[0][3] ~^ image[0][9])} + {7'd0,(kernel[0][4] ~^ image[0][10])} + {7'd0,(kernel[1][0] ~^ image[1][6])} + {7'd0,(kernel[1][1] ~^ image[1][7])} + {7'd0,(kernel[1][2] ~^ image[1][8])} + {7'd0,(kernel[1][3] ~^ image[1][9])} + {7'd0,(kernel[1][4] ~^ image[1][10])} + {7'd0,(kernel[2][0] ~^ image[2][6])} + {7'd0,(kernel[2][1] ~^ image[2][7])} + {7'd0,(kernel[2][2] ~^ image[2][8])} + {7'd0,(kernel[2][3] ~^ image[2][9])} + {7'd0,(kernel[2][4] ~^ image[2][10])} + {7'd0,(kernel[3][0] ~^ image[3][6])} + {7'd0,(kernel[3][1] ~^ image[3][7])} + {7'd0,(kernel[3][2] ~^ image[3][8])} + {7'd0,(kernel[3][3] ~^ image[3][9])} + {7'd0,(kernel[3][4] ~^ image[3][10])} + {7'd0,(kernel[4][0] ~^ image[4][6])} + {7'd0,(kernel[4][1] ~^ image[4][7])} + {7'd0,(kernel[4][2] ~^ image[4][8])} + {7'd0,(kernel[4][3] ~^ image[4][9])} + {7'd0,(kernel[4][4] ~^ image[4][10])};
assign out_fmap[0][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][7])} + {7'd0,(kernel[0][1] ~^ image[0][8])} + {7'd0,(kernel[0][2] ~^ image[0][9])} + {7'd0,(kernel[0][3] ~^ image[0][10])} + {7'd0,(kernel[0][4] ~^ image[0][11])} + {7'd0,(kernel[1][0] ~^ image[1][7])} + {7'd0,(kernel[1][1] ~^ image[1][8])} + {7'd0,(kernel[1][2] ~^ image[1][9])} + {7'd0,(kernel[1][3] ~^ image[1][10])} + {7'd0,(kernel[1][4] ~^ image[1][11])} + {7'd0,(kernel[2][0] ~^ image[2][7])} + {7'd0,(kernel[2][1] ~^ image[2][8])} + {7'd0,(kernel[2][2] ~^ image[2][9])} + {7'd0,(kernel[2][3] ~^ image[2][10])} + {7'd0,(kernel[2][4] ~^ image[2][11])} + {7'd0,(kernel[3][0] ~^ image[3][7])} + {7'd0,(kernel[3][1] ~^ image[3][8])} + {7'd0,(kernel[3][2] ~^ image[3][9])} + {7'd0,(kernel[3][3] ~^ image[3][10])} + {7'd0,(kernel[3][4] ~^ image[3][11])} + {7'd0,(kernel[4][0] ~^ image[4][7])} + {7'd0,(kernel[4][1] ~^ image[4][8])} + {7'd0,(kernel[4][2] ~^ image[4][9])} + {7'd0,(kernel[4][3] ~^ image[4][10])} + {7'd0,(kernel[4][4] ~^ image[4][11])};
assign out_fmap[1][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][0])} + {7'd0,(kernel[0][1] ~^ image[1][1])} + {7'd0,(kernel[0][2] ~^ image[1][2])} + {7'd0,(kernel[0][3] ~^ image[1][3])} + {7'd0,(kernel[0][4] ~^ image[1][4])} + {7'd0,(kernel[1][0] ~^ image[2][0])} + {7'd0,(kernel[1][1] ~^ image[2][1])} + {7'd0,(kernel[1][2] ~^ image[2][2])} + {7'd0,(kernel[1][3] ~^ image[2][3])} + {7'd0,(kernel[1][4] ~^ image[2][4])} + {7'd0,(kernel[2][0] ~^ image[3][0])} + {7'd0,(kernel[2][1] ~^ image[3][1])} + {7'd0,(kernel[2][2] ~^ image[3][2])} + {7'd0,(kernel[2][3] ~^ image[3][3])} + {7'd0,(kernel[2][4] ~^ image[3][4])} + {7'd0,(kernel[3][0] ~^ image[4][0])} + {7'd0,(kernel[3][1] ~^ image[4][1])} + {7'd0,(kernel[3][2] ~^ image[4][2])} + {7'd0,(kernel[3][3] ~^ image[4][3])} + {7'd0,(kernel[3][4] ~^ image[4][4])} + {7'd0,(kernel[4][0] ~^ image[5][0])} + {7'd0,(kernel[4][1] ~^ image[5][1])} + {7'd0,(kernel[4][2] ~^ image[5][2])} + {7'd0,(kernel[4][3] ~^ image[5][3])} + {7'd0,(kernel[4][4] ~^ image[5][4])};
assign out_fmap[1][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][1])} + {7'd0,(kernel[0][1] ~^ image[1][2])} + {7'd0,(kernel[0][2] ~^ image[1][3])} + {7'd0,(kernel[0][3] ~^ image[1][4])} + {7'd0,(kernel[0][4] ~^ image[1][5])} + {7'd0,(kernel[1][0] ~^ image[2][1])} + {7'd0,(kernel[1][1] ~^ image[2][2])} + {7'd0,(kernel[1][2] ~^ image[2][3])} + {7'd0,(kernel[1][3] ~^ image[2][4])} + {7'd0,(kernel[1][4] ~^ image[2][5])} + {7'd0,(kernel[2][0] ~^ image[3][1])} + {7'd0,(kernel[2][1] ~^ image[3][2])} + {7'd0,(kernel[2][2] ~^ image[3][3])} + {7'd0,(kernel[2][3] ~^ image[3][4])} + {7'd0,(kernel[2][4] ~^ image[3][5])} + {7'd0,(kernel[3][0] ~^ image[4][1])} + {7'd0,(kernel[3][1] ~^ image[4][2])} + {7'd0,(kernel[3][2] ~^ image[4][3])} + {7'd0,(kernel[3][3] ~^ image[4][4])} + {7'd0,(kernel[3][4] ~^ image[4][5])} + {7'd0,(kernel[4][0] ~^ image[5][1])} + {7'd0,(kernel[4][1] ~^ image[5][2])} + {7'd0,(kernel[4][2] ~^ image[5][3])} + {7'd0,(kernel[4][3] ~^ image[5][4])} + {7'd0,(kernel[4][4] ~^ image[5][5])};
assign out_fmap[1][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][2])} + {7'd0,(kernel[0][1] ~^ image[1][3])} + {7'd0,(kernel[0][2] ~^ image[1][4])} + {7'd0,(kernel[0][3] ~^ image[1][5])} + {7'd0,(kernel[0][4] ~^ image[1][6])} + {7'd0,(kernel[1][0] ~^ image[2][2])} + {7'd0,(kernel[1][1] ~^ image[2][3])} + {7'd0,(kernel[1][2] ~^ image[2][4])} + {7'd0,(kernel[1][3] ~^ image[2][5])} + {7'd0,(kernel[1][4] ~^ image[2][6])} + {7'd0,(kernel[2][0] ~^ image[3][2])} + {7'd0,(kernel[2][1] ~^ image[3][3])} + {7'd0,(kernel[2][2] ~^ image[3][4])} + {7'd0,(kernel[2][3] ~^ image[3][5])} + {7'd0,(kernel[2][4] ~^ image[3][6])} + {7'd0,(kernel[3][0] ~^ image[4][2])} + {7'd0,(kernel[3][1] ~^ image[4][3])} + {7'd0,(kernel[3][2] ~^ image[4][4])} + {7'd0,(kernel[3][3] ~^ image[4][5])} + {7'd0,(kernel[3][4] ~^ image[4][6])} + {7'd0,(kernel[4][0] ~^ image[5][2])} + {7'd0,(kernel[4][1] ~^ image[5][3])} + {7'd0,(kernel[4][2] ~^ image[5][4])} + {7'd0,(kernel[4][3] ~^ image[5][5])} + {7'd0,(kernel[4][4] ~^ image[5][6])};
assign out_fmap[1][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][3])} + {7'd0,(kernel[0][1] ~^ image[1][4])} + {7'd0,(kernel[0][2] ~^ image[1][5])} + {7'd0,(kernel[0][3] ~^ image[1][6])} + {7'd0,(kernel[0][4] ~^ image[1][7])} + {7'd0,(kernel[1][0] ~^ image[2][3])} + {7'd0,(kernel[1][1] ~^ image[2][4])} + {7'd0,(kernel[1][2] ~^ image[2][5])} + {7'd0,(kernel[1][3] ~^ image[2][6])} + {7'd0,(kernel[1][4] ~^ image[2][7])} + {7'd0,(kernel[2][0] ~^ image[3][3])} + {7'd0,(kernel[2][1] ~^ image[3][4])} + {7'd0,(kernel[2][2] ~^ image[3][5])} + {7'd0,(kernel[2][3] ~^ image[3][6])} + {7'd0,(kernel[2][4] ~^ image[3][7])} + {7'd0,(kernel[3][0] ~^ image[4][3])} + {7'd0,(kernel[3][1] ~^ image[4][4])} + {7'd0,(kernel[3][2] ~^ image[4][5])} + {7'd0,(kernel[3][3] ~^ image[4][6])} + {7'd0,(kernel[3][4] ~^ image[4][7])} + {7'd0,(kernel[4][0] ~^ image[5][3])} + {7'd0,(kernel[4][1] ~^ image[5][4])} + {7'd0,(kernel[4][2] ~^ image[5][5])} + {7'd0,(kernel[4][3] ~^ image[5][6])} + {7'd0,(kernel[4][4] ~^ image[5][7])};
assign out_fmap[1][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][4])} + {7'd0,(kernel[0][1] ~^ image[1][5])} + {7'd0,(kernel[0][2] ~^ image[1][6])} + {7'd0,(kernel[0][3] ~^ image[1][7])} + {7'd0,(kernel[0][4] ~^ image[1][8])} + {7'd0,(kernel[1][0] ~^ image[2][4])} + {7'd0,(kernel[1][1] ~^ image[2][5])} + {7'd0,(kernel[1][2] ~^ image[2][6])} + {7'd0,(kernel[1][3] ~^ image[2][7])} + {7'd0,(kernel[1][4] ~^ image[2][8])} + {7'd0,(kernel[2][0] ~^ image[3][4])} + {7'd0,(kernel[2][1] ~^ image[3][5])} + {7'd0,(kernel[2][2] ~^ image[3][6])} + {7'd0,(kernel[2][3] ~^ image[3][7])} + {7'd0,(kernel[2][4] ~^ image[3][8])} + {7'd0,(kernel[3][0] ~^ image[4][4])} + {7'd0,(kernel[3][1] ~^ image[4][5])} + {7'd0,(kernel[3][2] ~^ image[4][6])} + {7'd0,(kernel[3][3] ~^ image[4][7])} + {7'd0,(kernel[3][4] ~^ image[4][8])} + {7'd0,(kernel[4][0] ~^ image[5][4])} + {7'd0,(kernel[4][1] ~^ image[5][5])} + {7'd0,(kernel[4][2] ~^ image[5][6])} + {7'd0,(kernel[4][3] ~^ image[5][7])} + {7'd0,(kernel[4][4] ~^ image[5][8])};
assign out_fmap[1][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][5])} + {7'd0,(kernel[0][1] ~^ image[1][6])} + {7'd0,(kernel[0][2] ~^ image[1][7])} + {7'd0,(kernel[0][3] ~^ image[1][8])} + {7'd0,(kernel[0][4] ~^ image[1][9])} + {7'd0,(kernel[1][0] ~^ image[2][5])} + {7'd0,(kernel[1][1] ~^ image[2][6])} + {7'd0,(kernel[1][2] ~^ image[2][7])} + {7'd0,(kernel[1][3] ~^ image[2][8])} + {7'd0,(kernel[1][4] ~^ image[2][9])} + {7'd0,(kernel[2][0] ~^ image[3][5])} + {7'd0,(kernel[2][1] ~^ image[3][6])} + {7'd0,(kernel[2][2] ~^ image[3][7])} + {7'd0,(kernel[2][3] ~^ image[3][8])} + {7'd0,(kernel[2][4] ~^ image[3][9])} + {7'd0,(kernel[3][0] ~^ image[4][5])} + {7'd0,(kernel[3][1] ~^ image[4][6])} + {7'd0,(kernel[3][2] ~^ image[4][7])} + {7'd0,(kernel[3][3] ~^ image[4][8])} + {7'd0,(kernel[3][4] ~^ image[4][9])} + {7'd0,(kernel[4][0] ~^ image[5][5])} + {7'd0,(kernel[4][1] ~^ image[5][6])} + {7'd0,(kernel[4][2] ~^ image[5][7])} + {7'd0,(kernel[4][3] ~^ image[5][8])} + {7'd0,(kernel[4][4] ~^ image[5][9])};
assign out_fmap[1][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][6])} + {7'd0,(kernel[0][1] ~^ image[1][7])} + {7'd0,(kernel[0][2] ~^ image[1][8])} + {7'd0,(kernel[0][3] ~^ image[1][9])} + {7'd0,(kernel[0][4] ~^ image[1][10])} + {7'd0,(kernel[1][0] ~^ image[2][6])} + {7'd0,(kernel[1][1] ~^ image[2][7])} + {7'd0,(kernel[1][2] ~^ image[2][8])} + {7'd0,(kernel[1][3] ~^ image[2][9])} + {7'd0,(kernel[1][4] ~^ image[2][10])} + {7'd0,(kernel[2][0] ~^ image[3][6])} + {7'd0,(kernel[2][1] ~^ image[3][7])} + {7'd0,(kernel[2][2] ~^ image[3][8])} + {7'd0,(kernel[2][3] ~^ image[3][9])} + {7'd0,(kernel[2][4] ~^ image[3][10])} + {7'd0,(kernel[3][0] ~^ image[4][6])} + {7'd0,(kernel[3][1] ~^ image[4][7])} + {7'd0,(kernel[3][2] ~^ image[4][8])} + {7'd0,(kernel[3][3] ~^ image[4][9])} + {7'd0,(kernel[3][4] ~^ image[4][10])} + {7'd0,(kernel[4][0] ~^ image[5][6])} + {7'd0,(kernel[4][1] ~^ image[5][7])} + {7'd0,(kernel[4][2] ~^ image[5][8])} + {7'd0,(kernel[4][3] ~^ image[5][9])} + {7'd0,(kernel[4][4] ~^ image[5][10])};
assign out_fmap[1][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][7])} + {7'd0,(kernel[0][1] ~^ image[1][8])} + {7'd0,(kernel[0][2] ~^ image[1][9])} + {7'd0,(kernel[0][3] ~^ image[1][10])} + {7'd0,(kernel[0][4] ~^ image[1][11])} + {7'd0,(kernel[1][0] ~^ image[2][7])} + {7'd0,(kernel[1][1] ~^ image[2][8])} + {7'd0,(kernel[1][2] ~^ image[2][9])} + {7'd0,(kernel[1][3] ~^ image[2][10])} + {7'd0,(kernel[1][4] ~^ image[2][11])} + {7'd0,(kernel[2][0] ~^ image[3][7])} + {7'd0,(kernel[2][1] ~^ image[3][8])} + {7'd0,(kernel[2][2] ~^ image[3][9])} + {7'd0,(kernel[2][3] ~^ image[3][10])} + {7'd0,(kernel[2][4] ~^ image[3][11])} + {7'd0,(kernel[3][0] ~^ image[4][7])} + {7'd0,(kernel[3][1] ~^ image[4][8])} + {7'd0,(kernel[3][2] ~^ image[4][9])} + {7'd0,(kernel[3][3] ~^ image[4][10])} + {7'd0,(kernel[3][4] ~^ image[4][11])} + {7'd0,(kernel[4][0] ~^ image[5][7])} + {7'd0,(kernel[4][1] ~^ image[5][8])} + {7'd0,(kernel[4][2] ~^ image[5][9])} + {7'd0,(kernel[4][3] ~^ image[5][10])} + {7'd0,(kernel[4][4] ~^ image[5][11])};
assign out_fmap[2][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][0])} + {7'd0,(kernel[0][1] ~^ image[2][1])} + {7'd0,(kernel[0][2] ~^ image[2][2])} + {7'd0,(kernel[0][3] ~^ image[2][3])} + {7'd0,(kernel[0][4] ~^ image[2][4])} + {7'd0,(kernel[1][0] ~^ image[3][0])} + {7'd0,(kernel[1][1] ~^ image[3][1])} + {7'd0,(kernel[1][2] ~^ image[3][2])} + {7'd0,(kernel[1][3] ~^ image[3][3])} + {7'd0,(kernel[1][4] ~^ image[3][4])} + {7'd0,(kernel[2][0] ~^ image[4][0])} + {7'd0,(kernel[2][1] ~^ image[4][1])} + {7'd0,(kernel[2][2] ~^ image[4][2])} + {7'd0,(kernel[2][3] ~^ image[4][3])} + {7'd0,(kernel[2][4] ~^ image[4][4])} + {7'd0,(kernel[3][0] ~^ image[5][0])} + {7'd0,(kernel[3][1] ~^ image[5][1])} + {7'd0,(kernel[3][2] ~^ image[5][2])} + {7'd0,(kernel[3][3] ~^ image[5][3])} + {7'd0,(kernel[3][4] ~^ image[5][4])} + {7'd0,(kernel[4][0] ~^ image[6][0])} + {7'd0,(kernel[4][1] ~^ image[6][1])} + {7'd0,(kernel[4][2] ~^ image[6][2])} + {7'd0,(kernel[4][3] ~^ image[6][3])} + {7'd0,(kernel[4][4] ~^ image[6][4])};
assign out_fmap[2][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][1])} + {7'd0,(kernel[0][1] ~^ image[2][2])} + {7'd0,(kernel[0][2] ~^ image[2][3])} + {7'd0,(kernel[0][3] ~^ image[2][4])} + {7'd0,(kernel[0][4] ~^ image[2][5])} + {7'd0,(kernel[1][0] ~^ image[3][1])} + {7'd0,(kernel[1][1] ~^ image[3][2])} + {7'd0,(kernel[1][2] ~^ image[3][3])} + {7'd0,(kernel[1][3] ~^ image[3][4])} + {7'd0,(kernel[1][4] ~^ image[3][5])} + {7'd0,(kernel[2][0] ~^ image[4][1])} + {7'd0,(kernel[2][1] ~^ image[4][2])} + {7'd0,(kernel[2][2] ~^ image[4][3])} + {7'd0,(kernel[2][3] ~^ image[4][4])} + {7'd0,(kernel[2][4] ~^ image[4][5])} + {7'd0,(kernel[3][0] ~^ image[5][1])} + {7'd0,(kernel[3][1] ~^ image[5][2])} + {7'd0,(kernel[3][2] ~^ image[5][3])} + {7'd0,(kernel[3][3] ~^ image[5][4])} + {7'd0,(kernel[3][4] ~^ image[5][5])} + {7'd0,(kernel[4][0] ~^ image[6][1])} + {7'd0,(kernel[4][1] ~^ image[6][2])} + {7'd0,(kernel[4][2] ~^ image[6][3])} + {7'd0,(kernel[4][3] ~^ image[6][4])} + {7'd0,(kernel[4][4] ~^ image[6][5])};
assign out_fmap[2][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][2])} + {7'd0,(kernel[0][1] ~^ image[2][3])} + {7'd0,(kernel[0][2] ~^ image[2][4])} + {7'd0,(kernel[0][3] ~^ image[2][5])} + {7'd0,(kernel[0][4] ~^ image[2][6])} + {7'd0,(kernel[1][0] ~^ image[3][2])} + {7'd0,(kernel[1][1] ~^ image[3][3])} + {7'd0,(kernel[1][2] ~^ image[3][4])} + {7'd0,(kernel[1][3] ~^ image[3][5])} + {7'd0,(kernel[1][4] ~^ image[3][6])} + {7'd0,(kernel[2][0] ~^ image[4][2])} + {7'd0,(kernel[2][1] ~^ image[4][3])} + {7'd0,(kernel[2][2] ~^ image[4][4])} + {7'd0,(kernel[2][3] ~^ image[4][5])} + {7'd0,(kernel[2][4] ~^ image[4][6])} + {7'd0,(kernel[3][0] ~^ image[5][2])} + {7'd0,(kernel[3][1] ~^ image[5][3])} + {7'd0,(kernel[3][2] ~^ image[5][4])} + {7'd0,(kernel[3][3] ~^ image[5][5])} + {7'd0,(kernel[3][4] ~^ image[5][6])} + {7'd0,(kernel[4][0] ~^ image[6][2])} + {7'd0,(kernel[4][1] ~^ image[6][3])} + {7'd0,(kernel[4][2] ~^ image[6][4])} + {7'd0,(kernel[4][3] ~^ image[6][5])} + {7'd0,(kernel[4][4] ~^ image[6][6])};
assign out_fmap[2][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][3])} + {7'd0,(kernel[0][1] ~^ image[2][4])} + {7'd0,(kernel[0][2] ~^ image[2][5])} + {7'd0,(kernel[0][3] ~^ image[2][6])} + {7'd0,(kernel[0][4] ~^ image[2][7])} + {7'd0,(kernel[1][0] ~^ image[3][3])} + {7'd0,(kernel[1][1] ~^ image[3][4])} + {7'd0,(kernel[1][2] ~^ image[3][5])} + {7'd0,(kernel[1][3] ~^ image[3][6])} + {7'd0,(kernel[1][4] ~^ image[3][7])} + {7'd0,(kernel[2][0] ~^ image[4][3])} + {7'd0,(kernel[2][1] ~^ image[4][4])} + {7'd0,(kernel[2][2] ~^ image[4][5])} + {7'd0,(kernel[2][3] ~^ image[4][6])} + {7'd0,(kernel[2][4] ~^ image[4][7])} + {7'd0,(kernel[3][0] ~^ image[5][3])} + {7'd0,(kernel[3][1] ~^ image[5][4])} + {7'd0,(kernel[3][2] ~^ image[5][5])} + {7'd0,(kernel[3][3] ~^ image[5][6])} + {7'd0,(kernel[3][4] ~^ image[5][7])} + {7'd0,(kernel[4][0] ~^ image[6][3])} + {7'd0,(kernel[4][1] ~^ image[6][4])} + {7'd0,(kernel[4][2] ~^ image[6][5])} + {7'd0,(kernel[4][3] ~^ image[6][6])} + {7'd0,(kernel[4][4] ~^ image[6][7])};
assign out_fmap[2][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][4])} + {7'd0,(kernel[0][1] ~^ image[2][5])} + {7'd0,(kernel[0][2] ~^ image[2][6])} + {7'd0,(kernel[0][3] ~^ image[2][7])} + {7'd0,(kernel[0][4] ~^ image[2][8])} + {7'd0,(kernel[1][0] ~^ image[3][4])} + {7'd0,(kernel[1][1] ~^ image[3][5])} + {7'd0,(kernel[1][2] ~^ image[3][6])} + {7'd0,(kernel[1][3] ~^ image[3][7])} + {7'd0,(kernel[1][4] ~^ image[3][8])} + {7'd0,(kernel[2][0] ~^ image[4][4])} + {7'd0,(kernel[2][1] ~^ image[4][5])} + {7'd0,(kernel[2][2] ~^ image[4][6])} + {7'd0,(kernel[2][3] ~^ image[4][7])} + {7'd0,(kernel[2][4] ~^ image[4][8])} + {7'd0,(kernel[3][0] ~^ image[5][4])} + {7'd0,(kernel[3][1] ~^ image[5][5])} + {7'd0,(kernel[3][2] ~^ image[5][6])} + {7'd0,(kernel[3][3] ~^ image[5][7])} + {7'd0,(kernel[3][4] ~^ image[5][8])} + {7'd0,(kernel[4][0] ~^ image[6][4])} + {7'd0,(kernel[4][1] ~^ image[6][5])} + {7'd0,(kernel[4][2] ~^ image[6][6])} + {7'd0,(kernel[4][3] ~^ image[6][7])} + {7'd0,(kernel[4][4] ~^ image[6][8])};
assign out_fmap[2][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][5])} + {7'd0,(kernel[0][1] ~^ image[2][6])} + {7'd0,(kernel[0][2] ~^ image[2][7])} + {7'd0,(kernel[0][3] ~^ image[2][8])} + {7'd0,(kernel[0][4] ~^ image[2][9])} + {7'd0,(kernel[1][0] ~^ image[3][5])} + {7'd0,(kernel[1][1] ~^ image[3][6])} + {7'd0,(kernel[1][2] ~^ image[3][7])} + {7'd0,(kernel[1][3] ~^ image[3][8])} + {7'd0,(kernel[1][4] ~^ image[3][9])} + {7'd0,(kernel[2][0] ~^ image[4][5])} + {7'd0,(kernel[2][1] ~^ image[4][6])} + {7'd0,(kernel[2][2] ~^ image[4][7])} + {7'd0,(kernel[2][3] ~^ image[4][8])} + {7'd0,(kernel[2][4] ~^ image[4][9])} + {7'd0,(kernel[3][0] ~^ image[5][5])} + {7'd0,(kernel[3][1] ~^ image[5][6])} + {7'd0,(kernel[3][2] ~^ image[5][7])} + {7'd0,(kernel[3][3] ~^ image[5][8])} + {7'd0,(kernel[3][4] ~^ image[5][9])} + {7'd0,(kernel[4][0] ~^ image[6][5])} + {7'd0,(kernel[4][1] ~^ image[6][6])} + {7'd0,(kernel[4][2] ~^ image[6][7])} + {7'd0,(kernel[4][3] ~^ image[6][8])} + {7'd0,(kernel[4][4] ~^ image[6][9])};
assign out_fmap[2][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][6])} + {7'd0,(kernel[0][1] ~^ image[2][7])} + {7'd0,(kernel[0][2] ~^ image[2][8])} + {7'd0,(kernel[0][3] ~^ image[2][9])} + {7'd0,(kernel[0][4] ~^ image[2][10])} + {7'd0,(kernel[1][0] ~^ image[3][6])} + {7'd0,(kernel[1][1] ~^ image[3][7])} + {7'd0,(kernel[1][2] ~^ image[3][8])} + {7'd0,(kernel[1][3] ~^ image[3][9])} + {7'd0,(kernel[1][4] ~^ image[3][10])} + {7'd0,(kernel[2][0] ~^ image[4][6])} + {7'd0,(kernel[2][1] ~^ image[4][7])} + {7'd0,(kernel[2][2] ~^ image[4][8])} + {7'd0,(kernel[2][3] ~^ image[4][9])} + {7'd0,(kernel[2][4] ~^ image[4][10])} + {7'd0,(kernel[3][0] ~^ image[5][6])} + {7'd0,(kernel[3][1] ~^ image[5][7])} + {7'd0,(kernel[3][2] ~^ image[5][8])} + {7'd0,(kernel[3][3] ~^ image[5][9])} + {7'd0,(kernel[3][4] ~^ image[5][10])} + {7'd0,(kernel[4][0] ~^ image[6][6])} + {7'd0,(kernel[4][1] ~^ image[6][7])} + {7'd0,(kernel[4][2] ~^ image[6][8])} + {7'd0,(kernel[4][3] ~^ image[6][9])} + {7'd0,(kernel[4][4] ~^ image[6][10])};
assign out_fmap[2][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][7])} + {7'd0,(kernel[0][1] ~^ image[2][8])} + {7'd0,(kernel[0][2] ~^ image[2][9])} + {7'd0,(kernel[0][3] ~^ image[2][10])} + {7'd0,(kernel[0][4] ~^ image[2][11])} + {7'd0,(kernel[1][0] ~^ image[3][7])} + {7'd0,(kernel[1][1] ~^ image[3][8])} + {7'd0,(kernel[1][2] ~^ image[3][9])} + {7'd0,(kernel[1][3] ~^ image[3][10])} + {7'd0,(kernel[1][4] ~^ image[3][11])} + {7'd0,(kernel[2][0] ~^ image[4][7])} + {7'd0,(kernel[2][1] ~^ image[4][8])} + {7'd0,(kernel[2][2] ~^ image[4][9])} + {7'd0,(kernel[2][3] ~^ image[4][10])} + {7'd0,(kernel[2][4] ~^ image[4][11])} + {7'd0,(kernel[3][0] ~^ image[5][7])} + {7'd0,(kernel[3][1] ~^ image[5][8])} + {7'd0,(kernel[3][2] ~^ image[5][9])} + {7'd0,(kernel[3][3] ~^ image[5][10])} + {7'd0,(kernel[3][4] ~^ image[5][11])} + {7'd0,(kernel[4][0] ~^ image[6][7])} + {7'd0,(kernel[4][1] ~^ image[6][8])} + {7'd0,(kernel[4][2] ~^ image[6][9])} + {7'd0,(kernel[4][3] ~^ image[6][10])} + {7'd0,(kernel[4][4] ~^ image[6][11])};
assign out_fmap[3][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][0])} + {7'd0,(kernel[0][1] ~^ image[3][1])} + {7'd0,(kernel[0][2] ~^ image[3][2])} + {7'd0,(kernel[0][3] ~^ image[3][3])} + {7'd0,(kernel[0][4] ~^ image[3][4])} + {7'd0,(kernel[1][0] ~^ image[4][0])} + {7'd0,(kernel[1][1] ~^ image[4][1])} + {7'd0,(kernel[1][2] ~^ image[4][2])} + {7'd0,(kernel[1][3] ~^ image[4][3])} + {7'd0,(kernel[1][4] ~^ image[4][4])} + {7'd0,(kernel[2][0] ~^ image[5][0])} + {7'd0,(kernel[2][1] ~^ image[5][1])} + {7'd0,(kernel[2][2] ~^ image[5][2])} + {7'd0,(kernel[2][3] ~^ image[5][3])} + {7'd0,(kernel[2][4] ~^ image[5][4])} + {7'd0,(kernel[3][0] ~^ image[6][0])} + {7'd0,(kernel[3][1] ~^ image[6][1])} + {7'd0,(kernel[3][2] ~^ image[6][2])} + {7'd0,(kernel[3][3] ~^ image[6][3])} + {7'd0,(kernel[3][4] ~^ image[6][4])} + {7'd0,(kernel[4][0] ~^ image[7][0])} + {7'd0,(kernel[4][1] ~^ image[7][1])} + {7'd0,(kernel[4][2] ~^ image[7][2])} + {7'd0,(kernel[4][3] ~^ image[7][3])} + {7'd0,(kernel[4][4] ~^ image[7][4])};
assign out_fmap[3][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][1])} + {7'd0,(kernel[0][1] ~^ image[3][2])} + {7'd0,(kernel[0][2] ~^ image[3][3])} + {7'd0,(kernel[0][3] ~^ image[3][4])} + {7'd0,(kernel[0][4] ~^ image[3][5])} + {7'd0,(kernel[1][0] ~^ image[4][1])} + {7'd0,(kernel[1][1] ~^ image[4][2])} + {7'd0,(kernel[1][2] ~^ image[4][3])} + {7'd0,(kernel[1][3] ~^ image[4][4])} + {7'd0,(kernel[1][4] ~^ image[4][5])} + {7'd0,(kernel[2][0] ~^ image[5][1])} + {7'd0,(kernel[2][1] ~^ image[5][2])} + {7'd0,(kernel[2][2] ~^ image[5][3])} + {7'd0,(kernel[2][3] ~^ image[5][4])} + {7'd0,(kernel[2][4] ~^ image[5][5])} + {7'd0,(kernel[3][0] ~^ image[6][1])} + {7'd0,(kernel[3][1] ~^ image[6][2])} + {7'd0,(kernel[3][2] ~^ image[6][3])} + {7'd0,(kernel[3][3] ~^ image[6][4])} + {7'd0,(kernel[3][4] ~^ image[6][5])} + {7'd0,(kernel[4][0] ~^ image[7][1])} + {7'd0,(kernel[4][1] ~^ image[7][2])} + {7'd0,(kernel[4][2] ~^ image[7][3])} + {7'd0,(kernel[4][3] ~^ image[7][4])} + {7'd0,(kernel[4][4] ~^ image[7][5])};
assign out_fmap[3][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][2])} + {7'd0,(kernel[0][1] ~^ image[3][3])} + {7'd0,(kernel[0][2] ~^ image[3][4])} + {7'd0,(kernel[0][3] ~^ image[3][5])} + {7'd0,(kernel[0][4] ~^ image[3][6])} + {7'd0,(kernel[1][0] ~^ image[4][2])} + {7'd0,(kernel[1][1] ~^ image[4][3])} + {7'd0,(kernel[1][2] ~^ image[4][4])} + {7'd0,(kernel[1][3] ~^ image[4][5])} + {7'd0,(kernel[1][4] ~^ image[4][6])} + {7'd0,(kernel[2][0] ~^ image[5][2])} + {7'd0,(kernel[2][1] ~^ image[5][3])} + {7'd0,(kernel[2][2] ~^ image[5][4])} + {7'd0,(kernel[2][3] ~^ image[5][5])} + {7'd0,(kernel[2][4] ~^ image[5][6])} + {7'd0,(kernel[3][0] ~^ image[6][2])} + {7'd0,(kernel[3][1] ~^ image[6][3])} + {7'd0,(kernel[3][2] ~^ image[6][4])} + {7'd0,(kernel[3][3] ~^ image[6][5])} + {7'd0,(kernel[3][4] ~^ image[6][6])} + {7'd0,(kernel[4][0] ~^ image[7][2])} + {7'd0,(kernel[4][1] ~^ image[7][3])} + {7'd0,(kernel[4][2] ~^ image[7][4])} + {7'd0,(kernel[4][3] ~^ image[7][5])} + {7'd0,(kernel[4][4] ~^ image[7][6])};
assign out_fmap[3][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][3])} + {7'd0,(kernel[0][1] ~^ image[3][4])} + {7'd0,(kernel[0][2] ~^ image[3][5])} + {7'd0,(kernel[0][3] ~^ image[3][6])} + {7'd0,(kernel[0][4] ~^ image[3][7])} + {7'd0,(kernel[1][0] ~^ image[4][3])} + {7'd0,(kernel[1][1] ~^ image[4][4])} + {7'd0,(kernel[1][2] ~^ image[4][5])} + {7'd0,(kernel[1][3] ~^ image[4][6])} + {7'd0,(kernel[1][4] ~^ image[4][7])} + {7'd0,(kernel[2][0] ~^ image[5][3])} + {7'd0,(kernel[2][1] ~^ image[5][4])} + {7'd0,(kernel[2][2] ~^ image[5][5])} + {7'd0,(kernel[2][3] ~^ image[5][6])} + {7'd0,(kernel[2][4] ~^ image[5][7])} + {7'd0,(kernel[3][0] ~^ image[6][3])} + {7'd0,(kernel[3][1] ~^ image[6][4])} + {7'd0,(kernel[3][2] ~^ image[6][5])} + {7'd0,(kernel[3][3] ~^ image[6][6])} + {7'd0,(kernel[3][4] ~^ image[6][7])} + {7'd0,(kernel[4][0] ~^ image[7][3])} + {7'd0,(kernel[4][1] ~^ image[7][4])} + {7'd0,(kernel[4][2] ~^ image[7][5])} + {7'd0,(kernel[4][3] ~^ image[7][6])} + {7'd0,(kernel[4][4] ~^ image[7][7])};
assign out_fmap[3][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][4])} + {7'd0,(kernel[0][1] ~^ image[3][5])} + {7'd0,(kernel[0][2] ~^ image[3][6])} + {7'd0,(kernel[0][3] ~^ image[3][7])} + {7'd0,(kernel[0][4] ~^ image[3][8])} + {7'd0,(kernel[1][0] ~^ image[4][4])} + {7'd0,(kernel[1][1] ~^ image[4][5])} + {7'd0,(kernel[1][2] ~^ image[4][6])} + {7'd0,(kernel[1][3] ~^ image[4][7])} + {7'd0,(kernel[1][4] ~^ image[4][8])} + {7'd0,(kernel[2][0] ~^ image[5][4])} + {7'd0,(kernel[2][1] ~^ image[5][5])} + {7'd0,(kernel[2][2] ~^ image[5][6])} + {7'd0,(kernel[2][3] ~^ image[5][7])} + {7'd0,(kernel[2][4] ~^ image[5][8])} + {7'd0,(kernel[3][0] ~^ image[6][4])} + {7'd0,(kernel[3][1] ~^ image[6][5])} + {7'd0,(kernel[3][2] ~^ image[6][6])} + {7'd0,(kernel[3][3] ~^ image[6][7])} + {7'd0,(kernel[3][4] ~^ image[6][8])} + {7'd0,(kernel[4][0] ~^ image[7][4])} + {7'd0,(kernel[4][1] ~^ image[7][5])} + {7'd0,(kernel[4][2] ~^ image[7][6])} + {7'd0,(kernel[4][3] ~^ image[7][7])} + {7'd0,(kernel[4][4] ~^ image[7][8])};
assign out_fmap[3][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][5])} + {7'd0,(kernel[0][1] ~^ image[3][6])} + {7'd0,(kernel[0][2] ~^ image[3][7])} + {7'd0,(kernel[0][3] ~^ image[3][8])} + {7'd0,(kernel[0][4] ~^ image[3][9])} + {7'd0,(kernel[1][0] ~^ image[4][5])} + {7'd0,(kernel[1][1] ~^ image[4][6])} + {7'd0,(kernel[1][2] ~^ image[4][7])} + {7'd0,(kernel[1][3] ~^ image[4][8])} + {7'd0,(kernel[1][4] ~^ image[4][9])} + {7'd0,(kernel[2][0] ~^ image[5][5])} + {7'd0,(kernel[2][1] ~^ image[5][6])} + {7'd0,(kernel[2][2] ~^ image[5][7])} + {7'd0,(kernel[2][3] ~^ image[5][8])} + {7'd0,(kernel[2][4] ~^ image[5][9])} + {7'd0,(kernel[3][0] ~^ image[6][5])} + {7'd0,(kernel[3][1] ~^ image[6][6])} + {7'd0,(kernel[3][2] ~^ image[6][7])} + {7'd0,(kernel[3][3] ~^ image[6][8])} + {7'd0,(kernel[3][4] ~^ image[6][9])} + {7'd0,(kernel[4][0] ~^ image[7][5])} + {7'd0,(kernel[4][1] ~^ image[7][6])} + {7'd0,(kernel[4][2] ~^ image[7][7])} + {7'd0,(kernel[4][3] ~^ image[7][8])} + {7'd0,(kernel[4][4] ~^ image[7][9])};
assign out_fmap[3][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][6])} + {7'd0,(kernel[0][1] ~^ image[3][7])} + {7'd0,(kernel[0][2] ~^ image[3][8])} + {7'd0,(kernel[0][3] ~^ image[3][9])} + {7'd0,(kernel[0][4] ~^ image[3][10])} + {7'd0,(kernel[1][0] ~^ image[4][6])} + {7'd0,(kernel[1][1] ~^ image[4][7])} + {7'd0,(kernel[1][2] ~^ image[4][8])} + {7'd0,(kernel[1][3] ~^ image[4][9])} + {7'd0,(kernel[1][4] ~^ image[4][10])} + {7'd0,(kernel[2][0] ~^ image[5][6])} + {7'd0,(kernel[2][1] ~^ image[5][7])} + {7'd0,(kernel[2][2] ~^ image[5][8])} + {7'd0,(kernel[2][3] ~^ image[5][9])} + {7'd0,(kernel[2][4] ~^ image[5][10])} + {7'd0,(kernel[3][0] ~^ image[6][6])} + {7'd0,(kernel[3][1] ~^ image[6][7])} + {7'd0,(kernel[3][2] ~^ image[6][8])} + {7'd0,(kernel[3][3] ~^ image[6][9])} + {7'd0,(kernel[3][4] ~^ image[6][10])} + {7'd0,(kernel[4][0] ~^ image[7][6])} + {7'd0,(kernel[4][1] ~^ image[7][7])} + {7'd0,(kernel[4][2] ~^ image[7][8])} + {7'd0,(kernel[4][3] ~^ image[7][9])} + {7'd0,(kernel[4][4] ~^ image[7][10])};
assign out_fmap[3][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][7])} + {7'd0,(kernel[0][1] ~^ image[3][8])} + {7'd0,(kernel[0][2] ~^ image[3][9])} + {7'd0,(kernel[0][3] ~^ image[3][10])} + {7'd0,(kernel[0][4] ~^ image[3][11])} + {7'd0,(kernel[1][0] ~^ image[4][7])} + {7'd0,(kernel[1][1] ~^ image[4][8])} + {7'd0,(kernel[1][2] ~^ image[4][9])} + {7'd0,(kernel[1][3] ~^ image[4][10])} + {7'd0,(kernel[1][4] ~^ image[4][11])} + {7'd0,(kernel[2][0] ~^ image[5][7])} + {7'd0,(kernel[2][1] ~^ image[5][8])} + {7'd0,(kernel[2][2] ~^ image[5][9])} + {7'd0,(kernel[2][3] ~^ image[5][10])} + {7'd0,(kernel[2][4] ~^ image[5][11])} + {7'd0,(kernel[3][0] ~^ image[6][7])} + {7'd0,(kernel[3][1] ~^ image[6][8])} + {7'd0,(kernel[3][2] ~^ image[6][9])} + {7'd0,(kernel[3][3] ~^ image[6][10])} + {7'd0,(kernel[3][4] ~^ image[6][11])} + {7'd0,(kernel[4][0] ~^ image[7][7])} + {7'd0,(kernel[4][1] ~^ image[7][8])} + {7'd0,(kernel[4][2] ~^ image[7][9])} + {7'd0,(kernel[4][3] ~^ image[7][10])} + {7'd0,(kernel[4][4] ~^ image[7][11])};
assign out_fmap[4][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][0])} + {7'd0,(kernel[0][1] ~^ image[4][1])} + {7'd0,(kernel[0][2] ~^ image[4][2])} + {7'd0,(kernel[0][3] ~^ image[4][3])} + {7'd0,(kernel[0][4] ~^ image[4][4])} + {7'd0,(kernel[1][0] ~^ image[5][0])} + {7'd0,(kernel[1][1] ~^ image[5][1])} + {7'd0,(kernel[1][2] ~^ image[5][2])} + {7'd0,(kernel[1][3] ~^ image[5][3])} + {7'd0,(kernel[1][4] ~^ image[5][4])} + {7'd0,(kernel[2][0] ~^ image[6][0])} + {7'd0,(kernel[2][1] ~^ image[6][1])} + {7'd0,(kernel[2][2] ~^ image[6][2])} + {7'd0,(kernel[2][3] ~^ image[6][3])} + {7'd0,(kernel[2][4] ~^ image[6][4])} + {7'd0,(kernel[3][0] ~^ image[7][0])} + {7'd0,(kernel[3][1] ~^ image[7][1])} + {7'd0,(kernel[3][2] ~^ image[7][2])} + {7'd0,(kernel[3][3] ~^ image[7][3])} + {7'd0,(kernel[3][4] ~^ image[7][4])} + {7'd0,(kernel[4][0] ~^ image[8][0])} + {7'd0,(kernel[4][1] ~^ image[8][1])} + {7'd0,(kernel[4][2] ~^ image[8][2])} + {7'd0,(kernel[4][3] ~^ image[8][3])} + {7'd0,(kernel[4][4] ~^ image[8][4])};
assign out_fmap[4][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][1])} + {7'd0,(kernel[0][1] ~^ image[4][2])} + {7'd0,(kernel[0][2] ~^ image[4][3])} + {7'd0,(kernel[0][3] ~^ image[4][4])} + {7'd0,(kernel[0][4] ~^ image[4][5])} + {7'd0,(kernel[1][0] ~^ image[5][1])} + {7'd0,(kernel[1][1] ~^ image[5][2])} + {7'd0,(kernel[1][2] ~^ image[5][3])} + {7'd0,(kernel[1][3] ~^ image[5][4])} + {7'd0,(kernel[1][4] ~^ image[5][5])} + {7'd0,(kernel[2][0] ~^ image[6][1])} + {7'd0,(kernel[2][1] ~^ image[6][2])} + {7'd0,(kernel[2][2] ~^ image[6][3])} + {7'd0,(kernel[2][3] ~^ image[6][4])} + {7'd0,(kernel[2][4] ~^ image[6][5])} + {7'd0,(kernel[3][0] ~^ image[7][1])} + {7'd0,(kernel[3][1] ~^ image[7][2])} + {7'd0,(kernel[3][2] ~^ image[7][3])} + {7'd0,(kernel[3][3] ~^ image[7][4])} + {7'd0,(kernel[3][4] ~^ image[7][5])} + {7'd0,(kernel[4][0] ~^ image[8][1])} + {7'd0,(kernel[4][1] ~^ image[8][2])} + {7'd0,(kernel[4][2] ~^ image[8][3])} + {7'd0,(kernel[4][3] ~^ image[8][4])} + {7'd0,(kernel[4][4] ~^ image[8][5])};
assign out_fmap[4][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][2])} + {7'd0,(kernel[0][1] ~^ image[4][3])} + {7'd0,(kernel[0][2] ~^ image[4][4])} + {7'd0,(kernel[0][3] ~^ image[4][5])} + {7'd0,(kernel[0][4] ~^ image[4][6])} + {7'd0,(kernel[1][0] ~^ image[5][2])} + {7'd0,(kernel[1][1] ~^ image[5][3])} + {7'd0,(kernel[1][2] ~^ image[5][4])} + {7'd0,(kernel[1][3] ~^ image[5][5])} + {7'd0,(kernel[1][4] ~^ image[5][6])} + {7'd0,(kernel[2][0] ~^ image[6][2])} + {7'd0,(kernel[2][1] ~^ image[6][3])} + {7'd0,(kernel[2][2] ~^ image[6][4])} + {7'd0,(kernel[2][3] ~^ image[6][5])} + {7'd0,(kernel[2][4] ~^ image[6][6])} + {7'd0,(kernel[3][0] ~^ image[7][2])} + {7'd0,(kernel[3][1] ~^ image[7][3])} + {7'd0,(kernel[3][2] ~^ image[7][4])} + {7'd0,(kernel[3][3] ~^ image[7][5])} + {7'd0,(kernel[3][4] ~^ image[7][6])} + {7'd0,(kernel[4][0] ~^ image[8][2])} + {7'd0,(kernel[4][1] ~^ image[8][3])} + {7'd0,(kernel[4][2] ~^ image[8][4])} + {7'd0,(kernel[4][3] ~^ image[8][5])} + {7'd0,(kernel[4][4] ~^ image[8][6])};
assign out_fmap[4][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][3])} + {7'd0,(kernel[0][1] ~^ image[4][4])} + {7'd0,(kernel[0][2] ~^ image[4][5])} + {7'd0,(kernel[0][3] ~^ image[4][6])} + {7'd0,(kernel[0][4] ~^ image[4][7])} + {7'd0,(kernel[1][0] ~^ image[5][3])} + {7'd0,(kernel[1][1] ~^ image[5][4])} + {7'd0,(kernel[1][2] ~^ image[5][5])} + {7'd0,(kernel[1][3] ~^ image[5][6])} + {7'd0,(kernel[1][4] ~^ image[5][7])} + {7'd0,(kernel[2][0] ~^ image[6][3])} + {7'd0,(kernel[2][1] ~^ image[6][4])} + {7'd0,(kernel[2][2] ~^ image[6][5])} + {7'd0,(kernel[2][3] ~^ image[6][6])} + {7'd0,(kernel[2][4] ~^ image[6][7])} + {7'd0,(kernel[3][0] ~^ image[7][3])} + {7'd0,(kernel[3][1] ~^ image[7][4])} + {7'd0,(kernel[3][2] ~^ image[7][5])} + {7'd0,(kernel[3][3] ~^ image[7][6])} + {7'd0,(kernel[3][4] ~^ image[7][7])} + {7'd0,(kernel[4][0] ~^ image[8][3])} + {7'd0,(kernel[4][1] ~^ image[8][4])} + {7'd0,(kernel[4][2] ~^ image[8][5])} + {7'd0,(kernel[4][3] ~^ image[8][6])} + {7'd0,(kernel[4][4] ~^ image[8][7])};
assign out_fmap[4][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][4])} + {7'd0,(kernel[0][1] ~^ image[4][5])} + {7'd0,(kernel[0][2] ~^ image[4][6])} + {7'd0,(kernel[0][3] ~^ image[4][7])} + {7'd0,(kernel[0][4] ~^ image[4][8])} + {7'd0,(kernel[1][0] ~^ image[5][4])} + {7'd0,(kernel[1][1] ~^ image[5][5])} + {7'd0,(kernel[1][2] ~^ image[5][6])} + {7'd0,(kernel[1][3] ~^ image[5][7])} + {7'd0,(kernel[1][4] ~^ image[5][8])} + {7'd0,(kernel[2][0] ~^ image[6][4])} + {7'd0,(kernel[2][1] ~^ image[6][5])} + {7'd0,(kernel[2][2] ~^ image[6][6])} + {7'd0,(kernel[2][3] ~^ image[6][7])} + {7'd0,(kernel[2][4] ~^ image[6][8])} + {7'd0,(kernel[3][0] ~^ image[7][4])} + {7'd0,(kernel[3][1] ~^ image[7][5])} + {7'd0,(kernel[3][2] ~^ image[7][6])} + {7'd0,(kernel[3][3] ~^ image[7][7])} + {7'd0,(kernel[3][4] ~^ image[7][8])} + {7'd0,(kernel[4][0] ~^ image[8][4])} + {7'd0,(kernel[4][1] ~^ image[8][5])} + {7'd0,(kernel[4][2] ~^ image[8][6])} + {7'd0,(kernel[4][3] ~^ image[8][7])} + {7'd0,(kernel[4][4] ~^ image[8][8])};
assign out_fmap[4][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][5])} + {7'd0,(kernel[0][1] ~^ image[4][6])} + {7'd0,(kernel[0][2] ~^ image[4][7])} + {7'd0,(kernel[0][3] ~^ image[4][8])} + {7'd0,(kernel[0][4] ~^ image[4][9])} + {7'd0,(kernel[1][0] ~^ image[5][5])} + {7'd0,(kernel[1][1] ~^ image[5][6])} + {7'd0,(kernel[1][2] ~^ image[5][7])} + {7'd0,(kernel[1][3] ~^ image[5][8])} + {7'd0,(kernel[1][4] ~^ image[5][9])} + {7'd0,(kernel[2][0] ~^ image[6][5])} + {7'd0,(kernel[2][1] ~^ image[6][6])} + {7'd0,(kernel[2][2] ~^ image[6][7])} + {7'd0,(kernel[2][3] ~^ image[6][8])} + {7'd0,(kernel[2][4] ~^ image[6][9])} + {7'd0,(kernel[3][0] ~^ image[7][5])} + {7'd0,(kernel[3][1] ~^ image[7][6])} + {7'd0,(kernel[3][2] ~^ image[7][7])} + {7'd0,(kernel[3][3] ~^ image[7][8])} + {7'd0,(kernel[3][4] ~^ image[7][9])} + {7'd0,(kernel[4][0] ~^ image[8][5])} + {7'd0,(kernel[4][1] ~^ image[8][6])} + {7'd0,(kernel[4][2] ~^ image[8][7])} + {7'd0,(kernel[4][3] ~^ image[8][8])} + {7'd0,(kernel[4][4] ~^ image[8][9])};
assign out_fmap[4][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][6])} + {7'd0,(kernel[0][1] ~^ image[4][7])} + {7'd0,(kernel[0][2] ~^ image[4][8])} + {7'd0,(kernel[0][3] ~^ image[4][9])} + {7'd0,(kernel[0][4] ~^ image[4][10])} + {7'd0,(kernel[1][0] ~^ image[5][6])} + {7'd0,(kernel[1][1] ~^ image[5][7])} + {7'd0,(kernel[1][2] ~^ image[5][8])} + {7'd0,(kernel[1][3] ~^ image[5][9])} + {7'd0,(kernel[1][4] ~^ image[5][10])} + {7'd0,(kernel[2][0] ~^ image[6][6])} + {7'd0,(kernel[2][1] ~^ image[6][7])} + {7'd0,(kernel[2][2] ~^ image[6][8])} + {7'd0,(kernel[2][3] ~^ image[6][9])} + {7'd0,(kernel[2][4] ~^ image[6][10])} + {7'd0,(kernel[3][0] ~^ image[7][6])} + {7'd0,(kernel[3][1] ~^ image[7][7])} + {7'd0,(kernel[3][2] ~^ image[7][8])} + {7'd0,(kernel[3][3] ~^ image[7][9])} + {7'd0,(kernel[3][4] ~^ image[7][10])} + {7'd0,(kernel[4][0] ~^ image[8][6])} + {7'd0,(kernel[4][1] ~^ image[8][7])} + {7'd0,(kernel[4][2] ~^ image[8][8])} + {7'd0,(kernel[4][3] ~^ image[8][9])} + {7'd0,(kernel[4][4] ~^ image[8][10])};
assign out_fmap[4][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][7])} + {7'd0,(kernel[0][1] ~^ image[4][8])} + {7'd0,(kernel[0][2] ~^ image[4][9])} + {7'd0,(kernel[0][3] ~^ image[4][10])} + {7'd0,(kernel[0][4] ~^ image[4][11])} + {7'd0,(kernel[1][0] ~^ image[5][7])} + {7'd0,(kernel[1][1] ~^ image[5][8])} + {7'd0,(kernel[1][2] ~^ image[5][9])} + {7'd0,(kernel[1][3] ~^ image[5][10])} + {7'd0,(kernel[1][4] ~^ image[5][11])} + {7'd0,(kernel[2][0] ~^ image[6][7])} + {7'd0,(kernel[2][1] ~^ image[6][8])} + {7'd0,(kernel[2][2] ~^ image[6][9])} + {7'd0,(kernel[2][3] ~^ image[6][10])} + {7'd0,(kernel[2][4] ~^ image[6][11])} + {7'd0,(kernel[3][0] ~^ image[7][7])} + {7'd0,(kernel[3][1] ~^ image[7][8])} + {7'd0,(kernel[3][2] ~^ image[7][9])} + {7'd0,(kernel[3][3] ~^ image[7][10])} + {7'd0,(kernel[3][4] ~^ image[7][11])} + {7'd0,(kernel[4][0] ~^ image[8][7])} + {7'd0,(kernel[4][1] ~^ image[8][8])} + {7'd0,(kernel[4][2] ~^ image[8][9])} + {7'd0,(kernel[4][3] ~^ image[8][10])} + {7'd0,(kernel[4][4] ~^ image[8][11])};
assign out_fmap[5][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][0])} + {7'd0,(kernel[0][1] ~^ image[5][1])} + {7'd0,(kernel[0][2] ~^ image[5][2])} + {7'd0,(kernel[0][3] ~^ image[5][3])} + {7'd0,(kernel[0][4] ~^ image[5][4])} + {7'd0,(kernel[1][0] ~^ image[6][0])} + {7'd0,(kernel[1][1] ~^ image[6][1])} + {7'd0,(kernel[1][2] ~^ image[6][2])} + {7'd0,(kernel[1][3] ~^ image[6][3])} + {7'd0,(kernel[1][4] ~^ image[6][4])} + {7'd0,(kernel[2][0] ~^ image[7][0])} + {7'd0,(kernel[2][1] ~^ image[7][1])} + {7'd0,(kernel[2][2] ~^ image[7][2])} + {7'd0,(kernel[2][3] ~^ image[7][3])} + {7'd0,(kernel[2][4] ~^ image[7][4])} + {7'd0,(kernel[3][0] ~^ image[8][0])} + {7'd0,(kernel[3][1] ~^ image[8][1])} + {7'd0,(kernel[3][2] ~^ image[8][2])} + {7'd0,(kernel[3][3] ~^ image[8][3])} + {7'd0,(kernel[3][4] ~^ image[8][4])} + {7'd0,(kernel[4][0] ~^ image[9][0])} + {7'd0,(kernel[4][1] ~^ image[9][1])} + {7'd0,(kernel[4][2] ~^ image[9][2])} + {7'd0,(kernel[4][3] ~^ image[9][3])} + {7'd0,(kernel[4][4] ~^ image[9][4])};
assign out_fmap[5][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][1])} + {7'd0,(kernel[0][1] ~^ image[5][2])} + {7'd0,(kernel[0][2] ~^ image[5][3])} + {7'd0,(kernel[0][3] ~^ image[5][4])} + {7'd0,(kernel[0][4] ~^ image[5][5])} + {7'd0,(kernel[1][0] ~^ image[6][1])} + {7'd0,(kernel[1][1] ~^ image[6][2])} + {7'd0,(kernel[1][2] ~^ image[6][3])} + {7'd0,(kernel[1][3] ~^ image[6][4])} + {7'd0,(kernel[1][4] ~^ image[6][5])} + {7'd0,(kernel[2][0] ~^ image[7][1])} + {7'd0,(kernel[2][1] ~^ image[7][2])} + {7'd0,(kernel[2][2] ~^ image[7][3])} + {7'd0,(kernel[2][3] ~^ image[7][4])} + {7'd0,(kernel[2][4] ~^ image[7][5])} + {7'd0,(kernel[3][0] ~^ image[8][1])} + {7'd0,(kernel[3][1] ~^ image[8][2])} + {7'd0,(kernel[3][2] ~^ image[8][3])} + {7'd0,(kernel[3][3] ~^ image[8][4])} + {7'd0,(kernel[3][4] ~^ image[8][5])} + {7'd0,(kernel[4][0] ~^ image[9][1])} + {7'd0,(kernel[4][1] ~^ image[9][2])} + {7'd0,(kernel[4][2] ~^ image[9][3])} + {7'd0,(kernel[4][3] ~^ image[9][4])} + {7'd0,(kernel[4][4] ~^ image[9][5])};
assign out_fmap[5][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][2])} + {7'd0,(kernel[0][1] ~^ image[5][3])} + {7'd0,(kernel[0][2] ~^ image[5][4])} + {7'd0,(kernel[0][3] ~^ image[5][5])} + {7'd0,(kernel[0][4] ~^ image[5][6])} + {7'd0,(kernel[1][0] ~^ image[6][2])} + {7'd0,(kernel[1][1] ~^ image[6][3])} + {7'd0,(kernel[1][2] ~^ image[6][4])} + {7'd0,(kernel[1][3] ~^ image[6][5])} + {7'd0,(kernel[1][4] ~^ image[6][6])} + {7'd0,(kernel[2][0] ~^ image[7][2])} + {7'd0,(kernel[2][1] ~^ image[7][3])} + {7'd0,(kernel[2][2] ~^ image[7][4])} + {7'd0,(kernel[2][3] ~^ image[7][5])} + {7'd0,(kernel[2][4] ~^ image[7][6])} + {7'd0,(kernel[3][0] ~^ image[8][2])} + {7'd0,(kernel[3][1] ~^ image[8][3])} + {7'd0,(kernel[3][2] ~^ image[8][4])} + {7'd0,(kernel[3][3] ~^ image[8][5])} + {7'd0,(kernel[3][4] ~^ image[8][6])} + {7'd0,(kernel[4][0] ~^ image[9][2])} + {7'd0,(kernel[4][1] ~^ image[9][3])} + {7'd0,(kernel[4][2] ~^ image[9][4])} + {7'd0,(kernel[4][3] ~^ image[9][5])} + {7'd0,(kernel[4][4] ~^ image[9][6])};
assign out_fmap[5][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][3])} + {7'd0,(kernel[0][1] ~^ image[5][4])} + {7'd0,(kernel[0][2] ~^ image[5][5])} + {7'd0,(kernel[0][3] ~^ image[5][6])} + {7'd0,(kernel[0][4] ~^ image[5][7])} + {7'd0,(kernel[1][0] ~^ image[6][3])} + {7'd0,(kernel[1][1] ~^ image[6][4])} + {7'd0,(kernel[1][2] ~^ image[6][5])} + {7'd0,(kernel[1][3] ~^ image[6][6])} + {7'd0,(kernel[1][4] ~^ image[6][7])} + {7'd0,(kernel[2][0] ~^ image[7][3])} + {7'd0,(kernel[2][1] ~^ image[7][4])} + {7'd0,(kernel[2][2] ~^ image[7][5])} + {7'd0,(kernel[2][3] ~^ image[7][6])} + {7'd0,(kernel[2][4] ~^ image[7][7])} + {7'd0,(kernel[3][0] ~^ image[8][3])} + {7'd0,(kernel[3][1] ~^ image[8][4])} + {7'd0,(kernel[3][2] ~^ image[8][5])} + {7'd0,(kernel[3][3] ~^ image[8][6])} + {7'd0,(kernel[3][4] ~^ image[8][7])} + {7'd0,(kernel[4][0] ~^ image[9][3])} + {7'd0,(kernel[4][1] ~^ image[9][4])} + {7'd0,(kernel[4][2] ~^ image[9][5])} + {7'd0,(kernel[4][3] ~^ image[9][6])} + {7'd0,(kernel[4][4] ~^ image[9][7])};
assign out_fmap[5][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][4])} + {7'd0,(kernel[0][1] ~^ image[5][5])} + {7'd0,(kernel[0][2] ~^ image[5][6])} + {7'd0,(kernel[0][3] ~^ image[5][7])} + {7'd0,(kernel[0][4] ~^ image[5][8])} + {7'd0,(kernel[1][0] ~^ image[6][4])} + {7'd0,(kernel[1][1] ~^ image[6][5])} + {7'd0,(kernel[1][2] ~^ image[6][6])} + {7'd0,(kernel[1][3] ~^ image[6][7])} + {7'd0,(kernel[1][4] ~^ image[6][8])} + {7'd0,(kernel[2][0] ~^ image[7][4])} + {7'd0,(kernel[2][1] ~^ image[7][5])} + {7'd0,(kernel[2][2] ~^ image[7][6])} + {7'd0,(kernel[2][3] ~^ image[7][7])} + {7'd0,(kernel[2][4] ~^ image[7][8])} + {7'd0,(kernel[3][0] ~^ image[8][4])} + {7'd0,(kernel[3][1] ~^ image[8][5])} + {7'd0,(kernel[3][2] ~^ image[8][6])} + {7'd0,(kernel[3][3] ~^ image[8][7])} + {7'd0,(kernel[3][4] ~^ image[8][8])} + {7'd0,(kernel[4][0] ~^ image[9][4])} + {7'd0,(kernel[4][1] ~^ image[9][5])} + {7'd0,(kernel[4][2] ~^ image[9][6])} + {7'd0,(kernel[4][3] ~^ image[9][7])} + {7'd0,(kernel[4][4] ~^ image[9][8])};
assign out_fmap[5][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][5])} + {7'd0,(kernel[0][1] ~^ image[5][6])} + {7'd0,(kernel[0][2] ~^ image[5][7])} + {7'd0,(kernel[0][3] ~^ image[5][8])} + {7'd0,(kernel[0][4] ~^ image[5][9])} + {7'd0,(kernel[1][0] ~^ image[6][5])} + {7'd0,(kernel[1][1] ~^ image[6][6])} + {7'd0,(kernel[1][2] ~^ image[6][7])} + {7'd0,(kernel[1][3] ~^ image[6][8])} + {7'd0,(kernel[1][4] ~^ image[6][9])} + {7'd0,(kernel[2][0] ~^ image[7][5])} + {7'd0,(kernel[2][1] ~^ image[7][6])} + {7'd0,(kernel[2][2] ~^ image[7][7])} + {7'd0,(kernel[2][3] ~^ image[7][8])} + {7'd0,(kernel[2][4] ~^ image[7][9])} + {7'd0,(kernel[3][0] ~^ image[8][5])} + {7'd0,(kernel[3][1] ~^ image[8][6])} + {7'd0,(kernel[3][2] ~^ image[8][7])} + {7'd0,(kernel[3][3] ~^ image[8][8])} + {7'd0,(kernel[3][4] ~^ image[8][9])} + {7'd0,(kernel[4][0] ~^ image[9][5])} + {7'd0,(kernel[4][1] ~^ image[9][6])} + {7'd0,(kernel[4][2] ~^ image[9][7])} + {7'd0,(kernel[4][3] ~^ image[9][8])} + {7'd0,(kernel[4][4] ~^ image[9][9])};
assign out_fmap[5][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][6])} + {7'd0,(kernel[0][1] ~^ image[5][7])} + {7'd0,(kernel[0][2] ~^ image[5][8])} + {7'd0,(kernel[0][3] ~^ image[5][9])} + {7'd0,(kernel[0][4] ~^ image[5][10])} + {7'd0,(kernel[1][0] ~^ image[6][6])} + {7'd0,(kernel[1][1] ~^ image[6][7])} + {7'd0,(kernel[1][2] ~^ image[6][8])} + {7'd0,(kernel[1][3] ~^ image[6][9])} + {7'd0,(kernel[1][4] ~^ image[6][10])} + {7'd0,(kernel[2][0] ~^ image[7][6])} + {7'd0,(kernel[2][1] ~^ image[7][7])} + {7'd0,(kernel[2][2] ~^ image[7][8])} + {7'd0,(kernel[2][3] ~^ image[7][9])} + {7'd0,(kernel[2][4] ~^ image[7][10])} + {7'd0,(kernel[3][0] ~^ image[8][6])} + {7'd0,(kernel[3][1] ~^ image[8][7])} + {7'd0,(kernel[3][2] ~^ image[8][8])} + {7'd0,(kernel[3][3] ~^ image[8][9])} + {7'd0,(kernel[3][4] ~^ image[8][10])} + {7'd0,(kernel[4][0] ~^ image[9][6])} + {7'd0,(kernel[4][1] ~^ image[9][7])} + {7'd0,(kernel[4][2] ~^ image[9][8])} + {7'd0,(kernel[4][3] ~^ image[9][9])} + {7'd0,(kernel[4][4] ~^ image[9][10])};
assign out_fmap[5][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][7])} + {7'd0,(kernel[0][1] ~^ image[5][8])} + {7'd0,(kernel[0][2] ~^ image[5][9])} + {7'd0,(kernel[0][3] ~^ image[5][10])} + {7'd0,(kernel[0][4] ~^ image[5][11])} + {7'd0,(kernel[1][0] ~^ image[6][7])} + {7'd0,(kernel[1][1] ~^ image[6][8])} + {7'd0,(kernel[1][2] ~^ image[6][9])} + {7'd0,(kernel[1][3] ~^ image[6][10])} + {7'd0,(kernel[1][4] ~^ image[6][11])} + {7'd0,(kernel[2][0] ~^ image[7][7])} + {7'd0,(kernel[2][1] ~^ image[7][8])} + {7'd0,(kernel[2][2] ~^ image[7][9])} + {7'd0,(kernel[2][3] ~^ image[7][10])} + {7'd0,(kernel[2][4] ~^ image[7][11])} + {7'd0,(kernel[3][0] ~^ image[8][7])} + {7'd0,(kernel[3][1] ~^ image[8][8])} + {7'd0,(kernel[3][2] ~^ image[8][9])} + {7'd0,(kernel[3][3] ~^ image[8][10])} + {7'd0,(kernel[3][4] ~^ image[8][11])} + {7'd0,(kernel[4][0] ~^ image[9][7])} + {7'd0,(kernel[4][1] ~^ image[9][8])} + {7'd0,(kernel[4][2] ~^ image[9][9])} + {7'd0,(kernel[4][3] ~^ image[9][10])} + {7'd0,(kernel[4][4] ~^ image[9][11])};
assign out_fmap[6][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][0])} + {7'd0,(kernel[0][1] ~^ image[6][1])} + {7'd0,(kernel[0][2] ~^ image[6][2])} + {7'd0,(kernel[0][3] ~^ image[6][3])} + {7'd0,(kernel[0][4] ~^ image[6][4])} + {7'd0,(kernel[1][0] ~^ image[7][0])} + {7'd0,(kernel[1][1] ~^ image[7][1])} + {7'd0,(kernel[1][2] ~^ image[7][2])} + {7'd0,(kernel[1][3] ~^ image[7][3])} + {7'd0,(kernel[1][4] ~^ image[7][4])} + {7'd0,(kernel[2][0] ~^ image[8][0])} + {7'd0,(kernel[2][1] ~^ image[8][1])} + {7'd0,(kernel[2][2] ~^ image[8][2])} + {7'd0,(kernel[2][3] ~^ image[8][3])} + {7'd0,(kernel[2][4] ~^ image[8][4])} + {7'd0,(kernel[3][0] ~^ image[9][0])} + {7'd0,(kernel[3][1] ~^ image[9][1])} + {7'd0,(kernel[3][2] ~^ image[9][2])} + {7'd0,(kernel[3][3] ~^ image[9][3])} + {7'd0,(kernel[3][4] ~^ image[9][4])} + {7'd0,(kernel[4][0] ~^ image[10][0])} + {7'd0,(kernel[4][1] ~^ image[10][1])} + {7'd0,(kernel[4][2] ~^ image[10][2])} + {7'd0,(kernel[4][3] ~^ image[10][3])} + {7'd0,(kernel[4][4] ~^ image[10][4])};
assign out_fmap[6][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][1])} + {7'd0,(kernel[0][1] ~^ image[6][2])} + {7'd0,(kernel[0][2] ~^ image[6][3])} + {7'd0,(kernel[0][3] ~^ image[6][4])} + {7'd0,(kernel[0][4] ~^ image[6][5])} + {7'd0,(kernel[1][0] ~^ image[7][1])} + {7'd0,(kernel[1][1] ~^ image[7][2])} + {7'd0,(kernel[1][2] ~^ image[7][3])} + {7'd0,(kernel[1][3] ~^ image[7][4])} + {7'd0,(kernel[1][4] ~^ image[7][5])} + {7'd0,(kernel[2][0] ~^ image[8][1])} + {7'd0,(kernel[2][1] ~^ image[8][2])} + {7'd0,(kernel[2][2] ~^ image[8][3])} + {7'd0,(kernel[2][3] ~^ image[8][4])} + {7'd0,(kernel[2][4] ~^ image[8][5])} + {7'd0,(kernel[3][0] ~^ image[9][1])} + {7'd0,(kernel[3][1] ~^ image[9][2])} + {7'd0,(kernel[3][2] ~^ image[9][3])} + {7'd0,(kernel[3][3] ~^ image[9][4])} + {7'd0,(kernel[3][4] ~^ image[9][5])} + {7'd0,(kernel[4][0] ~^ image[10][1])} + {7'd0,(kernel[4][1] ~^ image[10][2])} + {7'd0,(kernel[4][2] ~^ image[10][3])} + {7'd0,(kernel[4][3] ~^ image[10][4])} + {7'd0,(kernel[4][4] ~^ image[10][5])};
assign out_fmap[6][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][2])} + {7'd0,(kernel[0][1] ~^ image[6][3])} + {7'd0,(kernel[0][2] ~^ image[6][4])} + {7'd0,(kernel[0][3] ~^ image[6][5])} + {7'd0,(kernel[0][4] ~^ image[6][6])} + {7'd0,(kernel[1][0] ~^ image[7][2])} + {7'd0,(kernel[1][1] ~^ image[7][3])} + {7'd0,(kernel[1][2] ~^ image[7][4])} + {7'd0,(kernel[1][3] ~^ image[7][5])} + {7'd0,(kernel[1][4] ~^ image[7][6])} + {7'd0,(kernel[2][0] ~^ image[8][2])} + {7'd0,(kernel[2][1] ~^ image[8][3])} + {7'd0,(kernel[2][2] ~^ image[8][4])} + {7'd0,(kernel[2][3] ~^ image[8][5])} + {7'd0,(kernel[2][4] ~^ image[8][6])} + {7'd0,(kernel[3][0] ~^ image[9][2])} + {7'd0,(kernel[3][1] ~^ image[9][3])} + {7'd0,(kernel[3][2] ~^ image[9][4])} + {7'd0,(kernel[3][3] ~^ image[9][5])} + {7'd0,(kernel[3][4] ~^ image[9][6])} + {7'd0,(kernel[4][0] ~^ image[10][2])} + {7'd0,(kernel[4][1] ~^ image[10][3])} + {7'd0,(kernel[4][2] ~^ image[10][4])} + {7'd0,(kernel[4][3] ~^ image[10][5])} + {7'd0,(kernel[4][4] ~^ image[10][6])};
assign out_fmap[6][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][3])} + {7'd0,(kernel[0][1] ~^ image[6][4])} + {7'd0,(kernel[0][2] ~^ image[6][5])} + {7'd0,(kernel[0][3] ~^ image[6][6])} + {7'd0,(kernel[0][4] ~^ image[6][7])} + {7'd0,(kernel[1][0] ~^ image[7][3])} + {7'd0,(kernel[1][1] ~^ image[7][4])} + {7'd0,(kernel[1][2] ~^ image[7][5])} + {7'd0,(kernel[1][3] ~^ image[7][6])} + {7'd0,(kernel[1][4] ~^ image[7][7])} + {7'd0,(kernel[2][0] ~^ image[8][3])} + {7'd0,(kernel[2][1] ~^ image[8][4])} + {7'd0,(kernel[2][2] ~^ image[8][5])} + {7'd0,(kernel[2][3] ~^ image[8][6])} + {7'd0,(kernel[2][4] ~^ image[8][7])} + {7'd0,(kernel[3][0] ~^ image[9][3])} + {7'd0,(kernel[3][1] ~^ image[9][4])} + {7'd0,(kernel[3][2] ~^ image[9][5])} + {7'd0,(kernel[3][3] ~^ image[9][6])} + {7'd0,(kernel[3][4] ~^ image[9][7])} + {7'd0,(kernel[4][0] ~^ image[10][3])} + {7'd0,(kernel[4][1] ~^ image[10][4])} + {7'd0,(kernel[4][2] ~^ image[10][5])} + {7'd0,(kernel[4][3] ~^ image[10][6])} + {7'd0,(kernel[4][4] ~^ image[10][7])};
assign out_fmap[6][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][4])} + {7'd0,(kernel[0][1] ~^ image[6][5])} + {7'd0,(kernel[0][2] ~^ image[6][6])} + {7'd0,(kernel[0][3] ~^ image[6][7])} + {7'd0,(kernel[0][4] ~^ image[6][8])} + {7'd0,(kernel[1][0] ~^ image[7][4])} + {7'd0,(kernel[1][1] ~^ image[7][5])} + {7'd0,(kernel[1][2] ~^ image[7][6])} + {7'd0,(kernel[1][3] ~^ image[7][7])} + {7'd0,(kernel[1][4] ~^ image[7][8])} + {7'd0,(kernel[2][0] ~^ image[8][4])} + {7'd0,(kernel[2][1] ~^ image[8][5])} + {7'd0,(kernel[2][2] ~^ image[8][6])} + {7'd0,(kernel[2][3] ~^ image[8][7])} + {7'd0,(kernel[2][4] ~^ image[8][8])} + {7'd0,(kernel[3][0] ~^ image[9][4])} + {7'd0,(kernel[3][1] ~^ image[9][5])} + {7'd0,(kernel[3][2] ~^ image[9][6])} + {7'd0,(kernel[3][3] ~^ image[9][7])} + {7'd0,(kernel[3][4] ~^ image[9][8])} + {7'd0,(kernel[4][0] ~^ image[10][4])} + {7'd0,(kernel[4][1] ~^ image[10][5])} + {7'd0,(kernel[4][2] ~^ image[10][6])} + {7'd0,(kernel[4][3] ~^ image[10][7])} + {7'd0,(kernel[4][4] ~^ image[10][8])};
assign out_fmap[6][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][5])} + {7'd0,(kernel[0][1] ~^ image[6][6])} + {7'd0,(kernel[0][2] ~^ image[6][7])} + {7'd0,(kernel[0][3] ~^ image[6][8])} + {7'd0,(kernel[0][4] ~^ image[6][9])} + {7'd0,(kernel[1][0] ~^ image[7][5])} + {7'd0,(kernel[1][1] ~^ image[7][6])} + {7'd0,(kernel[1][2] ~^ image[7][7])} + {7'd0,(kernel[1][3] ~^ image[7][8])} + {7'd0,(kernel[1][4] ~^ image[7][9])} + {7'd0,(kernel[2][0] ~^ image[8][5])} + {7'd0,(kernel[2][1] ~^ image[8][6])} + {7'd0,(kernel[2][2] ~^ image[8][7])} + {7'd0,(kernel[2][3] ~^ image[8][8])} + {7'd0,(kernel[2][4] ~^ image[8][9])} + {7'd0,(kernel[3][0] ~^ image[9][5])} + {7'd0,(kernel[3][1] ~^ image[9][6])} + {7'd0,(kernel[3][2] ~^ image[9][7])} + {7'd0,(kernel[3][3] ~^ image[9][8])} + {7'd0,(kernel[3][4] ~^ image[9][9])} + {7'd0,(kernel[4][0] ~^ image[10][5])} + {7'd0,(kernel[4][1] ~^ image[10][6])} + {7'd0,(kernel[4][2] ~^ image[10][7])} + {7'd0,(kernel[4][3] ~^ image[10][8])} + {7'd0,(kernel[4][4] ~^ image[10][9])};
assign out_fmap[6][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][6])} + {7'd0,(kernel[0][1] ~^ image[6][7])} + {7'd0,(kernel[0][2] ~^ image[6][8])} + {7'd0,(kernel[0][3] ~^ image[6][9])} + {7'd0,(kernel[0][4] ~^ image[6][10])} + {7'd0,(kernel[1][0] ~^ image[7][6])} + {7'd0,(kernel[1][1] ~^ image[7][7])} + {7'd0,(kernel[1][2] ~^ image[7][8])} + {7'd0,(kernel[1][3] ~^ image[7][9])} + {7'd0,(kernel[1][4] ~^ image[7][10])} + {7'd0,(kernel[2][0] ~^ image[8][6])} + {7'd0,(kernel[2][1] ~^ image[8][7])} + {7'd0,(kernel[2][2] ~^ image[8][8])} + {7'd0,(kernel[2][3] ~^ image[8][9])} + {7'd0,(kernel[2][4] ~^ image[8][10])} + {7'd0,(kernel[3][0] ~^ image[9][6])} + {7'd0,(kernel[3][1] ~^ image[9][7])} + {7'd0,(kernel[3][2] ~^ image[9][8])} + {7'd0,(kernel[3][3] ~^ image[9][9])} + {7'd0,(kernel[3][4] ~^ image[9][10])} + {7'd0,(kernel[4][0] ~^ image[10][6])} + {7'd0,(kernel[4][1] ~^ image[10][7])} + {7'd0,(kernel[4][2] ~^ image[10][8])} + {7'd0,(kernel[4][3] ~^ image[10][9])} + {7'd0,(kernel[4][4] ~^ image[10][10])};
assign out_fmap[6][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][7])} + {7'd0,(kernel[0][1] ~^ image[6][8])} + {7'd0,(kernel[0][2] ~^ image[6][9])} + {7'd0,(kernel[0][3] ~^ image[6][10])} + {7'd0,(kernel[0][4] ~^ image[6][11])} + {7'd0,(kernel[1][0] ~^ image[7][7])} + {7'd0,(kernel[1][1] ~^ image[7][8])} + {7'd0,(kernel[1][2] ~^ image[7][9])} + {7'd0,(kernel[1][3] ~^ image[7][10])} + {7'd0,(kernel[1][4] ~^ image[7][11])} + {7'd0,(kernel[2][0] ~^ image[8][7])} + {7'd0,(kernel[2][1] ~^ image[8][8])} + {7'd0,(kernel[2][2] ~^ image[8][9])} + {7'd0,(kernel[2][3] ~^ image[8][10])} + {7'd0,(kernel[2][4] ~^ image[8][11])} + {7'd0,(kernel[3][0] ~^ image[9][7])} + {7'd0,(kernel[3][1] ~^ image[9][8])} + {7'd0,(kernel[3][2] ~^ image[9][9])} + {7'd0,(kernel[3][3] ~^ image[9][10])} + {7'd0,(kernel[3][4] ~^ image[9][11])} + {7'd0,(kernel[4][0] ~^ image[10][7])} + {7'd0,(kernel[4][1] ~^ image[10][8])} + {7'd0,(kernel[4][2] ~^ image[10][9])} + {7'd0,(kernel[4][3] ~^ image[10][10])} + {7'd0,(kernel[4][4] ~^ image[10][11])};
assign out_fmap[7][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][0])} + {7'd0,(kernel[0][1] ~^ image[7][1])} + {7'd0,(kernel[0][2] ~^ image[7][2])} + {7'd0,(kernel[0][3] ~^ image[7][3])} + {7'd0,(kernel[0][4] ~^ image[7][4])} + {7'd0,(kernel[1][0] ~^ image[8][0])} + {7'd0,(kernel[1][1] ~^ image[8][1])} + {7'd0,(kernel[1][2] ~^ image[8][2])} + {7'd0,(kernel[1][3] ~^ image[8][3])} + {7'd0,(kernel[1][4] ~^ image[8][4])} + {7'd0,(kernel[2][0] ~^ image[9][0])} + {7'd0,(kernel[2][1] ~^ image[9][1])} + {7'd0,(kernel[2][2] ~^ image[9][2])} + {7'd0,(kernel[2][3] ~^ image[9][3])} + {7'd0,(kernel[2][4] ~^ image[9][4])} + {7'd0,(kernel[3][0] ~^ image[10][0])} + {7'd0,(kernel[3][1] ~^ image[10][1])} + {7'd0,(kernel[3][2] ~^ image[10][2])} + {7'd0,(kernel[3][3] ~^ image[10][3])} + {7'd0,(kernel[3][4] ~^ image[10][4])} + {7'd0,(kernel[4][0] ~^ image[11][0])} + {7'd0,(kernel[4][1] ~^ image[11][1])} + {7'd0,(kernel[4][2] ~^ image[11][2])} + {7'd0,(kernel[4][3] ~^ image[11][3])} + {7'd0,(kernel[4][4] ~^ image[11][4])};
assign out_fmap[7][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][1])} + {7'd0,(kernel[0][1] ~^ image[7][2])} + {7'd0,(kernel[0][2] ~^ image[7][3])} + {7'd0,(kernel[0][3] ~^ image[7][4])} + {7'd0,(kernel[0][4] ~^ image[7][5])} + {7'd0,(kernel[1][0] ~^ image[8][1])} + {7'd0,(kernel[1][1] ~^ image[8][2])} + {7'd0,(kernel[1][2] ~^ image[8][3])} + {7'd0,(kernel[1][3] ~^ image[8][4])} + {7'd0,(kernel[1][4] ~^ image[8][5])} + {7'd0,(kernel[2][0] ~^ image[9][1])} + {7'd0,(kernel[2][1] ~^ image[9][2])} + {7'd0,(kernel[2][2] ~^ image[9][3])} + {7'd0,(kernel[2][3] ~^ image[9][4])} + {7'd0,(kernel[2][4] ~^ image[9][5])} + {7'd0,(kernel[3][0] ~^ image[10][1])} + {7'd0,(kernel[3][1] ~^ image[10][2])} + {7'd0,(kernel[3][2] ~^ image[10][3])} + {7'd0,(kernel[3][3] ~^ image[10][4])} + {7'd0,(kernel[3][4] ~^ image[10][5])} + {7'd0,(kernel[4][0] ~^ image[11][1])} + {7'd0,(kernel[4][1] ~^ image[11][2])} + {7'd0,(kernel[4][2] ~^ image[11][3])} + {7'd0,(kernel[4][3] ~^ image[11][4])} + {7'd0,(kernel[4][4] ~^ image[11][5])};
assign out_fmap[7][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][2])} + {7'd0,(kernel[0][1] ~^ image[7][3])} + {7'd0,(kernel[0][2] ~^ image[7][4])} + {7'd0,(kernel[0][3] ~^ image[7][5])} + {7'd0,(kernel[0][4] ~^ image[7][6])} + {7'd0,(kernel[1][0] ~^ image[8][2])} + {7'd0,(kernel[1][1] ~^ image[8][3])} + {7'd0,(kernel[1][2] ~^ image[8][4])} + {7'd0,(kernel[1][3] ~^ image[8][5])} + {7'd0,(kernel[1][4] ~^ image[8][6])} + {7'd0,(kernel[2][0] ~^ image[9][2])} + {7'd0,(kernel[2][1] ~^ image[9][3])} + {7'd0,(kernel[2][2] ~^ image[9][4])} + {7'd0,(kernel[2][3] ~^ image[9][5])} + {7'd0,(kernel[2][4] ~^ image[9][6])} + {7'd0,(kernel[3][0] ~^ image[10][2])} + {7'd0,(kernel[3][1] ~^ image[10][3])} + {7'd0,(kernel[3][2] ~^ image[10][4])} + {7'd0,(kernel[3][3] ~^ image[10][5])} + {7'd0,(kernel[3][4] ~^ image[10][6])} + {7'd0,(kernel[4][0] ~^ image[11][2])} + {7'd0,(kernel[4][1] ~^ image[11][3])} + {7'd0,(kernel[4][2] ~^ image[11][4])} + {7'd0,(kernel[4][3] ~^ image[11][5])} + {7'd0,(kernel[4][4] ~^ image[11][6])};
assign out_fmap[7][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][3])} + {7'd0,(kernel[0][1] ~^ image[7][4])} + {7'd0,(kernel[0][2] ~^ image[7][5])} + {7'd0,(kernel[0][3] ~^ image[7][6])} + {7'd0,(kernel[0][4] ~^ image[7][7])} + {7'd0,(kernel[1][0] ~^ image[8][3])} + {7'd0,(kernel[1][1] ~^ image[8][4])} + {7'd0,(kernel[1][2] ~^ image[8][5])} + {7'd0,(kernel[1][3] ~^ image[8][6])} + {7'd0,(kernel[1][4] ~^ image[8][7])} + {7'd0,(kernel[2][0] ~^ image[9][3])} + {7'd0,(kernel[2][1] ~^ image[9][4])} + {7'd0,(kernel[2][2] ~^ image[9][5])} + {7'd0,(kernel[2][3] ~^ image[9][6])} + {7'd0,(kernel[2][4] ~^ image[9][7])} + {7'd0,(kernel[3][0] ~^ image[10][3])} + {7'd0,(kernel[3][1] ~^ image[10][4])} + {7'd0,(kernel[3][2] ~^ image[10][5])} + {7'd0,(kernel[3][3] ~^ image[10][6])} + {7'd0,(kernel[3][4] ~^ image[10][7])} + {7'd0,(kernel[4][0] ~^ image[11][3])} + {7'd0,(kernel[4][1] ~^ image[11][4])} + {7'd0,(kernel[4][2] ~^ image[11][5])} + {7'd0,(kernel[4][3] ~^ image[11][6])} + {7'd0,(kernel[4][4] ~^ image[11][7])};
assign out_fmap[7][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][4])} + {7'd0,(kernel[0][1] ~^ image[7][5])} + {7'd0,(kernel[0][2] ~^ image[7][6])} + {7'd0,(kernel[0][3] ~^ image[7][7])} + {7'd0,(kernel[0][4] ~^ image[7][8])} + {7'd0,(kernel[1][0] ~^ image[8][4])} + {7'd0,(kernel[1][1] ~^ image[8][5])} + {7'd0,(kernel[1][2] ~^ image[8][6])} + {7'd0,(kernel[1][3] ~^ image[8][7])} + {7'd0,(kernel[1][4] ~^ image[8][8])} + {7'd0,(kernel[2][0] ~^ image[9][4])} + {7'd0,(kernel[2][1] ~^ image[9][5])} + {7'd0,(kernel[2][2] ~^ image[9][6])} + {7'd0,(kernel[2][3] ~^ image[9][7])} + {7'd0,(kernel[2][4] ~^ image[9][8])} + {7'd0,(kernel[3][0] ~^ image[10][4])} + {7'd0,(kernel[3][1] ~^ image[10][5])} + {7'd0,(kernel[3][2] ~^ image[10][6])} + {7'd0,(kernel[3][3] ~^ image[10][7])} + {7'd0,(kernel[3][4] ~^ image[10][8])} + {7'd0,(kernel[4][0] ~^ image[11][4])} + {7'd0,(kernel[4][1] ~^ image[11][5])} + {7'd0,(kernel[4][2] ~^ image[11][6])} + {7'd0,(kernel[4][3] ~^ image[11][7])} + {7'd0,(kernel[4][4] ~^ image[11][8])};
assign out_fmap[7][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][5])} + {7'd0,(kernel[0][1] ~^ image[7][6])} + {7'd0,(kernel[0][2] ~^ image[7][7])} + {7'd0,(kernel[0][3] ~^ image[7][8])} + {7'd0,(kernel[0][4] ~^ image[7][9])} + {7'd0,(kernel[1][0] ~^ image[8][5])} + {7'd0,(kernel[1][1] ~^ image[8][6])} + {7'd0,(kernel[1][2] ~^ image[8][7])} + {7'd0,(kernel[1][3] ~^ image[8][8])} + {7'd0,(kernel[1][4] ~^ image[8][9])} + {7'd0,(kernel[2][0] ~^ image[9][5])} + {7'd0,(kernel[2][1] ~^ image[9][6])} + {7'd0,(kernel[2][2] ~^ image[9][7])} + {7'd0,(kernel[2][3] ~^ image[9][8])} + {7'd0,(kernel[2][4] ~^ image[9][9])} + {7'd0,(kernel[3][0] ~^ image[10][5])} + {7'd0,(kernel[3][1] ~^ image[10][6])} + {7'd0,(kernel[3][2] ~^ image[10][7])} + {7'd0,(kernel[3][3] ~^ image[10][8])} + {7'd0,(kernel[3][4] ~^ image[10][9])} + {7'd0,(kernel[4][0] ~^ image[11][5])} + {7'd0,(kernel[4][1] ~^ image[11][6])} + {7'd0,(kernel[4][2] ~^ image[11][7])} + {7'd0,(kernel[4][3] ~^ image[11][8])} + {7'd0,(kernel[4][4] ~^ image[11][9])};
assign out_fmap[7][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][6])} + {7'd0,(kernel[0][1] ~^ image[7][7])} + {7'd0,(kernel[0][2] ~^ image[7][8])} + {7'd0,(kernel[0][3] ~^ image[7][9])} + {7'd0,(kernel[0][4] ~^ image[7][10])} + {7'd0,(kernel[1][0] ~^ image[8][6])} + {7'd0,(kernel[1][1] ~^ image[8][7])} + {7'd0,(kernel[1][2] ~^ image[8][8])} + {7'd0,(kernel[1][3] ~^ image[8][9])} + {7'd0,(kernel[1][4] ~^ image[8][10])} + {7'd0,(kernel[2][0] ~^ image[9][6])} + {7'd0,(kernel[2][1] ~^ image[9][7])} + {7'd0,(kernel[2][2] ~^ image[9][8])} + {7'd0,(kernel[2][3] ~^ image[9][9])} + {7'd0,(kernel[2][4] ~^ image[9][10])} + {7'd0,(kernel[3][0] ~^ image[10][6])} + {7'd0,(kernel[3][1] ~^ image[10][7])} + {7'd0,(kernel[3][2] ~^ image[10][8])} + {7'd0,(kernel[3][3] ~^ image[10][9])} + {7'd0,(kernel[3][4] ~^ image[10][10])} + {7'd0,(kernel[4][0] ~^ image[11][6])} + {7'd0,(kernel[4][1] ~^ image[11][7])} + {7'd0,(kernel[4][2] ~^ image[11][8])} + {7'd0,(kernel[4][3] ~^ image[11][9])} + {7'd0,(kernel[4][4] ~^ image[11][10])};
assign out_fmap[7][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][7])} + {7'd0,(kernel[0][1] ~^ image[7][8])} + {7'd0,(kernel[0][2] ~^ image[7][9])} + {7'd0,(kernel[0][3] ~^ image[7][10])} + {7'd0,(kernel[0][4] ~^ image[7][11])} + {7'd0,(kernel[1][0] ~^ image[8][7])} + {7'd0,(kernel[1][1] ~^ image[8][8])} + {7'd0,(kernel[1][2] ~^ image[8][9])} + {7'd0,(kernel[1][3] ~^ image[8][10])} + {7'd0,(kernel[1][4] ~^ image[8][11])} + {7'd0,(kernel[2][0] ~^ image[9][7])} + {7'd0,(kernel[2][1] ~^ image[9][8])} + {7'd0,(kernel[2][2] ~^ image[9][9])} + {7'd0,(kernel[2][3] ~^ image[9][10])} + {7'd0,(kernel[2][4] ~^ image[9][11])} + {7'd0,(kernel[3][0] ~^ image[10][7])} + {7'd0,(kernel[3][1] ~^ image[10][8])} + {7'd0,(kernel[3][2] ~^ image[10][9])} + {7'd0,(kernel[3][3] ~^ image[10][10])} + {7'd0,(kernel[3][4] ~^ image[10][11])} + {7'd0,(kernel[4][0] ~^ image[11][7])} + {7'd0,(kernel[4][1] ~^ image[11][8])} + {7'd0,(kernel[4][2] ~^ image[11][9])} + {7'd0,(kernel[4][3] ~^ image[11][10])} + {7'd0,(kernel[4][4] ~^ image[11][11])};

endmodule