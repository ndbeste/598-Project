module convchan2
    #( parameter bW = 8 )
    ( 
    input  logic          image     [0:11][0:11],
    input  logic          kernel    [0:4] [0:4],
    output logic [bW-1:0] out_fmap  [0:7][0:7]
    );

assign out_fmap[0][0] = kernel[0][0] ~^ image[0][0] + kernel[0][1] ~^ image[0][1] + kernel[0][2] ~^ image[0][2] + kernel[0][3] ~^ image[0][3] + kernel[0][4] ~^ image[0][4] + kernel[1][0] ~^ image[1][0] + kernel[1][1] ~^ image[1][1] + kernel[1][2] ~^ image[1][2] + kernel[1][3] ~^ image[1][3] + kernel[1][4] ~^ image[1][4] + kernel[2][0] ~^ image[2][0] + kernel[2][1] ~^ image[2][1] + kernel[2][2] ~^ image[2][2] + kernel[2][3] ~^ image[2][3] + kernel[2][4] ~^ image[2][4] + kernel[3][0] ~^ image[3][0] + kernel[3][1] ~^ image[3][1] + kernel[3][2] ~^ image[3][2] + kernel[3][3] ~^ image[3][3] + kernel[3][4] ~^ image[3][4] + kernel[4][0] ~^ image[4][0] + kernel[4][1] ~^ image[4][1] + kernel[4][2] ~^ image[4][2] + kernel[4][3] ~^ image[4][3] + kernel[4][4] ~^ image[4][4];
assign out_fmap[0][1] = kernel[0][0] ~^ image[0][1] + kernel[0][1] ~^ image[0][2] + kernel[0][2] ~^ image[0][3] + kernel[0][3] ~^ image[0][4] + kernel[0][4] ~^ image[0][5] + kernel[1][0] ~^ image[1][1] + kernel[1][1] ~^ image[1][2] + kernel[1][2] ~^ image[1][3] + kernel[1][3] ~^ image[1][4] + kernel[1][4] ~^ image[1][5] + kernel[2][0] ~^ image[2][1] + kernel[2][1] ~^ image[2][2] + kernel[2][2] ~^ image[2][3] + kernel[2][3] ~^ image[2][4] + kernel[2][4] ~^ image[2][5] + kernel[3][0] ~^ image[3][1] + kernel[3][1] ~^ image[3][2] + kernel[3][2] ~^ image[3][3] + kernel[3][3] ~^ image[3][4] + kernel[3][4] ~^ image[3][5] + kernel[4][0] ~^ image[4][1] + kernel[4][1] ~^ image[4][2] + kernel[4][2] ~^ image[4][3] + kernel[4][3] ~^ image[4][4] + kernel[4][4] ~^ image[4][5];
assign out_fmap[0][2] = kernel[0][0] ~^ image[0][2] + kernel[0][1] ~^ image[0][3] + kernel[0][2] ~^ image[0][4] + kernel[0][3] ~^ image[0][5] + kernel[0][4] ~^ image[0][6] + kernel[1][0] ~^ image[1][2] + kernel[1][1] ~^ image[1][3] + kernel[1][2] ~^ image[1][4] + kernel[1][3] ~^ image[1][5] + kernel[1][4] ~^ image[1][6] + kernel[2][0] ~^ image[2][2] + kernel[2][1] ~^ image[2][3] + kernel[2][2] ~^ image[2][4] + kernel[2][3] ~^ image[2][5] + kernel[2][4] ~^ image[2][6] + kernel[3][0] ~^ image[3][2] + kernel[3][1] ~^ image[3][3] + kernel[3][2] ~^ image[3][4] + kernel[3][3] ~^ image[3][5] + kernel[3][4] ~^ image[3][6] + kernel[4][0] ~^ image[4][2] + kernel[4][1] ~^ image[4][3] + kernel[4][2] ~^ image[4][4] + kernel[4][3] ~^ image[4][5] + kernel[4][4] ~^ image[4][6];
assign out_fmap[0][3] = kernel[0][0] ~^ image[0][3] + kernel[0][1] ~^ image[0][4] + kernel[0][2] ~^ image[0][5] + kernel[0][3] ~^ image[0][6] + kernel[0][4] ~^ image[0][7] + kernel[1][0] ~^ image[1][3] + kernel[1][1] ~^ image[1][4] + kernel[1][2] ~^ image[1][5] + kernel[1][3] ~^ image[1][6] + kernel[1][4] ~^ image[1][7] + kernel[2][0] ~^ image[2][3] + kernel[2][1] ~^ image[2][4] + kernel[2][2] ~^ image[2][5] + kernel[2][3] ~^ image[2][6] + kernel[2][4] ~^ image[2][7] + kernel[3][0] ~^ image[3][3] + kernel[3][1] ~^ image[3][4] + kernel[3][2] ~^ image[3][5] + kernel[3][3] ~^ image[3][6] + kernel[3][4] ~^ image[3][7] + kernel[4][0] ~^ image[4][3] + kernel[4][1] ~^ image[4][4] + kernel[4][2] ~^ image[4][5] + kernel[4][3] ~^ image[4][6] + kernel[4][4] ~^ image[4][7];
assign out_fmap[0][4] = kernel[0][0] ~^ image[0][4] + kernel[0][1] ~^ image[0][5] + kernel[0][2] ~^ image[0][6] + kernel[0][3] ~^ image[0][7] + kernel[0][4] ~^ image[0][8] + kernel[1][0] ~^ image[1][4] + kernel[1][1] ~^ image[1][5] + kernel[1][2] ~^ image[1][6] + kernel[1][3] ~^ image[1][7] + kernel[1][4] ~^ image[1][8] + kernel[2][0] ~^ image[2][4] + kernel[2][1] ~^ image[2][5] + kernel[2][2] ~^ image[2][6] + kernel[2][3] ~^ image[2][7] + kernel[2][4] ~^ image[2][8] + kernel[3][0] ~^ image[3][4] + kernel[3][1] ~^ image[3][5] + kernel[3][2] ~^ image[3][6] + kernel[3][3] ~^ image[3][7] + kernel[3][4] ~^ image[3][8] + kernel[4][0] ~^ image[4][4] + kernel[4][1] ~^ image[4][5] + kernel[4][2] ~^ image[4][6] + kernel[4][3] ~^ image[4][7] + kernel[4][4] ~^ image[4][8];
assign out_fmap[0][5] = kernel[0][0] ~^ image[0][5] + kernel[0][1] ~^ image[0][6] + kernel[0][2] ~^ image[0][7] + kernel[0][3] ~^ image[0][8] + kernel[0][4] ~^ image[0][9] + kernel[1][0] ~^ image[1][5] + kernel[1][1] ~^ image[1][6] + kernel[1][2] ~^ image[1][7] + kernel[1][3] ~^ image[1][8] + kernel[1][4] ~^ image[1][9] + kernel[2][0] ~^ image[2][5] + kernel[2][1] ~^ image[2][6] + kernel[2][2] ~^ image[2][7] + kernel[2][3] ~^ image[2][8] + kernel[2][4] ~^ image[2][9] + kernel[3][0] ~^ image[3][5] + kernel[3][1] ~^ image[3][6] + kernel[3][2] ~^ image[3][7] + kernel[3][3] ~^ image[3][8] + kernel[3][4] ~^ image[3][9] + kernel[4][0] ~^ image[4][5] + kernel[4][1] ~^ image[4][6] + kernel[4][2] ~^ image[4][7] + kernel[4][3] ~^ image[4][8] + kernel[4][4] ~^ image[4][9];
assign out_fmap[0][6] = kernel[0][0] ~^ image[0][6] + kernel[0][1] ~^ image[0][7] + kernel[0][2] ~^ image[0][8] + kernel[0][3] ~^ image[0][9] + kernel[0][4] ~^ image[0][10] + kernel[1][0] ~^ image[1][6] + kernel[1][1] ~^ image[1][7] + kernel[1][2] ~^ image[1][8] + kernel[1][3] ~^ image[1][9] + kernel[1][4] ~^ image[1][10] + kernel[2][0] ~^ image[2][6] + kernel[2][1] ~^ image[2][7] + kernel[2][2] ~^ image[2][8] + kernel[2][3] ~^ image[2][9] + kernel[2][4] ~^ image[2][10] + kernel[3][0] ~^ image[3][6] + kernel[3][1] ~^ image[3][7] + kernel[3][2] ~^ image[3][8] + kernel[3][3] ~^ image[3][9] + kernel[3][4] ~^ image[3][10] + kernel[4][0] ~^ image[4][6] + kernel[4][1] ~^ image[4][7] + kernel[4][2] ~^ image[4][8] + kernel[4][3] ~^ image[4][9] + kernel[4][4] ~^ image[4][10];
assign out_fmap[0][7] = kernel[0][0] ~^ image[0][7] + kernel[0][1] ~^ image[0][8] + kernel[0][2] ~^ image[0][9] + kernel[0][3] ~^ image[0][10] + kernel[0][4] ~^ image[0][11] + kernel[1][0] ~^ image[1][7] + kernel[1][1] ~^ image[1][8] + kernel[1][2] ~^ image[1][9] + kernel[1][3] ~^ image[1][10] + kernel[1][4] ~^ image[1][11] + kernel[2][0] ~^ image[2][7] + kernel[2][1] ~^ image[2][8] + kernel[2][2] ~^ image[2][9] + kernel[2][3] ~^ image[2][10] + kernel[2][4] ~^ image[2][11] + kernel[3][0] ~^ image[3][7] + kernel[3][1] ~^ image[3][8] + kernel[3][2] ~^ image[3][9] + kernel[3][3] ~^ image[3][10] + kernel[3][4] ~^ image[3][11] + kernel[4][0] ~^ image[4][7] + kernel[4][1] ~^ image[4][8] + kernel[4][2] ~^ image[4][9] + kernel[4][3] ~^ image[4][10] + kernel[4][4] ~^ image[4][11];
assign out_fmap[1][0] = kernel[0][0] ~^ image[1][0] + kernel[0][1] ~^ image[1][1] + kernel[0][2] ~^ image[1][2] + kernel[0][3] ~^ image[1][3] + kernel[0][4] ~^ image[1][4] + kernel[1][0] ~^ image[2][0] + kernel[1][1] ~^ image[2][1] + kernel[1][2] ~^ image[2][2] + kernel[1][3] ~^ image[2][3] + kernel[1][4] ~^ image[2][4] + kernel[2][0] ~^ image[3][0] + kernel[2][1] ~^ image[3][1] + kernel[2][2] ~^ image[3][2] + kernel[2][3] ~^ image[3][3] + kernel[2][4] ~^ image[3][4] + kernel[3][0] ~^ image[4][0] + kernel[3][1] ~^ image[4][1] + kernel[3][2] ~^ image[4][2] + kernel[3][3] ~^ image[4][3] + kernel[3][4] ~^ image[4][4] + kernel[4][0] ~^ image[5][0] + kernel[4][1] ~^ image[5][1] + kernel[4][2] ~^ image[5][2] + kernel[4][3] ~^ image[5][3] + kernel[4][4] ~^ image[5][4];
assign out_fmap[1][1] = kernel[0][0] ~^ image[1][1] + kernel[0][1] ~^ image[1][2] + kernel[0][2] ~^ image[1][3] + kernel[0][3] ~^ image[1][4] + kernel[0][4] ~^ image[1][5] + kernel[1][0] ~^ image[2][1] + kernel[1][1] ~^ image[2][2] + kernel[1][2] ~^ image[2][3] + kernel[1][3] ~^ image[2][4] + kernel[1][4] ~^ image[2][5] + kernel[2][0] ~^ image[3][1] + kernel[2][1] ~^ image[3][2] + kernel[2][2] ~^ image[3][3] + kernel[2][3] ~^ image[3][4] + kernel[2][4] ~^ image[3][5] + kernel[3][0] ~^ image[4][1] + kernel[3][1] ~^ image[4][2] + kernel[3][2] ~^ image[4][3] + kernel[3][3] ~^ image[4][4] + kernel[3][4] ~^ image[4][5] + kernel[4][0] ~^ image[5][1] + kernel[4][1] ~^ image[5][2] + kernel[4][2] ~^ image[5][3] + kernel[4][3] ~^ image[5][4] + kernel[4][4] ~^ image[5][5];
assign out_fmap[1][2] = kernel[0][0] ~^ image[1][2] + kernel[0][1] ~^ image[1][3] + kernel[0][2] ~^ image[1][4] + kernel[0][3] ~^ image[1][5] + kernel[0][4] ~^ image[1][6] + kernel[1][0] ~^ image[2][2] + kernel[1][1] ~^ image[2][3] + kernel[1][2] ~^ image[2][4] + kernel[1][3] ~^ image[2][5] + kernel[1][4] ~^ image[2][6] + kernel[2][0] ~^ image[3][2] + kernel[2][1] ~^ image[3][3] + kernel[2][2] ~^ image[3][4] + kernel[2][3] ~^ image[3][5] + kernel[2][4] ~^ image[3][6] + kernel[3][0] ~^ image[4][2] + kernel[3][1] ~^ image[4][3] + kernel[3][2] ~^ image[4][4] + kernel[3][3] ~^ image[4][5] + kernel[3][4] ~^ image[4][6] + kernel[4][0] ~^ image[5][2] + kernel[4][1] ~^ image[5][3] + kernel[4][2] ~^ image[5][4] + kernel[4][3] ~^ image[5][5] + kernel[4][4] ~^ image[5][6];
assign out_fmap[1][3] = kernel[0][0] ~^ image[1][3] + kernel[0][1] ~^ image[1][4] + kernel[0][2] ~^ image[1][5] + kernel[0][3] ~^ image[1][6] + kernel[0][4] ~^ image[1][7] + kernel[1][0] ~^ image[2][3] + kernel[1][1] ~^ image[2][4] + kernel[1][2] ~^ image[2][5] + kernel[1][3] ~^ image[2][6] + kernel[1][4] ~^ image[2][7] + kernel[2][0] ~^ image[3][3] + kernel[2][1] ~^ image[3][4] + kernel[2][2] ~^ image[3][5] + kernel[2][3] ~^ image[3][6] + kernel[2][4] ~^ image[3][7] + kernel[3][0] ~^ image[4][3] + kernel[3][1] ~^ image[4][4] + kernel[3][2] ~^ image[4][5] + kernel[3][3] ~^ image[4][6] + kernel[3][4] ~^ image[4][7] + kernel[4][0] ~^ image[5][3] + kernel[4][1] ~^ image[5][4] + kernel[4][2] ~^ image[5][5] + kernel[4][3] ~^ image[5][6] + kernel[4][4] ~^ image[5][7];
assign out_fmap[1][4] = kernel[0][0] ~^ image[1][4] + kernel[0][1] ~^ image[1][5] + kernel[0][2] ~^ image[1][6] + kernel[0][3] ~^ image[1][7] + kernel[0][4] ~^ image[1][8] + kernel[1][0] ~^ image[2][4] + kernel[1][1] ~^ image[2][5] + kernel[1][2] ~^ image[2][6] + kernel[1][3] ~^ image[2][7] + kernel[1][4] ~^ image[2][8] + kernel[2][0] ~^ image[3][4] + kernel[2][1] ~^ image[3][5] + kernel[2][2] ~^ image[3][6] + kernel[2][3] ~^ image[3][7] + kernel[2][4] ~^ image[3][8] + kernel[3][0] ~^ image[4][4] + kernel[3][1] ~^ image[4][5] + kernel[3][2] ~^ image[4][6] + kernel[3][3] ~^ image[4][7] + kernel[3][4] ~^ image[4][8] + kernel[4][0] ~^ image[5][4] + kernel[4][1] ~^ image[5][5] + kernel[4][2] ~^ image[5][6] + kernel[4][3] ~^ image[5][7] + kernel[4][4] ~^ image[5][8];
assign out_fmap[1][5] = kernel[0][0] ~^ image[1][5] + kernel[0][1] ~^ image[1][6] + kernel[0][2] ~^ image[1][7] + kernel[0][3] ~^ image[1][8] + kernel[0][4] ~^ image[1][9] + kernel[1][0] ~^ image[2][5] + kernel[1][1] ~^ image[2][6] + kernel[1][2] ~^ image[2][7] + kernel[1][3] ~^ image[2][8] + kernel[1][4] ~^ image[2][9] + kernel[2][0] ~^ image[3][5] + kernel[2][1] ~^ image[3][6] + kernel[2][2] ~^ image[3][7] + kernel[2][3] ~^ image[3][8] + kernel[2][4] ~^ image[3][9] + kernel[3][0] ~^ image[4][5] + kernel[3][1] ~^ image[4][6] + kernel[3][2] ~^ image[4][7] + kernel[3][3] ~^ image[4][8] + kernel[3][4] ~^ image[4][9] + kernel[4][0] ~^ image[5][5] + kernel[4][1] ~^ image[5][6] + kernel[4][2] ~^ image[5][7] + kernel[4][3] ~^ image[5][8] + kernel[4][4] ~^ image[5][9];
assign out_fmap[1][6] = kernel[0][0] ~^ image[1][6] + kernel[0][1] ~^ image[1][7] + kernel[0][2] ~^ image[1][8] + kernel[0][3] ~^ image[1][9] + kernel[0][4] ~^ image[1][10] + kernel[1][0] ~^ image[2][6] + kernel[1][1] ~^ image[2][7] + kernel[1][2] ~^ image[2][8] + kernel[1][3] ~^ image[2][9] + kernel[1][4] ~^ image[2][10] + kernel[2][0] ~^ image[3][6] + kernel[2][1] ~^ image[3][7] + kernel[2][2] ~^ image[3][8] + kernel[2][3] ~^ image[3][9] + kernel[2][4] ~^ image[3][10] + kernel[3][0] ~^ image[4][6] + kernel[3][1] ~^ image[4][7] + kernel[3][2] ~^ image[4][8] + kernel[3][3] ~^ image[4][9] + kernel[3][4] ~^ image[4][10] + kernel[4][0] ~^ image[5][6] + kernel[4][1] ~^ image[5][7] + kernel[4][2] ~^ image[5][8] + kernel[4][3] ~^ image[5][9] + kernel[4][4] ~^ image[5][10];
assign out_fmap[1][7] = kernel[0][0] ~^ image[1][7] + kernel[0][1] ~^ image[1][8] + kernel[0][2] ~^ image[1][9] + kernel[0][3] ~^ image[1][10] + kernel[0][4] ~^ image[1][11] + kernel[1][0] ~^ image[2][7] + kernel[1][1] ~^ image[2][8] + kernel[1][2] ~^ image[2][9] + kernel[1][3] ~^ image[2][10] + kernel[1][4] ~^ image[2][11] + kernel[2][0] ~^ image[3][7] + kernel[2][1] ~^ image[3][8] + kernel[2][2] ~^ image[3][9] + kernel[2][3] ~^ image[3][10] + kernel[2][4] ~^ image[3][11] + kernel[3][0] ~^ image[4][7] + kernel[3][1] ~^ image[4][8] + kernel[3][2] ~^ image[4][9] + kernel[3][3] ~^ image[4][10] + kernel[3][4] ~^ image[4][11] + kernel[4][0] ~^ image[5][7] + kernel[4][1] ~^ image[5][8] + kernel[4][2] ~^ image[5][9] + kernel[4][3] ~^ image[5][10] + kernel[4][4] ~^ image[5][11];
assign out_fmap[2][0] = kernel[0][0] ~^ image[2][0] + kernel[0][1] ~^ image[2][1] + kernel[0][2] ~^ image[2][2] + kernel[0][3] ~^ image[2][3] + kernel[0][4] ~^ image[2][4] + kernel[1][0] ~^ image[3][0] + kernel[1][1] ~^ image[3][1] + kernel[1][2] ~^ image[3][2] + kernel[1][3] ~^ image[3][3] + kernel[1][4] ~^ image[3][4] + kernel[2][0] ~^ image[4][0] + kernel[2][1] ~^ image[4][1] + kernel[2][2] ~^ image[4][2] + kernel[2][3] ~^ image[4][3] + kernel[2][4] ~^ image[4][4] + kernel[3][0] ~^ image[5][0] + kernel[3][1] ~^ image[5][1] + kernel[3][2] ~^ image[5][2] + kernel[3][3] ~^ image[5][3] + kernel[3][4] ~^ image[5][4] + kernel[4][0] ~^ image[6][0] + kernel[4][1] ~^ image[6][1] + kernel[4][2] ~^ image[6][2] + kernel[4][3] ~^ image[6][3] + kernel[4][4] ~^ image[6][4];
assign out_fmap[2][1] = kernel[0][0] ~^ image[2][1] + kernel[0][1] ~^ image[2][2] + kernel[0][2] ~^ image[2][3] + kernel[0][3] ~^ image[2][4] + kernel[0][4] ~^ image[2][5] + kernel[1][0] ~^ image[3][1] + kernel[1][1] ~^ image[3][2] + kernel[1][2] ~^ image[3][3] + kernel[1][3] ~^ image[3][4] + kernel[1][4] ~^ image[3][5] + kernel[2][0] ~^ image[4][1] + kernel[2][1] ~^ image[4][2] + kernel[2][2] ~^ image[4][3] + kernel[2][3] ~^ image[4][4] + kernel[2][4] ~^ image[4][5] + kernel[3][0] ~^ image[5][1] + kernel[3][1] ~^ image[5][2] + kernel[3][2] ~^ image[5][3] + kernel[3][3] ~^ image[5][4] + kernel[3][4] ~^ image[5][5] + kernel[4][0] ~^ image[6][1] + kernel[4][1] ~^ image[6][2] + kernel[4][2] ~^ image[6][3] + kernel[4][3] ~^ image[6][4] + kernel[4][4] ~^ image[6][5];
assign out_fmap[2][2] = kernel[0][0] ~^ image[2][2] + kernel[0][1] ~^ image[2][3] + kernel[0][2] ~^ image[2][4] + kernel[0][3] ~^ image[2][5] + kernel[0][4] ~^ image[2][6] + kernel[1][0] ~^ image[3][2] + kernel[1][1] ~^ image[3][3] + kernel[1][2] ~^ image[3][4] + kernel[1][3] ~^ image[3][5] + kernel[1][4] ~^ image[3][6] + kernel[2][0] ~^ image[4][2] + kernel[2][1] ~^ image[4][3] + kernel[2][2] ~^ image[4][4] + kernel[2][3] ~^ image[4][5] + kernel[2][4] ~^ image[4][6] + kernel[3][0] ~^ image[5][2] + kernel[3][1] ~^ image[5][3] + kernel[3][2] ~^ image[5][4] + kernel[3][3] ~^ image[5][5] + kernel[3][4] ~^ image[5][6] + kernel[4][0] ~^ image[6][2] + kernel[4][1] ~^ image[6][3] + kernel[4][2] ~^ image[6][4] + kernel[4][3] ~^ image[6][5] + kernel[4][4] ~^ image[6][6];
assign out_fmap[2][3] = kernel[0][0] ~^ image[2][3] + kernel[0][1] ~^ image[2][4] + kernel[0][2] ~^ image[2][5] + kernel[0][3] ~^ image[2][6] + kernel[0][4] ~^ image[2][7] + kernel[1][0] ~^ image[3][3] + kernel[1][1] ~^ image[3][4] + kernel[1][2] ~^ image[3][5] + kernel[1][3] ~^ image[3][6] + kernel[1][4] ~^ image[3][7] + kernel[2][0] ~^ image[4][3] + kernel[2][1] ~^ image[4][4] + kernel[2][2] ~^ image[4][5] + kernel[2][3] ~^ image[4][6] + kernel[2][4] ~^ image[4][7] + kernel[3][0] ~^ image[5][3] + kernel[3][1] ~^ image[5][4] + kernel[3][2] ~^ image[5][5] + kernel[3][3] ~^ image[5][6] + kernel[3][4] ~^ image[5][7] + kernel[4][0] ~^ image[6][3] + kernel[4][1] ~^ image[6][4] + kernel[4][2] ~^ image[6][5] + kernel[4][3] ~^ image[6][6] + kernel[4][4] ~^ image[6][7];
assign out_fmap[2][4] = kernel[0][0] ~^ image[2][4] + kernel[0][1] ~^ image[2][5] + kernel[0][2] ~^ image[2][6] + kernel[0][3] ~^ image[2][7] + kernel[0][4] ~^ image[2][8] + kernel[1][0] ~^ image[3][4] + kernel[1][1] ~^ image[3][5] + kernel[1][2] ~^ image[3][6] + kernel[1][3] ~^ image[3][7] + kernel[1][4] ~^ image[3][8] + kernel[2][0] ~^ image[4][4] + kernel[2][1] ~^ image[4][5] + kernel[2][2] ~^ image[4][6] + kernel[2][3] ~^ image[4][7] + kernel[2][4] ~^ image[4][8] + kernel[3][0] ~^ image[5][4] + kernel[3][1] ~^ image[5][5] + kernel[3][2] ~^ image[5][6] + kernel[3][3] ~^ image[5][7] + kernel[3][4] ~^ image[5][8] + kernel[4][0] ~^ image[6][4] + kernel[4][1] ~^ image[6][5] + kernel[4][2] ~^ image[6][6] + kernel[4][3] ~^ image[6][7] + kernel[4][4] ~^ image[6][8];
assign out_fmap[2][5] = kernel[0][0] ~^ image[2][5] + kernel[0][1] ~^ image[2][6] + kernel[0][2] ~^ image[2][7] + kernel[0][3] ~^ image[2][8] + kernel[0][4] ~^ image[2][9] + kernel[1][0] ~^ image[3][5] + kernel[1][1] ~^ image[3][6] + kernel[1][2] ~^ image[3][7] + kernel[1][3] ~^ image[3][8] + kernel[1][4] ~^ image[3][9] + kernel[2][0] ~^ image[4][5] + kernel[2][1] ~^ image[4][6] + kernel[2][2] ~^ image[4][7] + kernel[2][3] ~^ image[4][8] + kernel[2][4] ~^ image[4][9] + kernel[3][0] ~^ image[5][5] + kernel[3][1] ~^ image[5][6] + kernel[3][2] ~^ image[5][7] + kernel[3][3] ~^ image[5][8] + kernel[3][4] ~^ image[5][9] + kernel[4][0] ~^ image[6][5] + kernel[4][1] ~^ image[6][6] + kernel[4][2] ~^ image[6][7] + kernel[4][3] ~^ image[6][8] + kernel[4][4] ~^ image[6][9];
assign out_fmap[2][6] = kernel[0][0] ~^ image[2][6] + kernel[0][1] ~^ image[2][7] + kernel[0][2] ~^ image[2][8] + kernel[0][3] ~^ image[2][9] + kernel[0][4] ~^ image[2][10] + kernel[1][0] ~^ image[3][6] + kernel[1][1] ~^ image[3][7] + kernel[1][2] ~^ image[3][8] + kernel[1][3] ~^ image[3][9] + kernel[1][4] ~^ image[3][10] + kernel[2][0] ~^ image[4][6] + kernel[2][1] ~^ image[4][7] + kernel[2][2] ~^ image[4][8] + kernel[2][3] ~^ image[4][9] + kernel[2][4] ~^ image[4][10] + kernel[3][0] ~^ image[5][6] + kernel[3][1] ~^ image[5][7] + kernel[3][2] ~^ image[5][8] + kernel[3][3] ~^ image[5][9] + kernel[3][4] ~^ image[5][10] + kernel[4][0] ~^ image[6][6] + kernel[4][1] ~^ image[6][7] + kernel[4][2] ~^ image[6][8] + kernel[4][3] ~^ image[6][9] + kernel[4][4] ~^ image[6][10];
assign out_fmap[2][7] = kernel[0][0] ~^ image[2][7] + kernel[0][1] ~^ image[2][8] + kernel[0][2] ~^ image[2][9] + kernel[0][3] ~^ image[2][10] + kernel[0][4] ~^ image[2][11] + kernel[1][0] ~^ image[3][7] + kernel[1][1] ~^ image[3][8] + kernel[1][2] ~^ image[3][9] + kernel[1][3] ~^ image[3][10] + kernel[1][4] ~^ image[3][11] + kernel[2][0] ~^ image[4][7] + kernel[2][1] ~^ image[4][8] + kernel[2][2] ~^ image[4][9] + kernel[2][3] ~^ image[4][10] + kernel[2][4] ~^ image[4][11] + kernel[3][0] ~^ image[5][7] + kernel[3][1] ~^ image[5][8] + kernel[3][2] ~^ image[5][9] + kernel[3][3] ~^ image[5][10] + kernel[3][4] ~^ image[5][11] + kernel[4][0] ~^ image[6][7] + kernel[4][1] ~^ image[6][8] + kernel[4][2] ~^ image[6][9] + kernel[4][3] ~^ image[6][10] + kernel[4][4] ~^ image[6][11];
assign out_fmap[3][0] = kernel[0][0] ~^ image[3][0] + kernel[0][1] ~^ image[3][1] + kernel[0][2] ~^ image[3][2] + kernel[0][3] ~^ image[3][3] + kernel[0][4] ~^ image[3][4] + kernel[1][0] ~^ image[4][0] + kernel[1][1] ~^ image[4][1] + kernel[1][2] ~^ image[4][2] + kernel[1][3] ~^ image[4][3] + kernel[1][4] ~^ image[4][4] + kernel[2][0] ~^ image[5][0] + kernel[2][1] ~^ image[5][1] + kernel[2][2] ~^ image[5][2] + kernel[2][3] ~^ image[5][3] + kernel[2][4] ~^ image[5][4] + kernel[3][0] ~^ image[6][0] + kernel[3][1] ~^ image[6][1] + kernel[3][2] ~^ image[6][2] + kernel[3][3] ~^ image[6][3] + kernel[3][4] ~^ image[6][4] + kernel[4][0] ~^ image[7][0] + kernel[4][1] ~^ image[7][1] + kernel[4][2] ~^ image[7][2] + kernel[4][3] ~^ image[7][3] + kernel[4][4] ~^ image[7][4];
assign out_fmap[3][1] = kernel[0][0] ~^ image[3][1] + kernel[0][1] ~^ image[3][2] + kernel[0][2] ~^ image[3][3] + kernel[0][3] ~^ image[3][4] + kernel[0][4] ~^ image[3][5] + kernel[1][0] ~^ image[4][1] + kernel[1][1] ~^ image[4][2] + kernel[1][2] ~^ image[4][3] + kernel[1][3] ~^ image[4][4] + kernel[1][4] ~^ image[4][5] + kernel[2][0] ~^ image[5][1] + kernel[2][1] ~^ image[5][2] + kernel[2][2] ~^ image[5][3] + kernel[2][3] ~^ image[5][4] + kernel[2][4] ~^ image[5][5] + kernel[3][0] ~^ image[6][1] + kernel[3][1] ~^ image[6][2] + kernel[3][2] ~^ image[6][3] + kernel[3][3] ~^ image[6][4] + kernel[3][4] ~^ image[6][5] + kernel[4][0] ~^ image[7][1] + kernel[4][1] ~^ image[7][2] + kernel[4][2] ~^ image[7][3] + kernel[4][3] ~^ image[7][4] + kernel[4][4] ~^ image[7][5];
assign out_fmap[3][2] = kernel[0][0] ~^ image[3][2] + kernel[0][1] ~^ image[3][3] + kernel[0][2] ~^ image[3][4] + kernel[0][3] ~^ image[3][5] + kernel[0][4] ~^ image[3][6] + kernel[1][0] ~^ image[4][2] + kernel[1][1] ~^ image[4][3] + kernel[1][2] ~^ image[4][4] + kernel[1][3] ~^ image[4][5] + kernel[1][4] ~^ image[4][6] + kernel[2][0] ~^ image[5][2] + kernel[2][1] ~^ image[5][3] + kernel[2][2] ~^ image[5][4] + kernel[2][3] ~^ image[5][5] + kernel[2][4] ~^ image[5][6] + kernel[3][0] ~^ image[6][2] + kernel[3][1] ~^ image[6][3] + kernel[3][2] ~^ image[6][4] + kernel[3][3] ~^ image[6][5] + kernel[3][4] ~^ image[6][6] + kernel[4][0] ~^ image[7][2] + kernel[4][1] ~^ image[7][3] + kernel[4][2] ~^ image[7][4] + kernel[4][3] ~^ image[7][5] + kernel[4][4] ~^ image[7][6];
assign out_fmap[3][3] = kernel[0][0] ~^ image[3][3] + kernel[0][1] ~^ image[3][4] + kernel[0][2] ~^ image[3][5] + kernel[0][3] ~^ image[3][6] + kernel[0][4] ~^ image[3][7] + kernel[1][0] ~^ image[4][3] + kernel[1][1] ~^ image[4][4] + kernel[1][2] ~^ image[4][5] + kernel[1][3] ~^ image[4][6] + kernel[1][4] ~^ image[4][7] + kernel[2][0] ~^ image[5][3] + kernel[2][1] ~^ image[5][4] + kernel[2][2] ~^ image[5][5] + kernel[2][3] ~^ image[5][6] + kernel[2][4] ~^ image[5][7] + kernel[3][0] ~^ image[6][3] + kernel[3][1] ~^ image[6][4] + kernel[3][2] ~^ image[6][5] + kernel[3][3] ~^ image[6][6] + kernel[3][4] ~^ image[6][7] + kernel[4][0] ~^ image[7][3] + kernel[4][1] ~^ image[7][4] + kernel[4][2] ~^ image[7][5] + kernel[4][3] ~^ image[7][6] + kernel[4][4] ~^ image[7][7];
assign out_fmap[3][4] = kernel[0][0] ~^ image[3][4] + kernel[0][1] ~^ image[3][5] + kernel[0][2] ~^ image[3][6] + kernel[0][3] ~^ image[3][7] + kernel[0][4] ~^ image[3][8] + kernel[1][0] ~^ image[4][4] + kernel[1][1] ~^ image[4][5] + kernel[1][2] ~^ image[4][6] + kernel[1][3] ~^ image[4][7] + kernel[1][4] ~^ image[4][8] + kernel[2][0] ~^ image[5][4] + kernel[2][1] ~^ image[5][5] + kernel[2][2] ~^ image[5][6] + kernel[2][3] ~^ image[5][7] + kernel[2][4] ~^ image[5][8] + kernel[3][0] ~^ image[6][4] + kernel[3][1] ~^ image[6][5] + kernel[3][2] ~^ image[6][6] + kernel[3][3] ~^ image[6][7] + kernel[3][4] ~^ image[6][8] + kernel[4][0] ~^ image[7][4] + kernel[4][1] ~^ image[7][5] + kernel[4][2] ~^ image[7][6] + kernel[4][3] ~^ image[7][7] + kernel[4][4] ~^ image[7][8];
assign out_fmap[3][5] = kernel[0][0] ~^ image[3][5] + kernel[0][1] ~^ image[3][6] + kernel[0][2] ~^ image[3][7] + kernel[0][3] ~^ image[3][8] + kernel[0][4] ~^ image[3][9] + kernel[1][0] ~^ image[4][5] + kernel[1][1] ~^ image[4][6] + kernel[1][2] ~^ image[4][7] + kernel[1][3] ~^ image[4][8] + kernel[1][4] ~^ image[4][9] + kernel[2][0] ~^ image[5][5] + kernel[2][1] ~^ image[5][6] + kernel[2][2] ~^ image[5][7] + kernel[2][3] ~^ image[5][8] + kernel[2][4] ~^ image[5][9] + kernel[3][0] ~^ image[6][5] + kernel[3][1] ~^ image[6][6] + kernel[3][2] ~^ image[6][7] + kernel[3][3] ~^ image[6][8] + kernel[3][4] ~^ image[6][9] + kernel[4][0] ~^ image[7][5] + kernel[4][1] ~^ image[7][6] + kernel[4][2] ~^ image[7][7] + kernel[4][3] ~^ image[7][8] + kernel[4][4] ~^ image[7][9];
assign out_fmap[3][6] = kernel[0][0] ~^ image[3][6] + kernel[0][1] ~^ image[3][7] + kernel[0][2] ~^ image[3][8] + kernel[0][3] ~^ image[3][9] + kernel[0][4] ~^ image[3][10] + kernel[1][0] ~^ image[4][6] + kernel[1][1] ~^ image[4][7] + kernel[1][2] ~^ image[4][8] + kernel[1][3] ~^ image[4][9] + kernel[1][4] ~^ image[4][10] + kernel[2][0] ~^ image[5][6] + kernel[2][1] ~^ image[5][7] + kernel[2][2] ~^ image[5][8] + kernel[2][3] ~^ image[5][9] + kernel[2][4] ~^ image[5][10] + kernel[3][0] ~^ image[6][6] + kernel[3][1] ~^ image[6][7] + kernel[3][2] ~^ image[6][8] + kernel[3][3] ~^ image[6][9] + kernel[3][4] ~^ image[6][10] + kernel[4][0] ~^ image[7][6] + kernel[4][1] ~^ image[7][7] + kernel[4][2] ~^ image[7][8] + kernel[4][3] ~^ image[7][9] + kernel[4][4] ~^ image[7][10];
assign out_fmap[3][7] = kernel[0][0] ~^ image[3][7] + kernel[0][1] ~^ image[3][8] + kernel[0][2] ~^ image[3][9] + kernel[0][3] ~^ image[3][10] + kernel[0][4] ~^ image[3][11] + kernel[1][0] ~^ image[4][7] + kernel[1][1] ~^ image[4][8] + kernel[1][2] ~^ image[4][9] + kernel[1][3] ~^ image[4][10] + kernel[1][4] ~^ image[4][11] + kernel[2][0] ~^ image[5][7] + kernel[2][1] ~^ image[5][8] + kernel[2][2] ~^ image[5][9] + kernel[2][3] ~^ image[5][10] + kernel[2][4] ~^ image[5][11] + kernel[3][0] ~^ image[6][7] + kernel[3][1] ~^ image[6][8] + kernel[3][2] ~^ image[6][9] + kernel[3][3] ~^ image[6][10] + kernel[3][4] ~^ image[6][11] + kernel[4][0] ~^ image[7][7] + kernel[4][1] ~^ image[7][8] + kernel[4][2] ~^ image[7][9] + kernel[4][3] ~^ image[7][10] + kernel[4][4] ~^ image[7][11];
assign out_fmap[4][0] = kernel[0][0] ~^ image[4][0] + kernel[0][1] ~^ image[4][1] + kernel[0][2] ~^ image[4][2] + kernel[0][3] ~^ image[4][3] + kernel[0][4] ~^ image[4][4] + kernel[1][0] ~^ image[5][0] + kernel[1][1] ~^ image[5][1] + kernel[1][2] ~^ image[5][2] + kernel[1][3] ~^ image[5][3] + kernel[1][4] ~^ image[5][4] + kernel[2][0] ~^ image[6][0] + kernel[2][1] ~^ image[6][1] + kernel[2][2] ~^ image[6][2] + kernel[2][3] ~^ image[6][3] + kernel[2][4] ~^ image[6][4] + kernel[3][0] ~^ image[7][0] + kernel[3][1] ~^ image[7][1] + kernel[3][2] ~^ image[7][2] + kernel[3][3] ~^ image[7][3] + kernel[3][4] ~^ image[7][4] + kernel[4][0] ~^ image[8][0] + kernel[4][1] ~^ image[8][1] + kernel[4][2] ~^ image[8][2] + kernel[4][3] ~^ image[8][3] + kernel[4][4] ~^ image[8][4];
assign out_fmap[4][1] = kernel[0][0] ~^ image[4][1] + kernel[0][1] ~^ image[4][2] + kernel[0][2] ~^ image[4][3] + kernel[0][3] ~^ image[4][4] + kernel[0][4] ~^ image[4][5] + kernel[1][0] ~^ image[5][1] + kernel[1][1] ~^ image[5][2] + kernel[1][2] ~^ image[5][3] + kernel[1][3] ~^ image[5][4] + kernel[1][4] ~^ image[5][5] + kernel[2][0] ~^ image[6][1] + kernel[2][1] ~^ image[6][2] + kernel[2][2] ~^ image[6][3] + kernel[2][3] ~^ image[6][4] + kernel[2][4] ~^ image[6][5] + kernel[3][0] ~^ image[7][1] + kernel[3][1] ~^ image[7][2] + kernel[3][2] ~^ image[7][3] + kernel[3][3] ~^ image[7][4] + kernel[3][4] ~^ image[7][5] + kernel[4][0] ~^ image[8][1] + kernel[4][1] ~^ image[8][2] + kernel[4][2] ~^ image[8][3] + kernel[4][3] ~^ image[8][4] + kernel[4][4] ~^ image[8][5];
assign out_fmap[4][2] = kernel[0][0] ~^ image[4][2] + kernel[0][1] ~^ image[4][3] + kernel[0][2] ~^ image[4][4] + kernel[0][3] ~^ image[4][5] + kernel[0][4] ~^ image[4][6] + kernel[1][0] ~^ image[5][2] + kernel[1][1] ~^ image[5][3] + kernel[1][2] ~^ image[5][4] + kernel[1][3] ~^ image[5][5] + kernel[1][4] ~^ image[5][6] + kernel[2][0] ~^ image[6][2] + kernel[2][1] ~^ image[6][3] + kernel[2][2] ~^ image[6][4] + kernel[2][3] ~^ image[6][5] + kernel[2][4] ~^ image[6][6] + kernel[3][0] ~^ image[7][2] + kernel[3][1] ~^ image[7][3] + kernel[3][2] ~^ image[7][4] + kernel[3][3] ~^ image[7][5] + kernel[3][4] ~^ image[7][6] + kernel[4][0] ~^ image[8][2] + kernel[4][1] ~^ image[8][3] + kernel[4][2] ~^ image[8][4] + kernel[4][3] ~^ image[8][5] + kernel[4][4] ~^ image[8][6];
assign out_fmap[4][3] = kernel[0][0] ~^ image[4][3] + kernel[0][1] ~^ image[4][4] + kernel[0][2] ~^ image[4][5] + kernel[0][3] ~^ image[4][6] + kernel[0][4] ~^ image[4][7] + kernel[1][0] ~^ image[5][3] + kernel[1][1] ~^ image[5][4] + kernel[1][2] ~^ image[5][5] + kernel[1][3] ~^ image[5][6] + kernel[1][4] ~^ image[5][7] + kernel[2][0] ~^ image[6][3] + kernel[2][1] ~^ image[6][4] + kernel[2][2] ~^ image[6][5] + kernel[2][3] ~^ image[6][6] + kernel[2][4] ~^ image[6][7] + kernel[3][0] ~^ image[7][3] + kernel[3][1] ~^ image[7][4] + kernel[3][2] ~^ image[7][5] + kernel[3][3] ~^ image[7][6] + kernel[3][4] ~^ image[7][7] + kernel[4][0] ~^ image[8][3] + kernel[4][1] ~^ image[8][4] + kernel[4][2] ~^ image[8][5] + kernel[4][3] ~^ image[8][6] + kernel[4][4] ~^ image[8][7];
assign out_fmap[4][4] = kernel[0][0] ~^ image[4][4] + kernel[0][1] ~^ image[4][5] + kernel[0][2] ~^ image[4][6] + kernel[0][3] ~^ image[4][7] + kernel[0][4] ~^ image[4][8] + kernel[1][0] ~^ image[5][4] + kernel[1][1] ~^ image[5][5] + kernel[1][2] ~^ image[5][6] + kernel[1][3] ~^ image[5][7] + kernel[1][4] ~^ image[5][8] + kernel[2][0] ~^ image[6][4] + kernel[2][1] ~^ image[6][5] + kernel[2][2] ~^ image[6][6] + kernel[2][3] ~^ image[6][7] + kernel[2][4] ~^ image[6][8] + kernel[3][0] ~^ image[7][4] + kernel[3][1] ~^ image[7][5] + kernel[3][2] ~^ image[7][6] + kernel[3][3] ~^ image[7][7] + kernel[3][4] ~^ image[7][8] + kernel[4][0] ~^ image[8][4] + kernel[4][1] ~^ image[8][5] + kernel[4][2] ~^ image[8][6] + kernel[4][3] ~^ image[8][7] + kernel[4][4] ~^ image[8][8];
assign out_fmap[4][5] = kernel[0][0] ~^ image[4][5] + kernel[0][1] ~^ image[4][6] + kernel[0][2] ~^ image[4][7] + kernel[0][3] ~^ image[4][8] + kernel[0][4] ~^ image[4][9] + kernel[1][0] ~^ image[5][5] + kernel[1][1] ~^ image[5][6] + kernel[1][2] ~^ image[5][7] + kernel[1][3] ~^ image[5][8] + kernel[1][4] ~^ image[5][9] + kernel[2][0] ~^ image[6][5] + kernel[2][1] ~^ image[6][6] + kernel[2][2] ~^ image[6][7] + kernel[2][3] ~^ image[6][8] + kernel[2][4] ~^ image[6][9] + kernel[3][0] ~^ image[7][5] + kernel[3][1] ~^ image[7][6] + kernel[3][2] ~^ image[7][7] + kernel[3][3] ~^ image[7][8] + kernel[3][4] ~^ image[7][9] + kernel[4][0] ~^ image[8][5] + kernel[4][1] ~^ image[8][6] + kernel[4][2] ~^ image[8][7] + kernel[4][3] ~^ image[8][8] + kernel[4][4] ~^ image[8][9];
assign out_fmap[4][6] = kernel[0][0] ~^ image[4][6] + kernel[0][1] ~^ image[4][7] + kernel[0][2] ~^ image[4][8] + kernel[0][3] ~^ image[4][9] + kernel[0][4] ~^ image[4][10] + kernel[1][0] ~^ image[5][6] + kernel[1][1] ~^ image[5][7] + kernel[1][2] ~^ image[5][8] + kernel[1][3] ~^ image[5][9] + kernel[1][4] ~^ image[5][10] + kernel[2][0] ~^ image[6][6] + kernel[2][1] ~^ image[6][7] + kernel[2][2] ~^ image[6][8] + kernel[2][3] ~^ image[6][9] + kernel[2][4] ~^ image[6][10] + kernel[3][0] ~^ image[7][6] + kernel[3][1] ~^ image[7][7] + kernel[3][2] ~^ image[7][8] + kernel[3][3] ~^ image[7][9] + kernel[3][4] ~^ image[7][10] + kernel[4][0] ~^ image[8][6] + kernel[4][1] ~^ image[8][7] + kernel[4][2] ~^ image[8][8] + kernel[4][3] ~^ image[8][9] + kernel[4][4] ~^ image[8][10];
assign out_fmap[4][7] = kernel[0][0] ~^ image[4][7] + kernel[0][1] ~^ image[4][8] + kernel[0][2] ~^ image[4][9] + kernel[0][3] ~^ image[4][10] + kernel[0][4] ~^ image[4][11] + kernel[1][0] ~^ image[5][7] + kernel[1][1] ~^ image[5][8] + kernel[1][2] ~^ image[5][9] + kernel[1][3] ~^ image[5][10] + kernel[1][4] ~^ image[5][11] + kernel[2][0] ~^ image[6][7] + kernel[2][1] ~^ image[6][8] + kernel[2][2] ~^ image[6][9] + kernel[2][3] ~^ image[6][10] + kernel[2][4] ~^ image[6][11] + kernel[3][0] ~^ image[7][7] + kernel[3][1] ~^ image[7][8] + kernel[3][2] ~^ image[7][9] + kernel[3][3] ~^ image[7][10] + kernel[3][4] ~^ image[7][11] + kernel[4][0] ~^ image[8][7] + kernel[4][1] ~^ image[8][8] + kernel[4][2] ~^ image[8][9] + kernel[4][3] ~^ image[8][10] + kernel[4][4] ~^ image[8][11];
assign out_fmap[5][0] = kernel[0][0] ~^ image[5][0] + kernel[0][1] ~^ image[5][1] + kernel[0][2] ~^ image[5][2] + kernel[0][3] ~^ image[5][3] + kernel[0][4] ~^ image[5][4] + kernel[1][0] ~^ image[6][0] + kernel[1][1] ~^ image[6][1] + kernel[1][2] ~^ image[6][2] + kernel[1][3] ~^ image[6][3] + kernel[1][4] ~^ image[6][4] + kernel[2][0] ~^ image[7][0] + kernel[2][1] ~^ image[7][1] + kernel[2][2] ~^ image[7][2] + kernel[2][3] ~^ image[7][3] + kernel[2][4] ~^ image[7][4] + kernel[3][0] ~^ image[8][0] + kernel[3][1] ~^ image[8][1] + kernel[3][2] ~^ image[8][2] + kernel[3][3] ~^ image[8][3] + kernel[3][4] ~^ image[8][4] + kernel[4][0] ~^ image[9][0] + kernel[4][1] ~^ image[9][1] + kernel[4][2] ~^ image[9][2] + kernel[4][3] ~^ image[9][3] + kernel[4][4] ~^ image[9][4];
assign out_fmap[5][1] = kernel[0][0] ~^ image[5][1] + kernel[0][1] ~^ image[5][2] + kernel[0][2] ~^ image[5][3] + kernel[0][3] ~^ image[5][4] + kernel[0][4] ~^ image[5][5] + kernel[1][0] ~^ image[6][1] + kernel[1][1] ~^ image[6][2] + kernel[1][2] ~^ image[6][3] + kernel[1][3] ~^ image[6][4] + kernel[1][4] ~^ image[6][5] + kernel[2][0] ~^ image[7][1] + kernel[2][1] ~^ image[7][2] + kernel[2][2] ~^ image[7][3] + kernel[2][3] ~^ image[7][4] + kernel[2][4] ~^ image[7][5] + kernel[3][0] ~^ image[8][1] + kernel[3][1] ~^ image[8][2] + kernel[3][2] ~^ image[8][3] + kernel[3][3] ~^ image[8][4] + kernel[3][4] ~^ image[8][5] + kernel[4][0] ~^ image[9][1] + kernel[4][1] ~^ image[9][2] + kernel[4][2] ~^ image[9][3] + kernel[4][3] ~^ image[9][4] + kernel[4][4] ~^ image[9][5];
assign out_fmap[5][2] = kernel[0][0] ~^ image[5][2] + kernel[0][1] ~^ image[5][3] + kernel[0][2] ~^ image[5][4] + kernel[0][3] ~^ image[5][5] + kernel[0][4] ~^ image[5][6] + kernel[1][0] ~^ image[6][2] + kernel[1][1] ~^ image[6][3] + kernel[1][2] ~^ image[6][4] + kernel[1][3] ~^ image[6][5] + kernel[1][4] ~^ image[6][6] + kernel[2][0] ~^ image[7][2] + kernel[2][1] ~^ image[7][3] + kernel[2][2] ~^ image[7][4] + kernel[2][3] ~^ image[7][5] + kernel[2][4] ~^ image[7][6] + kernel[3][0] ~^ image[8][2] + kernel[3][1] ~^ image[8][3] + kernel[3][2] ~^ image[8][4] + kernel[3][3] ~^ image[8][5] + kernel[3][4] ~^ image[8][6] + kernel[4][0] ~^ image[9][2] + kernel[4][1] ~^ image[9][3] + kernel[4][2] ~^ image[9][4] + kernel[4][3] ~^ image[9][5] + kernel[4][4] ~^ image[9][6];
assign out_fmap[5][3] = kernel[0][0] ~^ image[5][3] + kernel[0][1] ~^ image[5][4] + kernel[0][2] ~^ image[5][5] + kernel[0][3] ~^ image[5][6] + kernel[0][4] ~^ image[5][7] + kernel[1][0] ~^ image[6][3] + kernel[1][1] ~^ image[6][4] + kernel[1][2] ~^ image[6][5] + kernel[1][3] ~^ image[6][6] + kernel[1][4] ~^ image[6][7] + kernel[2][0] ~^ image[7][3] + kernel[2][1] ~^ image[7][4] + kernel[2][2] ~^ image[7][5] + kernel[2][3] ~^ image[7][6] + kernel[2][4] ~^ image[7][7] + kernel[3][0] ~^ image[8][3] + kernel[3][1] ~^ image[8][4] + kernel[3][2] ~^ image[8][5] + kernel[3][3] ~^ image[8][6] + kernel[3][4] ~^ image[8][7] + kernel[4][0] ~^ image[9][3] + kernel[4][1] ~^ image[9][4] + kernel[4][2] ~^ image[9][5] + kernel[4][3] ~^ image[9][6] + kernel[4][4] ~^ image[9][7];
assign out_fmap[5][4] = kernel[0][0] ~^ image[5][4] + kernel[0][1] ~^ image[5][5] + kernel[0][2] ~^ image[5][6] + kernel[0][3] ~^ image[5][7] + kernel[0][4] ~^ image[5][8] + kernel[1][0] ~^ image[6][4] + kernel[1][1] ~^ image[6][5] + kernel[1][2] ~^ image[6][6] + kernel[1][3] ~^ image[6][7] + kernel[1][4] ~^ image[6][8] + kernel[2][0] ~^ image[7][4] + kernel[2][1] ~^ image[7][5] + kernel[2][2] ~^ image[7][6] + kernel[2][3] ~^ image[7][7] + kernel[2][4] ~^ image[7][8] + kernel[3][0] ~^ image[8][4] + kernel[3][1] ~^ image[8][5] + kernel[3][2] ~^ image[8][6] + kernel[3][3] ~^ image[8][7] + kernel[3][4] ~^ image[8][8] + kernel[4][0] ~^ image[9][4] + kernel[4][1] ~^ image[9][5] + kernel[4][2] ~^ image[9][6] + kernel[4][3] ~^ image[9][7] + kernel[4][4] ~^ image[9][8];
assign out_fmap[5][5] = kernel[0][0] ~^ image[5][5] + kernel[0][1] ~^ image[5][6] + kernel[0][2] ~^ image[5][7] + kernel[0][3] ~^ image[5][8] + kernel[0][4] ~^ image[5][9] + kernel[1][0] ~^ image[6][5] + kernel[1][1] ~^ image[6][6] + kernel[1][2] ~^ image[6][7] + kernel[1][3] ~^ image[6][8] + kernel[1][4] ~^ image[6][9] + kernel[2][0] ~^ image[7][5] + kernel[2][1] ~^ image[7][6] + kernel[2][2] ~^ image[7][7] + kernel[2][3] ~^ image[7][8] + kernel[2][4] ~^ image[7][9] + kernel[3][0] ~^ image[8][5] + kernel[3][1] ~^ image[8][6] + kernel[3][2] ~^ image[8][7] + kernel[3][3] ~^ image[8][8] + kernel[3][4] ~^ image[8][9] + kernel[4][0] ~^ image[9][5] + kernel[4][1] ~^ image[9][6] + kernel[4][2] ~^ image[9][7] + kernel[4][3] ~^ image[9][8] + kernel[4][4] ~^ image[9][9];
assign out_fmap[5][6] = kernel[0][0] ~^ image[5][6] + kernel[0][1] ~^ image[5][7] + kernel[0][2] ~^ image[5][8] + kernel[0][3] ~^ image[5][9] + kernel[0][4] ~^ image[5][10] + kernel[1][0] ~^ image[6][6] + kernel[1][1] ~^ image[6][7] + kernel[1][2] ~^ image[6][8] + kernel[1][3] ~^ image[6][9] + kernel[1][4] ~^ image[6][10] + kernel[2][0] ~^ image[7][6] + kernel[2][1] ~^ image[7][7] + kernel[2][2] ~^ image[7][8] + kernel[2][3] ~^ image[7][9] + kernel[2][4] ~^ image[7][10] + kernel[3][0] ~^ image[8][6] + kernel[3][1] ~^ image[8][7] + kernel[3][2] ~^ image[8][8] + kernel[3][3] ~^ image[8][9] + kernel[3][4] ~^ image[8][10] + kernel[4][0] ~^ image[9][6] + kernel[4][1] ~^ image[9][7] + kernel[4][2] ~^ image[9][8] + kernel[4][3] ~^ image[9][9] + kernel[4][4] ~^ image[9][10];
assign out_fmap[5][7] = kernel[0][0] ~^ image[5][7] + kernel[0][1] ~^ image[5][8] + kernel[0][2] ~^ image[5][9] + kernel[0][3] ~^ image[5][10] + kernel[0][4] ~^ image[5][11] + kernel[1][0] ~^ image[6][7] + kernel[1][1] ~^ image[6][8] + kernel[1][2] ~^ image[6][9] + kernel[1][3] ~^ image[6][10] + kernel[1][4] ~^ image[6][11] + kernel[2][0] ~^ image[7][7] + kernel[2][1] ~^ image[7][8] + kernel[2][2] ~^ image[7][9] + kernel[2][3] ~^ image[7][10] + kernel[2][4] ~^ image[7][11] + kernel[3][0] ~^ image[8][7] + kernel[3][1] ~^ image[8][8] + kernel[3][2] ~^ image[8][9] + kernel[3][3] ~^ image[8][10] + kernel[3][4] ~^ image[8][11] + kernel[4][0] ~^ image[9][7] + kernel[4][1] ~^ image[9][8] + kernel[4][2] ~^ image[9][9] + kernel[4][3] ~^ image[9][10] + kernel[4][4] ~^ image[9][11];
assign out_fmap[6][0] = kernel[0][0] ~^ image[6][0] + kernel[0][1] ~^ image[6][1] + kernel[0][2] ~^ image[6][2] + kernel[0][3] ~^ image[6][3] + kernel[0][4] ~^ image[6][4] + kernel[1][0] ~^ image[7][0] + kernel[1][1] ~^ image[7][1] + kernel[1][2] ~^ image[7][2] + kernel[1][3] ~^ image[7][3] + kernel[1][4] ~^ image[7][4] + kernel[2][0] ~^ image[8][0] + kernel[2][1] ~^ image[8][1] + kernel[2][2] ~^ image[8][2] + kernel[2][3] ~^ image[8][3] + kernel[2][4] ~^ image[8][4] + kernel[3][0] ~^ image[9][0] + kernel[3][1] ~^ image[9][1] + kernel[3][2] ~^ image[9][2] + kernel[3][3] ~^ image[9][3] + kernel[3][4] ~^ image[9][4] + kernel[4][0] ~^ image[10][0] + kernel[4][1] ~^ image[10][1] + kernel[4][2] ~^ image[10][2] + kernel[4][3] ~^ image[10][3] + kernel[4][4] ~^ image[10][4];
assign out_fmap[6][1] = kernel[0][0] ~^ image[6][1] + kernel[0][1] ~^ image[6][2] + kernel[0][2] ~^ image[6][3] + kernel[0][3] ~^ image[6][4] + kernel[0][4] ~^ image[6][5] + kernel[1][0] ~^ image[7][1] + kernel[1][1] ~^ image[7][2] + kernel[1][2] ~^ image[7][3] + kernel[1][3] ~^ image[7][4] + kernel[1][4] ~^ image[7][5] + kernel[2][0] ~^ image[8][1] + kernel[2][1] ~^ image[8][2] + kernel[2][2] ~^ image[8][3] + kernel[2][3] ~^ image[8][4] + kernel[2][4] ~^ image[8][5] + kernel[3][0] ~^ image[9][1] + kernel[3][1] ~^ image[9][2] + kernel[3][2] ~^ image[9][3] + kernel[3][3] ~^ image[9][4] + kernel[3][4] ~^ image[9][5] + kernel[4][0] ~^ image[10][1] + kernel[4][1] ~^ image[10][2] + kernel[4][2] ~^ image[10][3] + kernel[4][3] ~^ image[10][4] + kernel[4][4] ~^ image[10][5];
assign out_fmap[6][2] = kernel[0][0] ~^ image[6][2] + kernel[0][1] ~^ image[6][3] + kernel[0][2] ~^ image[6][4] + kernel[0][3] ~^ image[6][5] + kernel[0][4] ~^ image[6][6] + kernel[1][0] ~^ image[7][2] + kernel[1][1] ~^ image[7][3] + kernel[1][2] ~^ image[7][4] + kernel[1][3] ~^ image[7][5] + kernel[1][4] ~^ image[7][6] + kernel[2][0] ~^ image[8][2] + kernel[2][1] ~^ image[8][3] + kernel[2][2] ~^ image[8][4] + kernel[2][3] ~^ image[8][5] + kernel[2][4] ~^ image[8][6] + kernel[3][0] ~^ image[9][2] + kernel[3][1] ~^ image[9][3] + kernel[3][2] ~^ image[9][4] + kernel[3][3] ~^ image[9][5] + kernel[3][4] ~^ image[9][6] + kernel[4][0] ~^ image[10][2] + kernel[4][1] ~^ image[10][3] + kernel[4][2] ~^ image[10][4] + kernel[4][3] ~^ image[10][5] + kernel[4][4] ~^ image[10][6];
assign out_fmap[6][3] = kernel[0][0] ~^ image[6][3] + kernel[0][1] ~^ image[6][4] + kernel[0][2] ~^ image[6][5] + kernel[0][3] ~^ image[6][6] + kernel[0][4] ~^ image[6][7] + kernel[1][0] ~^ image[7][3] + kernel[1][1] ~^ image[7][4] + kernel[1][2] ~^ image[7][5] + kernel[1][3] ~^ image[7][6] + kernel[1][4] ~^ image[7][7] + kernel[2][0] ~^ image[8][3] + kernel[2][1] ~^ image[8][4] + kernel[2][2] ~^ image[8][5] + kernel[2][3] ~^ image[8][6] + kernel[2][4] ~^ image[8][7] + kernel[3][0] ~^ image[9][3] + kernel[3][1] ~^ image[9][4] + kernel[3][2] ~^ image[9][5] + kernel[3][3] ~^ image[9][6] + kernel[3][4] ~^ image[9][7] + kernel[4][0] ~^ image[10][3] + kernel[4][1] ~^ image[10][4] + kernel[4][2] ~^ image[10][5] + kernel[4][3] ~^ image[10][6] + kernel[4][4] ~^ image[10][7];
assign out_fmap[6][4] = kernel[0][0] ~^ image[6][4] + kernel[0][1] ~^ image[6][5] + kernel[0][2] ~^ image[6][6] + kernel[0][3] ~^ image[6][7] + kernel[0][4] ~^ image[6][8] + kernel[1][0] ~^ image[7][4] + kernel[1][1] ~^ image[7][5] + kernel[1][2] ~^ image[7][6] + kernel[1][3] ~^ image[7][7] + kernel[1][4] ~^ image[7][8] + kernel[2][0] ~^ image[8][4] + kernel[2][1] ~^ image[8][5] + kernel[2][2] ~^ image[8][6] + kernel[2][3] ~^ image[8][7] + kernel[2][4] ~^ image[8][8] + kernel[3][0] ~^ image[9][4] + kernel[3][1] ~^ image[9][5] + kernel[3][2] ~^ image[9][6] + kernel[3][3] ~^ image[9][7] + kernel[3][4] ~^ image[9][8] + kernel[4][0] ~^ image[10][4] + kernel[4][1] ~^ image[10][5] + kernel[4][2] ~^ image[10][6] + kernel[4][3] ~^ image[10][7] + kernel[4][4] ~^ image[10][8];
assign out_fmap[6][5] = kernel[0][0] ~^ image[6][5] + kernel[0][1] ~^ image[6][6] + kernel[0][2] ~^ image[6][7] + kernel[0][3] ~^ image[6][8] + kernel[0][4] ~^ image[6][9] + kernel[1][0] ~^ image[7][5] + kernel[1][1] ~^ image[7][6] + kernel[1][2] ~^ image[7][7] + kernel[1][3] ~^ image[7][8] + kernel[1][4] ~^ image[7][9] + kernel[2][0] ~^ image[8][5] + kernel[2][1] ~^ image[8][6] + kernel[2][2] ~^ image[8][7] + kernel[2][3] ~^ image[8][8] + kernel[2][4] ~^ image[8][9] + kernel[3][0] ~^ image[9][5] + kernel[3][1] ~^ image[9][6] + kernel[3][2] ~^ image[9][7] + kernel[3][3] ~^ image[9][8] + kernel[3][4] ~^ image[9][9] + kernel[4][0] ~^ image[10][5] + kernel[4][1] ~^ image[10][6] + kernel[4][2] ~^ image[10][7] + kernel[4][3] ~^ image[10][8] + kernel[4][4] ~^ image[10][9];
assign out_fmap[6][6] = kernel[0][0] ~^ image[6][6] + kernel[0][1] ~^ image[6][7] + kernel[0][2] ~^ image[6][8] + kernel[0][3] ~^ image[6][9] + kernel[0][4] ~^ image[6][10] + kernel[1][0] ~^ image[7][6] + kernel[1][1] ~^ image[7][7] + kernel[1][2] ~^ image[7][8] + kernel[1][3] ~^ image[7][9] + kernel[1][4] ~^ image[7][10] + kernel[2][0] ~^ image[8][6] + kernel[2][1] ~^ image[8][7] + kernel[2][2] ~^ image[8][8] + kernel[2][3] ~^ image[8][9] + kernel[2][4] ~^ image[8][10] + kernel[3][0] ~^ image[9][6] + kernel[3][1] ~^ image[9][7] + kernel[3][2] ~^ image[9][8] + kernel[3][3] ~^ image[9][9] + kernel[3][4] ~^ image[9][10] + kernel[4][0] ~^ image[10][6] + kernel[4][1] ~^ image[10][7] + kernel[4][2] ~^ image[10][8] + kernel[4][3] ~^ image[10][9] + kernel[4][4] ~^ image[10][10];
assign out_fmap[6][7] = kernel[0][0] ~^ image[6][7] + kernel[0][1] ~^ image[6][8] + kernel[0][2] ~^ image[6][9] + kernel[0][3] ~^ image[6][10] + kernel[0][4] ~^ image[6][11] + kernel[1][0] ~^ image[7][7] + kernel[1][1] ~^ image[7][8] + kernel[1][2] ~^ image[7][9] + kernel[1][3] ~^ image[7][10] + kernel[1][4] ~^ image[7][11] + kernel[2][0] ~^ image[8][7] + kernel[2][1] ~^ image[8][8] + kernel[2][2] ~^ image[8][9] + kernel[2][3] ~^ image[8][10] + kernel[2][4] ~^ image[8][11] + kernel[3][0] ~^ image[9][7] + kernel[3][1] ~^ image[9][8] + kernel[3][2] ~^ image[9][9] + kernel[3][3] ~^ image[9][10] + kernel[3][4] ~^ image[9][11] + kernel[4][0] ~^ image[10][7] + kernel[4][1] ~^ image[10][8] + kernel[4][2] ~^ image[10][9] + kernel[4][3] ~^ image[10][10] + kernel[4][4] ~^ image[10][11];
assign out_fmap[7][0] = kernel[0][0] ~^ image[7][0] + kernel[0][1] ~^ image[7][1] + kernel[0][2] ~^ image[7][2] + kernel[0][3] ~^ image[7][3] + kernel[0][4] ~^ image[7][4] + kernel[1][0] ~^ image[8][0] + kernel[1][1] ~^ image[8][1] + kernel[1][2] ~^ image[8][2] + kernel[1][3] ~^ image[8][3] + kernel[1][4] ~^ image[8][4] + kernel[2][0] ~^ image[9][0] + kernel[2][1] ~^ image[9][1] + kernel[2][2] ~^ image[9][2] + kernel[2][3] ~^ image[9][3] + kernel[2][4] ~^ image[9][4] + kernel[3][0] ~^ image[10][0] + kernel[3][1] ~^ image[10][1] + kernel[3][2] ~^ image[10][2] + kernel[3][3] ~^ image[10][3] + kernel[3][4] ~^ image[10][4] + kernel[4][0] ~^ image[11][0] + kernel[4][1] ~^ image[11][1] + kernel[4][2] ~^ image[11][2] + kernel[4][3] ~^ image[11][3] + kernel[4][4] ~^ image[11][4];
assign out_fmap[7][1] = kernel[0][0] ~^ image[7][1] + kernel[0][1] ~^ image[7][2] + kernel[0][2] ~^ image[7][3] + kernel[0][3] ~^ image[7][4] + kernel[0][4] ~^ image[7][5] + kernel[1][0] ~^ image[8][1] + kernel[1][1] ~^ image[8][2] + kernel[1][2] ~^ image[8][3] + kernel[1][3] ~^ image[8][4] + kernel[1][4] ~^ image[8][5] + kernel[2][0] ~^ image[9][1] + kernel[2][1] ~^ image[9][2] + kernel[2][2] ~^ image[9][3] + kernel[2][3] ~^ image[9][4] + kernel[2][4] ~^ image[9][5] + kernel[3][0] ~^ image[10][1] + kernel[3][1] ~^ image[10][2] + kernel[3][2] ~^ image[10][3] + kernel[3][3] ~^ image[10][4] + kernel[3][4] ~^ image[10][5] + kernel[4][0] ~^ image[11][1] + kernel[4][1] ~^ image[11][2] + kernel[4][2] ~^ image[11][3] + kernel[4][3] ~^ image[11][4] + kernel[4][4] ~^ image[11][5];
assign out_fmap[7][2] = kernel[0][0] ~^ image[7][2] + kernel[0][1] ~^ image[7][3] + kernel[0][2] ~^ image[7][4] + kernel[0][3] ~^ image[7][5] + kernel[0][4] ~^ image[7][6] + kernel[1][0] ~^ image[8][2] + kernel[1][1] ~^ image[8][3] + kernel[1][2] ~^ image[8][4] + kernel[1][3] ~^ image[8][5] + kernel[1][4] ~^ image[8][6] + kernel[2][0] ~^ image[9][2] + kernel[2][1] ~^ image[9][3] + kernel[2][2] ~^ image[9][4] + kernel[2][3] ~^ image[9][5] + kernel[2][4] ~^ image[9][6] + kernel[3][0] ~^ image[10][2] + kernel[3][1] ~^ image[10][3] + kernel[3][2] ~^ image[10][4] + kernel[3][3] ~^ image[10][5] + kernel[3][4] ~^ image[10][6] + kernel[4][0] ~^ image[11][2] + kernel[4][1] ~^ image[11][3] + kernel[4][2] ~^ image[11][4] + kernel[4][3] ~^ image[11][5] + kernel[4][4] ~^ image[11][6];
assign out_fmap[7][3] = kernel[0][0] ~^ image[7][3] + kernel[0][1] ~^ image[7][4] + kernel[0][2] ~^ image[7][5] + kernel[0][3] ~^ image[7][6] + kernel[0][4] ~^ image[7][7] + kernel[1][0] ~^ image[8][3] + kernel[1][1] ~^ image[8][4] + kernel[1][2] ~^ image[8][5] + kernel[1][3] ~^ image[8][6] + kernel[1][4] ~^ image[8][7] + kernel[2][0] ~^ image[9][3] + kernel[2][1] ~^ image[9][4] + kernel[2][2] ~^ image[9][5] + kernel[2][3] ~^ image[9][6] + kernel[2][4] ~^ image[9][7] + kernel[3][0] ~^ image[10][3] + kernel[3][1] ~^ image[10][4] + kernel[3][2] ~^ image[10][5] + kernel[3][3] ~^ image[10][6] + kernel[3][4] ~^ image[10][7] + kernel[4][0] ~^ image[11][3] + kernel[4][1] ~^ image[11][4] + kernel[4][2] ~^ image[11][5] + kernel[4][3] ~^ image[11][6] + kernel[4][4] ~^ image[11][7];
assign out_fmap[7][4] = kernel[0][0] ~^ image[7][4] + kernel[0][1] ~^ image[7][5] + kernel[0][2] ~^ image[7][6] + kernel[0][3] ~^ image[7][7] + kernel[0][4] ~^ image[7][8] + kernel[1][0] ~^ image[8][4] + kernel[1][1] ~^ image[8][5] + kernel[1][2] ~^ image[8][6] + kernel[1][3] ~^ image[8][7] + kernel[1][4] ~^ image[8][8] + kernel[2][0] ~^ image[9][4] + kernel[2][1] ~^ image[9][5] + kernel[2][2] ~^ image[9][6] + kernel[2][3] ~^ image[9][7] + kernel[2][4] ~^ image[9][8] + kernel[3][0] ~^ image[10][4] + kernel[3][1] ~^ image[10][5] + kernel[3][2] ~^ image[10][6] + kernel[3][3] ~^ image[10][7] + kernel[3][4] ~^ image[10][8] + kernel[4][0] ~^ image[11][4] + kernel[4][1] ~^ image[11][5] + kernel[4][2] ~^ image[11][6] + kernel[4][3] ~^ image[11][7] + kernel[4][4] ~^ image[11][8];
assign out_fmap[7][5] = kernel[0][0] ~^ image[7][5] + kernel[0][1] ~^ image[7][6] + kernel[0][2] ~^ image[7][7] + kernel[0][3] ~^ image[7][8] + kernel[0][4] ~^ image[7][9] + kernel[1][0] ~^ image[8][5] + kernel[1][1] ~^ image[8][6] + kernel[1][2] ~^ image[8][7] + kernel[1][3] ~^ image[8][8] + kernel[1][4] ~^ image[8][9] + kernel[2][0] ~^ image[9][5] + kernel[2][1] ~^ image[9][6] + kernel[2][2] ~^ image[9][7] + kernel[2][3] ~^ image[9][8] + kernel[2][4] ~^ image[9][9] + kernel[3][0] ~^ image[10][5] + kernel[3][1] ~^ image[10][6] + kernel[3][2] ~^ image[10][7] + kernel[3][3] ~^ image[10][8] + kernel[3][4] ~^ image[10][9] + kernel[4][0] ~^ image[11][5] + kernel[4][1] ~^ image[11][6] + kernel[4][2] ~^ image[11][7] + kernel[4][3] ~^ image[11][8] + kernel[4][4] ~^ image[11][9];
assign out_fmap[7][6] = kernel[0][0] ~^ image[7][6] + kernel[0][1] ~^ image[7][7] + kernel[0][2] ~^ image[7][8] + kernel[0][3] ~^ image[7][9] + kernel[0][4] ~^ image[7][10] + kernel[1][0] ~^ image[8][6] + kernel[1][1] ~^ image[8][7] + kernel[1][2] ~^ image[8][8] + kernel[1][3] ~^ image[8][9] + kernel[1][4] ~^ image[8][10] + kernel[2][0] ~^ image[9][6] + kernel[2][1] ~^ image[9][7] + kernel[2][2] ~^ image[9][8] + kernel[2][3] ~^ image[9][9] + kernel[2][4] ~^ image[9][10] + kernel[3][0] ~^ image[10][6] + kernel[3][1] ~^ image[10][7] + kernel[3][2] ~^ image[10][8] + kernel[3][3] ~^ image[10][9] + kernel[3][4] ~^ image[10][10] + kernel[4][0] ~^ image[11][6] + kernel[4][1] ~^ image[11][7] + kernel[4][2] ~^ image[11][8] + kernel[4][3] ~^ image[11][9] + kernel[4][4] ~^ image[11][10];
assign out_fmap[7][7] = kernel[0][0] ~^ image[7][7] + kernel[0][1] ~^ image[7][8] + kernel[0][2] ~^ image[7][9] + kernel[0][3] ~^ image[7][10] + kernel[0][4] ~^ image[7][11] + kernel[1][0] ~^ image[8][7] + kernel[1][1] ~^ image[8][8] + kernel[1][2] ~^ image[8][9] + kernel[1][3] ~^ image[8][10] + kernel[1][4] ~^ image[8][11] + kernel[2][0] ~^ image[9][7] + kernel[2][1] ~^ image[9][8] + kernel[2][2] ~^ image[9][9] + kernel[2][3] ~^ image[9][10] + kernel[2][4] ~^ image[9][11] + kernel[3][0] ~^ image[10][7] + kernel[3][1] ~^ image[10][8] + kernel[3][2] ~^ image[10][9] + kernel[3][3] ~^ image[10][10] + kernel[3][4] ~^ image[10][11] + kernel[4][0] ~^ image[11][7] + kernel[4][1] ~^ image[11][8] + kernel[4][2] ~^ image[11][9] + kernel[4][3] ~^ image[11][10] + kernel[4][4] ~^ image[11][11];

endmodule