module conv_pool_pixel450
#(parameter chan = 18,
parameter bW = 9)
(
input logic image[0:chan*6*6-1],
input logic kernels[0:chan*5*5-1],
input logic [bW-1:0] offset,
output logic pixel);


logic [chan*5*5-1:0] image_slice1;
assign image_slice1 = {image[0*6*6+0*6+0],image[0*6*6+0*6+1],image[0*6*6+0*6+2],image[0*6*6+0*6+3],image[0*6*6+0*6+4],image[0*6*6+1*6+0],image[0*6*6+1*6+1],image[0*6*6+1*6+2],image[0*6*6+1*6+3],image[0*6*6+1*6+4],image[0*6*6+2*6+0],image[0*6*6+2*6+1],image[0*6*6+2*6+2],image[0*6*6+2*6+3],image[0*6*6+2*6+4],image[0*6*6+3*6+0],image[0*6*6+3*6+1],image[0*6*6+3*6+2],image[0*6*6+3*6+3],image[0*6*6+3*6+4],image[0*6*6+4*6+0],image[0*6*6+4*6+1],image[0*6*6+4*6+2],image[0*6*6+4*6+3],image[0*6*6+4*6+4],image[1*6*6+0*6+0],image[1*6*6+0*6+1],image[1*6*6+0*6+2],image[1*6*6+0*6+3],image[1*6*6+0*6+4],image[1*6*6+1*6+0],image[1*6*6+1*6+1],image[1*6*6+1*6+2],image[1*6*6+1*6+3],image[1*6*6+1*6+4],image[1*6*6+2*6+0],image[1*6*6+2*6+1],image[1*6*6+2*6+2],image[1*6*6+2*6+3],image[1*6*6+2*6+4],image[1*6*6+3*6+0],image[1*6*6+3*6+1],image[1*6*6+3*6+2],image[1*6*6+3*6+3],image[1*6*6+3*6+4],image[1*6*6+4*6+0],image[1*6*6+4*6+1],image[1*6*6+4*6+2],image[1*6*6+4*6+3],image[1*6*6+4*6+4],image[2*6*6+0*6+0],image[2*6*6+0*6+1],image[2*6*6+0*6+2],image[2*6*6+0*6+3],image[2*6*6+0*6+4],image[2*6*6+1*6+0],image[2*6*6+1*6+1],image[2*6*6+1*6+2],image[2*6*6+1*6+3],image[2*6*6+1*6+4],image[2*6*6+2*6+0],image[2*6*6+2*6+1],image[2*6*6+2*6+2],image[2*6*6+2*6+3],image[2*6*6+2*6+4],image[2*6*6+3*6+0],image[2*6*6+3*6+1],image[2*6*6+3*6+2],image[2*6*6+3*6+3],image[2*6*6+3*6+4],image[2*6*6+4*6+0],image[2*6*6+4*6+1],image[2*6*6+4*6+2],image[2*6*6+4*6+3],image[2*6*6+4*6+4],image[3*6*6+0*6+0],image[3*6*6+0*6+1],image[3*6*6+0*6+2],image[3*6*6+0*6+3],image[3*6*6+0*6+4],image[3*6*6+1*6+0],image[3*6*6+1*6+1],image[3*6*6+1*6+2],image[3*6*6+1*6+3],image[3*6*6+1*6+4],image[3*6*6+2*6+0],image[3*6*6+2*6+1],image[3*6*6+2*6+2],image[3*6*6+2*6+3],image[3*6*6+2*6+4],image[3*6*6+3*6+0],image[3*6*6+3*6+1],image[3*6*6+3*6+2],image[3*6*6+3*6+3],image[3*6*6+3*6+4],image[3*6*6+4*6+0],image[3*6*6+4*6+1],image[3*6*6+4*6+2],image[3*6*6+4*6+3],image[3*6*6+4*6+4],image[4*6*6+0*6+0],image[4*6*6+0*6+1],image[4*6*6+0*6+2],image[4*6*6+0*6+3],image[4*6*6+0*6+4],image[4*6*6+1*6+0],image[4*6*6+1*6+1],image[4*6*6+1*6+2],image[4*6*6+1*6+3],image[4*6*6+1*6+4],image[4*6*6+2*6+0],image[4*6*6+2*6+1],image[4*6*6+2*6+2],image[4*6*6+2*6+3],image[4*6*6+2*6+4],image[4*6*6+3*6+0],image[4*6*6+3*6+1],image[4*6*6+3*6+2],image[4*6*6+3*6+3],image[4*6*6+3*6+4],image[4*6*6+4*6+0],image[4*6*6+4*6+1],image[4*6*6+4*6+2],image[4*6*6+4*6+3],image[4*6*6+4*6+4],image[5*6*6+0*6+0],image[5*6*6+0*6+1],image[5*6*6+0*6+2],image[5*6*6+0*6+3],image[5*6*6+0*6+4],image[5*6*6+1*6+0],image[5*6*6+1*6+1],image[5*6*6+1*6+2],image[5*6*6+1*6+3],image[5*6*6+1*6+4],image[5*6*6+2*6+0],image[5*6*6+2*6+1],image[5*6*6+2*6+2],image[5*6*6+2*6+3],image[5*6*6+2*6+4],image[5*6*6+3*6+0],image[5*6*6+3*6+1],image[5*6*6+3*6+2],image[5*6*6+3*6+3],image[5*6*6+3*6+4],image[5*6*6+4*6+0],image[5*6*6+4*6+1],image[5*6*6+4*6+2],image[5*6*6+4*6+3],image[5*6*6+4*6+4],image[6*6*6+0*6+0],image[6*6*6+0*6+1],image[6*6*6+0*6+2],image[6*6*6+0*6+3],image[6*6*6+0*6+4],image[6*6*6+1*6+0],image[6*6*6+1*6+1],image[6*6*6+1*6+2],image[6*6*6+1*6+3],image[6*6*6+1*6+4],image[6*6*6+2*6+0],image[6*6*6+2*6+1],image[6*6*6+2*6+2],image[6*6*6+2*6+3],image[6*6*6+2*6+4],image[6*6*6+3*6+0],image[6*6*6+3*6+1],image[6*6*6+3*6+2],image[6*6*6+3*6+3],image[6*6*6+3*6+4],image[6*6*6+4*6+0],image[6*6*6+4*6+1],image[6*6*6+4*6+2],image[6*6*6+4*6+3],image[6*6*6+4*6+4],image[7*6*6+0*6+0],image[7*6*6+0*6+1],image[7*6*6+0*6+2],image[7*6*6+0*6+3],image[7*6*6+0*6+4],image[7*6*6+1*6+0],image[7*6*6+1*6+1],image[7*6*6+1*6+2],image[7*6*6+1*6+3],image[7*6*6+1*6+4],image[7*6*6+2*6+0],image[7*6*6+2*6+1],image[7*6*6+2*6+2],image[7*6*6+2*6+3],image[7*6*6+2*6+4],image[7*6*6+3*6+0],image[7*6*6+3*6+1],image[7*6*6+3*6+2],image[7*6*6+3*6+3],image[7*6*6+3*6+4],image[7*6*6+4*6+0],image[7*6*6+4*6+1],image[7*6*6+4*6+2],image[7*6*6+4*6+3],image[7*6*6+4*6+4],image[8*6*6+0*6+0],image[8*6*6+0*6+1],image[8*6*6+0*6+2],image[8*6*6+0*6+3],image[8*6*6+0*6+4],image[8*6*6+1*6+0],image[8*6*6+1*6+1],image[8*6*6+1*6+2],image[8*6*6+1*6+3],image[8*6*6+1*6+4],image[8*6*6+2*6+0],image[8*6*6+2*6+1],image[8*6*6+2*6+2],image[8*6*6+2*6+3],image[8*6*6+2*6+4],image[8*6*6+3*6+0],image[8*6*6+3*6+1],image[8*6*6+3*6+2],image[8*6*6+3*6+3],image[8*6*6+3*6+4],image[8*6*6+4*6+0],image[8*6*6+4*6+1],image[8*6*6+4*6+2],image[8*6*6+4*6+3],image[8*6*6+4*6+4],image[9*6*6+0*6+0],image[9*6*6+0*6+1],image[9*6*6+0*6+2],image[9*6*6+0*6+3],image[9*6*6+0*6+4],image[9*6*6+1*6+0],image[9*6*6+1*6+1],image[9*6*6+1*6+2],image[9*6*6+1*6+3],image[9*6*6+1*6+4],image[9*6*6+2*6+0],image[9*6*6+2*6+1],image[9*6*6+2*6+2],image[9*6*6+2*6+3],image[9*6*6+2*6+4],image[9*6*6+3*6+0],image[9*6*6+3*6+1],image[9*6*6+3*6+2],image[9*6*6+3*6+3],image[9*6*6+3*6+4],image[9*6*6+4*6+0],image[9*6*6+4*6+1],image[9*6*6+4*6+2],image[9*6*6+4*6+3],image[9*6*6+4*6+4],image[10*6*6+0*6+0],image[10*6*6+0*6+1],image[10*6*6+0*6+2],image[10*6*6+0*6+3],image[10*6*6+0*6+4],image[10*6*6+1*6+0],image[10*6*6+1*6+1],image[10*6*6+1*6+2],image[10*6*6+1*6+3],image[10*6*6+1*6+4],image[10*6*6+2*6+0],image[10*6*6+2*6+1],image[10*6*6+2*6+2],image[10*6*6+2*6+3],image[10*6*6+2*6+4],image[10*6*6+3*6+0],image[10*6*6+3*6+1],image[10*6*6+3*6+2],image[10*6*6+3*6+3],image[10*6*6+3*6+4],image[10*6*6+4*6+0],image[10*6*6+4*6+1],image[10*6*6+4*6+2],image[10*6*6+4*6+3],image[10*6*6+4*6+4],image[11*6*6+0*6+0],image[11*6*6+0*6+1],image[11*6*6+0*6+2],image[11*6*6+0*6+3],image[11*6*6+0*6+4],image[11*6*6+1*6+0],image[11*6*6+1*6+1],image[11*6*6+1*6+2],image[11*6*6+1*6+3],image[11*6*6+1*6+4],image[11*6*6+2*6+0],image[11*6*6+2*6+1],image[11*6*6+2*6+2],image[11*6*6+2*6+3],image[11*6*6+2*6+4],image[11*6*6+3*6+0],image[11*6*6+3*6+1],image[11*6*6+3*6+2],image[11*6*6+3*6+3],image[11*6*6+3*6+4],image[11*6*6+4*6+0],image[11*6*6+4*6+1],image[11*6*6+4*6+2],image[11*6*6+4*6+3],image[11*6*6+4*6+4],image[12*6*6+0*6+0],image[12*6*6+0*6+1],image[12*6*6+0*6+2],image[12*6*6+0*6+3],image[12*6*6+0*6+4],image[12*6*6+1*6+0],image[12*6*6+1*6+1],image[12*6*6+1*6+2],image[12*6*6+1*6+3],image[12*6*6+1*6+4],image[12*6*6+2*6+0],image[12*6*6+2*6+1],image[12*6*6+2*6+2],image[12*6*6+2*6+3],image[12*6*6+2*6+4],image[12*6*6+3*6+0],image[12*6*6+3*6+1],image[12*6*6+3*6+2],image[12*6*6+3*6+3],image[12*6*6+3*6+4],image[12*6*6+4*6+0],image[12*6*6+4*6+1],image[12*6*6+4*6+2],image[12*6*6+4*6+3],image[12*6*6+4*6+4],image[13*6*6+0*6+0],image[13*6*6+0*6+1],image[13*6*6+0*6+2],image[13*6*6+0*6+3],image[13*6*6+0*6+4],image[13*6*6+1*6+0],image[13*6*6+1*6+1],image[13*6*6+1*6+2],image[13*6*6+1*6+3],image[13*6*6+1*6+4],image[13*6*6+2*6+0],image[13*6*6+2*6+1],image[13*6*6+2*6+2],image[13*6*6+2*6+3],image[13*6*6+2*6+4],image[13*6*6+3*6+0],image[13*6*6+3*6+1],image[13*6*6+3*6+2],image[13*6*6+3*6+3],image[13*6*6+3*6+4],image[13*6*6+4*6+0],image[13*6*6+4*6+1],image[13*6*6+4*6+2],image[13*6*6+4*6+3],image[13*6*6+4*6+4],image[14*6*6+0*6+0],image[14*6*6+0*6+1],image[14*6*6+0*6+2],image[14*6*6+0*6+3],image[14*6*6+0*6+4],image[14*6*6+1*6+0],image[14*6*6+1*6+1],image[14*6*6+1*6+2],image[14*6*6+1*6+3],image[14*6*6+1*6+4],image[14*6*6+2*6+0],image[14*6*6+2*6+1],image[14*6*6+2*6+2],image[14*6*6+2*6+3],image[14*6*6+2*6+4],image[14*6*6+3*6+0],image[14*6*6+3*6+1],image[14*6*6+3*6+2],image[14*6*6+3*6+3],image[14*6*6+3*6+4],image[14*6*6+4*6+0],image[14*6*6+4*6+1],image[14*6*6+4*6+2],image[14*6*6+4*6+3],image[14*6*6+4*6+4],image[15*6*6+0*6+0],image[15*6*6+0*6+1],image[15*6*6+0*6+2],image[15*6*6+0*6+3],image[15*6*6+0*6+4],image[15*6*6+1*6+0],image[15*6*6+1*6+1],image[15*6*6+1*6+2],image[15*6*6+1*6+3],image[15*6*6+1*6+4],image[15*6*6+2*6+0],image[15*6*6+2*6+1],image[15*6*6+2*6+2],image[15*6*6+2*6+3],image[15*6*6+2*6+4],image[15*6*6+3*6+0],image[15*6*6+3*6+1],image[15*6*6+3*6+2],image[15*6*6+3*6+3],image[15*6*6+3*6+4],image[15*6*6+4*6+0],image[15*6*6+4*6+1],image[15*6*6+4*6+2],image[15*6*6+4*6+3],image[15*6*6+4*6+4],image[16*6*6+0*6+0],image[16*6*6+0*6+1],image[16*6*6+0*6+2],image[16*6*6+0*6+3],image[16*6*6+0*6+4],image[16*6*6+1*6+0],image[16*6*6+1*6+1],image[16*6*6+1*6+2],image[16*6*6+1*6+3],image[16*6*6+1*6+4],image[16*6*6+2*6+0],image[16*6*6+2*6+1],image[16*6*6+2*6+2],image[16*6*6+2*6+3],image[16*6*6+2*6+4],image[16*6*6+3*6+0],image[16*6*6+3*6+1],image[16*6*6+3*6+2],image[16*6*6+3*6+3],image[16*6*6+3*6+4],image[16*6*6+4*6+0],image[16*6*6+4*6+1],image[16*6*6+4*6+2],image[16*6*6+4*6+3],image[16*6*6+4*6+4],image[17*6*6+0*6+0],image[17*6*6+0*6+1],image[17*6*6+0*6+2],image[17*6*6+0*6+3],image[17*6*6+0*6+4],image[17*6*6+1*6+0],image[17*6*6+1*6+1],image[17*6*6+1*6+2],image[17*6*6+1*6+3],image[17*6*6+1*6+4],image[17*6*6+2*6+0],image[17*6*6+2*6+1],image[17*6*6+2*6+2],image[17*6*6+2*6+3],image[17*6*6+2*6+4],image[17*6*6+3*6+0],image[17*6*6+3*6+1],image[17*6*6+3*6+2],image[17*6*6+3*6+3],image[17*6*6+3*6+4],image[17*6*6+4*6+0],image[17*6*6+4*6+1],image[17*6*6+4*6+2],image[17*6*6+4*6+3],image[17*6*6+4*6+4]};
logic [chan*5*5-1:0] image_slice2;
assign image_slice2 = {image[0*6*6+0*6+1],image[0*6*6+0*6+2],image[0*6*6+0*6+3],image[0*6*6+0*6+4],image[0*6*6+0*6+5],image[0*6*6+1*6+1],image[0*6*6+1*6+2],image[0*6*6+1*6+3],image[0*6*6+1*6+4],image[0*6*6+1*6+5],image[0*6*6+2*6+1],image[0*6*6+2*6+2],image[0*6*6+2*6+3],image[0*6*6+2*6+4],image[0*6*6+2*6+5],image[0*6*6+3*6+1],image[0*6*6+3*6+2],image[0*6*6+3*6+3],image[0*6*6+3*6+4],image[0*6*6+3*6+5],image[0*6*6+4*6+1],image[0*6*6+4*6+2],image[0*6*6+4*6+3],image[0*6*6+4*6+4],image[0*6*6+4*6+5],image[1*6*6+0*6+1],image[1*6*6+0*6+2],image[1*6*6+0*6+3],image[1*6*6+0*6+4],image[1*6*6+0*6+5],image[1*6*6+1*6+1],image[1*6*6+1*6+2],image[1*6*6+1*6+3],image[1*6*6+1*6+4],image[1*6*6+1*6+5],image[1*6*6+2*6+1],image[1*6*6+2*6+2],image[1*6*6+2*6+3],image[1*6*6+2*6+4],image[1*6*6+2*6+5],image[1*6*6+3*6+1],image[1*6*6+3*6+2],image[1*6*6+3*6+3],image[1*6*6+3*6+4],image[1*6*6+3*6+5],image[1*6*6+4*6+1],image[1*6*6+4*6+2],image[1*6*6+4*6+3],image[1*6*6+4*6+4],image[1*6*6+4*6+5],image[2*6*6+0*6+1],image[2*6*6+0*6+2],image[2*6*6+0*6+3],image[2*6*6+0*6+4],image[2*6*6+0*6+5],image[2*6*6+1*6+1],image[2*6*6+1*6+2],image[2*6*6+1*6+3],image[2*6*6+1*6+4],image[2*6*6+1*6+5],image[2*6*6+2*6+1],image[2*6*6+2*6+2],image[2*6*6+2*6+3],image[2*6*6+2*6+4],image[2*6*6+2*6+5],image[2*6*6+3*6+1],image[2*6*6+3*6+2],image[2*6*6+3*6+3],image[2*6*6+3*6+4],image[2*6*6+3*6+5],image[2*6*6+4*6+1],image[2*6*6+4*6+2],image[2*6*6+4*6+3],image[2*6*6+4*6+4],image[2*6*6+4*6+5],image[3*6*6+0*6+1],image[3*6*6+0*6+2],image[3*6*6+0*6+3],image[3*6*6+0*6+4],image[3*6*6+0*6+5],image[3*6*6+1*6+1],image[3*6*6+1*6+2],image[3*6*6+1*6+3],image[3*6*6+1*6+4],image[3*6*6+1*6+5],image[3*6*6+2*6+1],image[3*6*6+2*6+2],image[3*6*6+2*6+3],image[3*6*6+2*6+4],image[3*6*6+2*6+5],image[3*6*6+3*6+1],image[3*6*6+3*6+2],image[3*6*6+3*6+3],image[3*6*6+3*6+4],image[3*6*6+3*6+5],image[3*6*6+4*6+1],image[3*6*6+4*6+2],image[3*6*6+4*6+3],image[3*6*6+4*6+4],image[3*6*6+4*6+5],image[4*6*6+0*6+1],image[4*6*6+0*6+2],image[4*6*6+0*6+3],image[4*6*6+0*6+4],image[4*6*6+0*6+5],image[4*6*6+1*6+1],image[4*6*6+1*6+2],image[4*6*6+1*6+3],image[4*6*6+1*6+4],image[4*6*6+1*6+5],image[4*6*6+2*6+1],image[4*6*6+2*6+2],image[4*6*6+2*6+3],image[4*6*6+2*6+4],image[4*6*6+2*6+5],image[4*6*6+3*6+1],image[4*6*6+3*6+2],image[4*6*6+3*6+3],image[4*6*6+3*6+4],image[4*6*6+3*6+5],image[4*6*6+4*6+1],image[4*6*6+4*6+2],image[4*6*6+4*6+3],image[4*6*6+4*6+4],image[4*6*6+4*6+5],image[5*6*6+0*6+1],image[5*6*6+0*6+2],image[5*6*6+0*6+3],image[5*6*6+0*6+4],image[5*6*6+0*6+5],image[5*6*6+1*6+1],image[5*6*6+1*6+2],image[5*6*6+1*6+3],image[5*6*6+1*6+4],image[5*6*6+1*6+5],image[5*6*6+2*6+1],image[5*6*6+2*6+2],image[5*6*6+2*6+3],image[5*6*6+2*6+4],image[5*6*6+2*6+5],image[5*6*6+3*6+1],image[5*6*6+3*6+2],image[5*6*6+3*6+3],image[5*6*6+3*6+4],image[5*6*6+3*6+5],image[5*6*6+4*6+1],image[5*6*6+4*6+2],image[5*6*6+4*6+3],image[5*6*6+4*6+4],image[5*6*6+4*6+5],image[6*6*6+0*6+1],image[6*6*6+0*6+2],image[6*6*6+0*6+3],image[6*6*6+0*6+4],image[6*6*6+0*6+5],image[6*6*6+1*6+1],image[6*6*6+1*6+2],image[6*6*6+1*6+3],image[6*6*6+1*6+4],image[6*6*6+1*6+5],image[6*6*6+2*6+1],image[6*6*6+2*6+2],image[6*6*6+2*6+3],image[6*6*6+2*6+4],image[6*6*6+2*6+5],image[6*6*6+3*6+1],image[6*6*6+3*6+2],image[6*6*6+3*6+3],image[6*6*6+3*6+4],image[6*6*6+3*6+5],image[6*6*6+4*6+1],image[6*6*6+4*6+2],image[6*6*6+4*6+3],image[6*6*6+4*6+4],image[6*6*6+4*6+5],image[7*6*6+0*6+1],image[7*6*6+0*6+2],image[7*6*6+0*6+3],image[7*6*6+0*6+4],image[7*6*6+0*6+5],image[7*6*6+1*6+1],image[7*6*6+1*6+2],image[7*6*6+1*6+3],image[7*6*6+1*6+4],image[7*6*6+1*6+5],image[7*6*6+2*6+1],image[7*6*6+2*6+2],image[7*6*6+2*6+3],image[7*6*6+2*6+4],image[7*6*6+2*6+5],image[7*6*6+3*6+1],image[7*6*6+3*6+2],image[7*6*6+3*6+3],image[7*6*6+3*6+4],image[7*6*6+3*6+5],image[7*6*6+4*6+1],image[7*6*6+4*6+2],image[7*6*6+4*6+3],image[7*6*6+4*6+4],image[7*6*6+4*6+5],image[8*6*6+0*6+1],image[8*6*6+0*6+2],image[8*6*6+0*6+3],image[8*6*6+0*6+4],image[8*6*6+0*6+5],image[8*6*6+1*6+1],image[8*6*6+1*6+2],image[8*6*6+1*6+3],image[8*6*6+1*6+4],image[8*6*6+1*6+5],image[8*6*6+2*6+1],image[8*6*6+2*6+2],image[8*6*6+2*6+3],image[8*6*6+2*6+4],image[8*6*6+2*6+5],image[8*6*6+3*6+1],image[8*6*6+3*6+2],image[8*6*6+3*6+3],image[8*6*6+3*6+4],image[8*6*6+3*6+5],image[8*6*6+4*6+1],image[8*6*6+4*6+2],image[8*6*6+4*6+3],image[8*6*6+4*6+4],image[8*6*6+4*6+5],image[9*6*6+0*6+1],image[9*6*6+0*6+2],image[9*6*6+0*6+3],image[9*6*6+0*6+4],image[9*6*6+0*6+5],image[9*6*6+1*6+1],image[9*6*6+1*6+2],image[9*6*6+1*6+3],image[9*6*6+1*6+4],image[9*6*6+1*6+5],image[9*6*6+2*6+1],image[9*6*6+2*6+2],image[9*6*6+2*6+3],image[9*6*6+2*6+4],image[9*6*6+2*6+5],image[9*6*6+3*6+1],image[9*6*6+3*6+2],image[9*6*6+3*6+3],image[9*6*6+3*6+4],image[9*6*6+3*6+5],image[9*6*6+4*6+1],image[9*6*6+4*6+2],image[9*6*6+4*6+3],image[9*6*6+4*6+4],image[9*6*6+4*6+5],image[10*6*6+0*6+1],image[10*6*6+0*6+2],image[10*6*6+0*6+3],image[10*6*6+0*6+4],image[10*6*6+0*6+5],image[10*6*6+1*6+1],image[10*6*6+1*6+2],image[10*6*6+1*6+3],image[10*6*6+1*6+4],image[10*6*6+1*6+5],image[10*6*6+2*6+1],image[10*6*6+2*6+2],image[10*6*6+2*6+3],image[10*6*6+2*6+4],image[10*6*6+2*6+5],image[10*6*6+3*6+1],image[10*6*6+3*6+2],image[10*6*6+3*6+3],image[10*6*6+3*6+4],image[10*6*6+3*6+5],image[10*6*6+4*6+1],image[10*6*6+4*6+2],image[10*6*6+4*6+3],image[10*6*6+4*6+4],image[10*6*6+4*6+5],image[11*6*6+0*6+1],image[11*6*6+0*6+2],image[11*6*6+0*6+3],image[11*6*6+0*6+4],image[11*6*6+0*6+5],image[11*6*6+1*6+1],image[11*6*6+1*6+2],image[11*6*6+1*6+3],image[11*6*6+1*6+4],image[11*6*6+1*6+5],image[11*6*6+2*6+1],image[11*6*6+2*6+2],image[11*6*6+2*6+3],image[11*6*6+2*6+4],image[11*6*6+2*6+5],image[11*6*6+3*6+1],image[11*6*6+3*6+2],image[11*6*6+3*6+3],image[11*6*6+3*6+4],image[11*6*6+3*6+5],image[11*6*6+4*6+1],image[11*6*6+4*6+2],image[11*6*6+4*6+3],image[11*6*6+4*6+4],image[11*6*6+4*6+5],image[12*6*6+0*6+1],image[12*6*6+0*6+2],image[12*6*6+0*6+3],image[12*6*6+0*6+4],image[12*6*6+0*6+5],image[12*6*6+1*6+1],image[12*6*6+1*6+2],image[12*6*6+1*6+3],image[12*6*6+1*6+4],image[12*6*6+1*6+5],image[12*6*6+2*6+1],image[12*6*6+2*6+2],image[12*6*6+2*6+3],image[12*6*6+2*6+4],image[12*6*6+2*6+5],image[12*6*6+3*6+1],image[12*6*6+3*6+2],image[12*6*6+3*6+3],image[12*6*6+3*6+4],image[12*6*6+3*6+5],image[12*6*6+4*6+1],image[12*6*6+4*6+2],image[12*6*6+4*6+3],image[12*6*6+4*6+4],image[12*6*6+4*6+5],image[13*6*6+0*6+1],image[13*6*6+0*6+2],image[13*6*6+0*6+3],image[13*6*6+0*6+4],image[13*6*6+0*6+5],image[13*6*6+1*6+1],image[13*6*6+1*6+2],image[13*6*6+1*6+3],image[13*6*6+1*6+4],image[13*6*6+1*6+5],image[13*6*6+2*6+1],image[13*6*6+2*6+2],image[13*6*6+2*6+3],image[13*6*6+2*6+4],image[13*6*6+2*6+5],image[13*6*6+3*6+1],image[13*6*6+3*6+2],image[13*6*6+3*6+3],image[13*6*6+3*6+4],image[13*6*6+3*6+5],image[13*6*6+4*6+1],image[13*6*6+4*6+2],image[13*6*6+4*6+3],image[13*6*6+4*6+4],image[13*6*6+4*6+5],image[14*6*6+0*6+1],image[14*6*6+0*6+2],image[14*6*6+0*6+3],image[14*6*6+0*6+4],image[14*6*6+0*6+5],image[14*6*6+1*6+1],image[14*6*6+1*6+2],image[14*6*6+1*6+3],image[14*6*6+1*6+4],image[14*6*6+1*6+5],image[14*6*6+2*6+1],image[14*6*6+2*6+2],image[14*6*6+2*6+3],image[14*6*6+2*6+4],image[14*6*6+2*6+5],image[14*6*6+3*6+1],image[14*6*6+3*6+2],image[14*6*6+3*6+3],image[14*6*6+3*6+4],image[14*6*6+3*6+5],image[14*6*6+4*6+1],image[14*6*6+4*6+2],image[14*6*6+4*6+3],image[14*6*6+4*6+4],image[14*6*6+4*6+5],image[15*6*6+0*6+1],image[15*6*6+0*6+2],image[15*6*6+0*6+3],image[15*6*6+0*6+4],image[15*6*6+0*6+5],image[15*6*6+1*6+1],image[15*6*6+1*6+2],image[15*6*6+1*6+3],image[15*6*6+1*6+4],image[15*6*6+1*6+5],image[15*6*6+2*6+1],image[15*6*6+2*6+2],image[15*6*6+2*6+3],image[15*6*6+2*6+4],image[15*6*6+2*6+5],image[15*6*6+3*6+1],image[15*6*6+3*6+2],image[15*6*6+3*6+3],image[15*6*6+3*6+4],image[15*6*6+3*6+5],image[15*6*6+4*6+1],image[15*6*6+4*6+2],image[15*6*6+4*6+3],image[15*6*6+4*6+4],image[15*6*6+4*6+5],image[16*6*6+0*6+1],image[16*6*6+0*6+2],image[16*6*6+0*6+3],image[16*6*6+0*6+4],image[16*6*6+0*6+5],image[16*6*6+1*6+1],image[16*6*6+1*6+2],image[16*6*6+1*6+3],image[16*6*6+1*6+4],image[16*6*6+1*6+5],image[16*6*6+2*6+1],image[16*6*6+2*6+2],image[16*6*6+2*6+3],image[16*6*6+2*6+4],image[16*6*6+2*6+5],image[16*6*6+3*6+1],image[16*6*6+3*6+2],image[16*6*6+3*6+3],image[16*6*6+3*6+4],image[16*6*6+3*6+5],image[16*6*6+4*6+1],image[16*6*6+4*6+2],image[16*6*6+4*6+3],image[16*6*6+4*6+4],image[16*6*6+4*6+5],image[17*6*6+0*6+1],image[17*6*6+0*6+2],image[17*6*6+0*6+3],image[17*6*6+0*6+4],image[17*6*6+0*6+5],image[17*6*6+1*6+1],image[17*6*6+1*6+2],image[17*6*6+1*6+3],image[17*6*6+1*6+4],image[17*6*6+1*6+5],image[17*6*6+2*6+1],image[17*6*6+2*6+2],image[17*6*6+2*6+3],image[17*6*6+2*6+4],image[17*6*6+2*6+5],image[17*6*6+3*6+1],image[17*6*6+3*6+2],image[17*6*6+3*6+3],image[17*6*6+3*6+4],image[17*6*6+3*6+5],image[17*6*6+4*6+1],image[17*6*6+4*6+2],image[17*6*6+4*6+3],image[17*6*6+4*6+4],image[17*6*6+4*6+5]};
logic [chan*5*5-1:0] image_slice3;
assign image_slice3 = {image[0*6*6+1*6+0],image[0*6*6+1*6+1],image[0*6*6+1*6+2],image[0*6*6+1*6+3],image[0*6*6+1*6+4],image[0*6*6+2*6+0],image[0*6*6+2*6+1],image[0*6*6+2*6+2],image[0*6*6+2*6+3],image[0*6*6+2*6+4],image[0*6*6+3*6+0],image[0*6*6+3*6+1],image[0*6*6+3*6+2],image[0*6*6+3*6+3],image[0*6*6+3*6+4],image[0*6*6+4*6+0],image[0*6*6+4*6+1],image[0*6*6+4*6+2],image[0*6*6+4*6+3],image[0*6*6+4*6+4],image[0*6*6+5*6+0],image[0*6*6+5*6+1],image[0*6*6+5*6+2],image[0*6*6+5*6+3],image[0*6*6+5*6+4],image[1*6*6+1*6+0],image[1*6*6+1*6+1],image[1*6*6+1*6+2],image[1*6*6+1*6+3],image[1*6*6+1*6+4],image[1*6*6+2*6+0],image[1*6*6+2*6+1],image[1*6*6+2*6+2],image[1*6*6+2*6+3],image[1*6*6+2*6+4],image[1*6*6+3*6+0],image[1*6*6+3*6+1],image[1*6*6+3*6+2],image[1*6*6+3*6+3],image[1*6*6+3*6+4],image[1*6*6+4*6+0],image[1*6*6+4*6+1],image[1*6*6+4*6+2],image[1*6*6+4*6+3],image[1*6*6+4*6+4],image[1*6*6+5*6+0],image[1*6*6+5*6+1],image[1*6*6+5*6+2],image[1*6*6+5*6+3],image[1*6*6+5*6+4],image[2*6*6+1*6+0],image[2*6*6+1*6+1],image[2*6*6+1*6+2],image[2*6*6+1*6+3],image[2*6*6+1*6+4],image[2*6*6+2*6+0],image[2*6*6+2*6+1],image[2*6*6+2*6+2],image[2*6*6+2*6+3],image[2*6*6+2*6+4],image[2*6*6+3*6+0],image[2*6*6+3*6+1],image[2*6*6+3*6+2],image[2*6*6+3*6+3],image[2*6*6+3*6+4],image[2*6*6+4*6+0],image[2*6*6+4*6+1],image[2*6*6+4*6+2],image[2*6*6+4*6+3],image[2*6*6+4*6+4],image[2*6*6+5*6+0],image[2*6*6+5*6+1],image[2*6*6+5*6+2],image[2*6*6+5*6+3],image[2*6*6+5*6+4],image[3*6*6+1*6+0],image[3*6*6+1*6+1],image[3*6*6+1*6+2],image[3*6*6+1*6+3],image[3*6*6+1*6+4],image[3*6*6+2*6+0],image[3*6*6+2*6+1],image[3*6*6+2*6+2],image[3*6*6+2*6+3],image[3*6*6+2*6+4],image[3*6*6+3*6+0],image[3*6*6+3*6+1],image[3*6*6+3*6+2],image[3*6*6+3*6+3],image[3*6*6+3*6+4],image[3*6*6+4*6+0],image[3*6*6+4*6+1],image[3*6*6+4*6+2],image[3*6*6+4*6+3],image[3*6*6+4*6+4],image[3*6*6+5*6+0],image[3*6*6+5*6+1],image[3*6*6+5*6+2],image[3*6*6+5*6+3],image[3*6*6+5*6+4],image[4*6*6+1*6+0],image[4*6*6+1*6+1],image[4*6*6+1*6+2],image[4*6*6+1*6+3],image[4*6*6+1*6+4],image[4*6*6+2*6+0],image[4*6*6+2*6+1],image[4*6*6+2*6+2],image[4*6*6+2*6+3],image[4*6*6+2*6+4],image[4*6*6+3*6+0],image[4*6*6+3*6+1],image[4*6*6+3*6+2],image[4*6*6+3*6+3],image[4*6*6+3*6+4],image[4*6*6+4*6+0],image[4*6*6+4*6+1],image[4*6*6+4*6+2],image[4*6*6+4*6+3],image[4*6*6+4*6+4],image[4*6*6+5*6+0],image[4*6*6+5*6+1],image[4*6*6+5*6+2],image[4*6*6+5*6+3],image[4*6*6+5*6+4],image[5*6*6+1*6+0],image[5*6*6+1*6+1],image[5*6*6+1*6+2],image[5*6*6+1*6+3],image[5*6*6+1*6+4],image[5*6*6+2*6+0],image[5*6*6+2*6+1],image[5*6*6+2*6+2],image[5*6*6+2*6+3],image[5*6*6+2*6+4],image[5*6*6+3*6+0],image[5*6*6+3*6+1],image[5*6*6+3*6+2],image[5*6*6+3*6+3],image[5*6*6+3*6+4],image[5*6*6+4*6+0],image[5*6*6+4*6+1],image[5*6*6+4*6+2],image[5*6*6+4*6+3],image[5*6*6+4*6+4],image[5*6*6+5*6+0],image[5*6*6+5*6+1],image[5*6*6+5*6+2],image[5*6*6+5*6+3],image[5*6*6+5*6+4],image[6*6*6+1*6+0],image[6*6*6+1*6+1],image[6*6*6+1*6+2],image[6*6*6+1*6+3],image[6*6*6+1*6+4],image[6*6*6+2*6+0],image[6*6*6+2*6+1],image[6*6*6+2*6+2],image[6*6*6+2*6+3],image[6*6*6+2*6+4],image[6*6*6+3*6+0],image[6*6*6+3*6+1],image[6*6*6+3*6+2],image[6*6*6+3*6+3],image[6*6*6+3*6+4],image[6*6*6+4*6+0],image[6*6*6+4*6+1],image[6*6*6+4*6+2],image[6*6*6+4*6+3],image[6*6*6+4*6+4],image[6*6*6+5*6+0],image[6*6*6+5*6+1],image[6*6*6+5*6+2],image[6*6*6+5*6+3],image[6*6*6+5*6+4],image[7*6*6+1*6+0],image[7*6*6+1*6+1],image[7*6*6+1*6+2],image[7*6*6+1*6+3],image[7*6*6+1*6+4],image[7*6*6+2*6+0],image[7*6*6+2*6+1],image[7*6*6+2*6+2],image[7*6*6+2*6+3],image[7*6*6+2*6+4],image[7*6*6+3*6+0],image[7*6*6+3*6+1],image[7*6*6+3*6+2],image[7*6*6+3*6+3],image[7*6*6+3*6+4],image[7*6*6+4*6+0],image[7*6*6+4*6+1],image[7*6*6+4*6+2],image[7*6*6+4*6+3],image[7*6*6+4*6+4],image[7*6*6+5*6+0],image[7*6*6+5*6+1],image[7*6*6+5*6+2],image[7*6*6+5*6+3],image[7*6*6+5*6+4],image[8*6*6+1*6+0],image[8*6*6+1*6+1],image[8*6*6+1*6+2],image[8*6*6+1*6+3],image[8*6*6+1*6+4],image[8*6*6+2*6+0],image[8*6*6+2*6+1],image[8*6*6+2*6+2],image[8*6*6+2*6+3],image[8*6*6+2*6+4],image[8*6*6+3*6+0],image[8*6*6+3*6+1],image[8*6*6+3*6+2],image[8*6*6+3*6+3],image[8*6*6+3*6+4],image[8*6*6+4*6+0],image[8*6*6+4*6+1],image[8*6*6+4*6+2],image[8*6*6+4*6+3],image[8*6*6+4*6+4],image[8*6*6+5*6+0],image[8*6*6+5*6+1],image[8*6*6+5*6+2],image[8*6*6+5*6+3],image[8*6*6+5*6+4],image[9*6*6+1*6+0],image[9*6*6+1*6+1],image[9*6*6+1*6+2],image[9*6*6+1*6+3],image[9*6*6+1*6+4],image[9*6*6+2*6+0],image[9*6*6+2*6+1],image[9*6*6+2*6+2],image[9*6*6+2*6+3],image[9*6*6+2*6+4],image[9*6*6+3*6+0],image[9*6*6+3*6+1],image[9*6*6+3*6+2],image[9*6*6+3*6+3],image[9*6*6+3*6+4],image[9*6*6+4*6+0],image[9*6*6+4*6+1],image[9*6*6+4*6+2],image[9*6*6+4*6+3],image[9*6*6+4*6+4],image[9*6*6+5*6+0],image[9*6*6+5*6+1],image[9*6*6+5*6+2],image[9*6*6+5*6+3],image[9*6*6+5*6+4],image[10*6*6+1*6+0],image[10*6*6+1*6+1],image[10*6*6+1*6+2],image[10*6*6+1*6+3],image[10*6*6+1*6+4],image[10*6*6+2*6+0],image[10*6*6+2*6+1],image[10*6*6+2*6+2],image[10*6*6+2*6+3],image[10*6*6+2*6+4],image[10*6*6+3*6+0],image[10*6*6+3*6+1],image[10*6*6+3*6+2],image[10*6*6+3*6+3],image[10*6*6+3*6+4],image[10*6*6+4*6+0],image[10*6*6+4*6+1],image[10*6*6+4*6+2],image[10*6*6+4*6+3],image[10*6*6+4*6+4],image[10*6*6+5*6+0],image[10*6*6+5*6+1],image[10*6*6+5*6+2],image[10*6*6+5*6+3],image[10*6*6+5*6+4],image[11*6*6+1*6+0],image[11*6*6+1*6+1],image[11*6*6+1*6+2],image[11*6*6+1*6+3],image[11*6*6+1*6+4],image[11*6*6+2*6+0],image[11*6*6+2*6+1],image[11*6*6+2*6+2],image[11*6*6+2*6+3],image[11*6*6+2*6+4],image[11*6*6+3*6+0],image[11*6*6+3*6+1],image[11*6*6+3*6+2],image[11*6*6+3*6+3],image[11*6*6+3*6+4],image[11*6*6+4*6+0],image[11*6*6+4*6+1],image[11*6*6+4*6+2],image[11*6*6+4*6+3],image[11*6*6+4*6+4],image[11*6*6+5*6+0],image[11*6*6+5*6+1],image[11*6*6+5*6+2],image[11*6*6+5*6+3],image[11*6*6+5*6+4],image[12*6*6+1*6+0],image[12*6*6+1*6+1],image[12*6*6+1*6+2],image[12*6*6+1*6+3],image[12*6*6+1*6+4],image[12*6*6+2*6+0],image[12*6*6+2*6+1],image[12*6*6+2*6+2],image[12*6*6+2*6+3],image[12*6*6+2*6+4],image[12*6*6+3*6+0],image[12*6*6+3*6+1],image[12*6*6+3*6+2],image[12*6*6+3*6+3],image[12*6*6+3*6+4],image[12*6*6+4*6+0],image[12*6*6+4*6+1],image[12*6*6+4*6+2],image[12*6*6+4*6+3],image[12*6*6+4*6+4],image[12*6*6+5*6+0],image[12*6*6+5*6+1],image[12*6*6+5*6+2],image[12*6*6+5*6+3],image[12*6*6+5*6+4],image[13*6*6+1*6+0],image[13*6*6+1*6+1],image[13*6*6+1*6+2],image[13*6*6+1*6+3],image[13*6*6+1*6+4],image[13*6*6+2*6+0],image[13*6*6+2*6+1],image[13*6*6+2*6+2],image[13*6*6+2*6+3],image[13*6*6+2*6+4],image[13*6*6+3*6+0],image[13*6*6+3*6+1],image[13*6*6+3*6+2],image[13*6*6+3*6+3],image[13*6*6+3*6+4],image[13*6*6+4*6+0],image[13*6*6+4*6+1],image[13*6*6+4*6+2],image[13*6*6+4*6+3],image[13*6*6+4*6+4],image[13*6*6+5*6+0],image[13*6*6+5*6+1],image[13*6*6+5*6+2],image[13*6*6+5*6+3],image[13*6*6+5*6+4],image[14*6*6+1*6+0],image[14*6*6+1*6+1],image[14*6*6+1*6+2],image[14*6*6+1*6+3],image[14*6*6+1*6+4],image[14*6*6+2*6+0],image[14*6*6+2*6+1],image[14*6*6+2*6+2],image[14*6*6+2*6+3],image[14*6*6+2*6+4],image[14*6*6+3*6+0],image[14*6*6+3*6+1],image[14*6*6+3*6+2],image[14*6*6+3*6+3],image[14*6*6+3*6+4],image[14*6*6+4*6+0],image[14*6*6+4*6+1],image[14*6*6+4*6+2],image[14*6*6+4*6+3],image[14*6*6+4*6+4],image[14*6*6+5*6+0],image[14*6*6+5*6+1],image[14*6*6+5*6+2],image[14*6*6+5*6+3],image[14*6*6+5*6+4],image[15*6*6+1*6+0],image[15*6*6+1*6+1],image[15*6*6+1*6+2],image[15*6*6+1*6+3],image[15*6*6+1*6+4],image[15*6*6+2*6+0],image[15*6*6+2*6+1],image[15*6*6+2*6+2],image[15*6*6+2*6+3],image[15*6*6+2*6+4],image[15*6*6+3*6+0],image[15*6*6+3*6+1],image[15*6*6+3*6+2],image[15*6*6+3*6+3],image[15*6*6+3*6+4],image[15*6*6+4*6+0],image[15*6*6+4*6+1],image[15*6*6+4*6+2],image[15*6*6+4*6+3],image[15*6*6+4*6+4],image[15*6*6+5*6+0],image[15*6*6+5*6+1],image[15*6*6+5*6+2],image[15*6*6+5*6+3],image[15*6*6+5*6+4],image[16*6*6+1*6+0],image[16*6*6+1*6+1],image[16*6*6+1*6+2],image[16*6*6+1*6+3],image[16*6*6+1*6+4],image[16*6*6+2*6+0],image[16*6*6+2*6+1],image[16*6*6+2*6+2],image[16*6*6+2*6+3],image[16*6*6+2*6+4],image[16*6*6+3*6+0],image[16*6*6+3*6+1],image[16*6*6+3*6+2],image[16*6*6+3*6+3],image[16*6*6+3*6+4],image[16*6*6+4*6+0],image[16*6*6+4*6+1],image[16*6*6+4*6+2],image[16*6*6+4*6+3],image[16*6*6+4*6+4],image[16*6*6+5*6+0],image[16*6*6+5*6+1],image[16*6*6+5*6+2],image[16*6*6+5*6+3],image[16*6*6+5*6+4],image[17*6*6+1*6+0],image[17*6*6+1*6+1],image[17*6*6+1*6+2],image[17*6*6+1*6+3],image[17*6*6+1*6+4],image[17*6*6+2*6+0],image[17*6*6+2*6+1],image[17*6*6+2*6+2],image[17*6*6+2*6+3],image[17*6*6+2*6+4],image[17*6*6+3*6+0],image[17*6*6+3*6+1],image[17*6*6+3*6+2],image[17*6*6+3*6+3],image[17*6*6+3*6+4],image[17*6*6+4*6+0],image[17*6*6+4*6+1],image[17*6*6+4*6+2],image[17*6*6+4*6+3],image[17*6*6+4*6+4],image[17*6*6+5*6+0],image[17*6*6+5*6+1],image[17*6*6+5*6+2],image[17*6*6+5*6+3],image[17*6*6+5*6+4]};
logic [chan*5*5-1:0] image_slice4;
assign image_slice4 = {image[0*6*6+1*6+1],image[0*6*6+1*6+2],image[0*6*6+1*6+3],image[0*6*6+1*6+4],image[0*6*6+1*6+5],image[0*6*6+2*6+1],image[0*6*6+2*6+2],image[0*6*6+2*6+3],image[0*6*6+2*6+4],image[0*6*6+2*6+5],image[0*6*6+3*6+1],image[0*6*6+3*6+2],image[0*6*6+3*6+3],image[0*6*6+3*6+4],image[0*6*6+3*6+5],image[0*6*6+4*6+1],image[0*6*6+4*6+2],image[0*6*6+4*6+3],image[0*6*6+4*6+4],image[0*6*6+4*6+5],image[0*6*6+5*6+1],image[0*6*6+5*6+2],image[0*6*6+5*6+3],image[0*6*6+5*6+4],image[0*6*6+5*6+5],image[1*6*6+1*6+1],image[1*6*6+1*6+2],image[1*6*6+1*6+3],image[1*6*6+1*6+4],image[1*6*6+1*6+5],image[1*6*6+2*6+1],image[1*6*6+2*6+2],image[1*6*6+2*6+3],image[1*6*6+2*6+4],image[1*6*6+2*6+5],image[1*6*6+3*6+1],image[1*6*6+3*6+2],image[1*6*6+3*6+3],image[1*6*6+3*6+4],image[1*6*6+3*6+5],image[1*6*6+4*6+1],image[1*6*6+4*6+2],image[1*6*6+4*6+3],image[1*6*6+4*6+4],image[1*6*6+4*6+5],image[1*6*6+5*6+1],image[1*6*6+5*6+2],image[1*6*6+5*6+3],image[1*6*6+5*6+4],image[1*6*6+5*6+5],image[2*6*6+1*6+1],image[2*6*6+1*6+2],image[2*6*6+1*6+3],image[2*6*6+1*6+4],image[2*6*6+1*6+5],image[2*6*6+2*6+1],image[2*6*6+2*6+2],image[2*6*6+2*6+3],image[2*6*6+2*6+4],image[2*6*6+2*6+5],image[2*6*6+3*6+1],image[2*6*6+3*6+2],image[2*6*6+3*6+3],image[2*6*6+3*6+4],image[2*6*6+3*6+5],image[2*6*6+4*6+1],image[2*6*6+4*6+2],image[2*6*6+4*6+3],image[2*6*6+4*6+4],image[2*6*6+4*6+5],image[2*6*6+5*6+1],image[2*6*6+5*6+2],image[2*6*6+5*6+3],image[2*6*6+5*6+4],image[2*6*6+5*6+5],image[3*6*6+1*6+1],image[3*6*6+1*6+2],image[3*6*6+1*6+3],image[3*6*6+1*6+4],image[3*6*6+1*6+5],image[3*6*6+2*6+1],image[3*6*6+2*6+2],image[3*6*6+2*6+3],image[3*6*6+2*6+4],image[3*6*6+2*6+5],image[3*6*6+3*6+1],image[3*6*6+3*6+2],image[3*6*6+3*6+3],image[3*6*6+3*6+4],image[3*6*6+3*6+5],image[3*6*6+4*6+1],image[3*6*6+4*6+2],image[3*6*6+4*6+3],image[3*6*6+4*6+4],image[3*6*6+4*6+5],image[3*6*6+5*6+1],image[3*6*6+5*6+2],image[3*6*6+5*6+3],image[3*6*6+5*6+4],image[3*6*6+5*6+5],image[4*6*6+1*6+1],image[4*6*6+1*6+2],image[4*6*6+1*6+3],image[4*6*6+1*6+4],image[4*6*6+1*6+5],image[4*6*6+2*6+1],image[4*6*6+2*6+2],image[4*6*6+2*6+3],image[4*6*6+2*6+4],image[4*6*6+2*6+5],image[4*6*6+3*6+1],image[4*6*6+3*6+2],image[4*6*6+3*6+3],image[4*6*6+3*6+4],image[4*6*6+3*6+5],image[4*6*6+4*6+1],image[4*6*6+4*6+2],image[4*6*6+4*6+3],image[4*6*6+4*6+4],image[4*6*6+4*6+5],image[4*6*6+5*6+1],image[4*6*6+5*6+2],image[4*6*6+5*6+3],image[4*6*6+5*6+4],image[4*6*6+5*6+5],image[5*6*6+1*6+1],image[5*6*6+1*6+2],image[5*6*6+1*6+3],image[5*6*6+1*6+4],image[5*6*6+1*6+5],image[5*6*6+2*6+1],image[5*6*6+2*6+2],image[5*6*6+2*6+3],image[5*6*6+2*6+4],image[5*6*6+2*6+5],image[5*6*6+3*6+1],image[5*6*6+3*6+2],image[5*6*6+3*6+3],image[5*6*6+3*6+4],image[5*6*6+3*6+5],image[5*6*6+4*6+1],image[5*6*6+4*6+2],image[5*6*6+4*6+3],image[5*6*6+4*6+4],image[5*6*6+4*6+5],image[5*6*6+5*6+1],image[5*6*6+5*6+2],image[5*6*6+5*6+3],image[5*6*6+5*6+4],image[5*6*6+5*6+5],image[6*6*6+1*6+1],image[6*6*6+1*6+2],image[6*6*6+1*6+3],image[6*6*6+1*6+4],image[6*6*6+1*6+5],image[6*6*6+2*6+1],image[6*6*6+2*6+2],image[6*6*6+2*6+3],image[6*6*6+2*6+4],image[6*6*6+2*6+5],image[6*6*6+3*6+1],image[6*6*6+3*6+2],image[6*6*6+3*6+3],image[6*6*6+3*6+4],image[6*6*6+3*6+5],image[6*6*6+4*6+1],image[6*6*6+4*6+2],image[6*6*6+4*6+3],image[6*6*6+4*6+4],image[6*6*6+4*6+5],image[6*6*6+5*6+1],image[6*6*6+5*6+2],image[6*6*6+5*6+3],image[6*6*6+5*6+4],image[6*6*6+5*6+5],image[7*6*6+1*6+1],image[7*6*6+1*6+2],image[7*6*6+1*6+3],image[7*6*6+1*6+4],image[7*6*6+1*6+5],image[7*6*6+2*6+1],image[7*6*6+2*6+2],image[7*6*6+2*6+3],image[7*6*6+2*6+4],image[7*6*6+2*6+5],image[7*6*6+3*6+1],image[7*6*6+3*6+2],image[7*6*6+3*6+3],image[7*6*6+3*6+4],image[7*6*6+3*6+5],image[7*6*6+4*6+1],image[7*6*6+4*6+2],image[7*6*6+4*6+3],image[7*6*6+4*6+4],image[7*6*6+4*6+5],image[7*6*6+5*6+1],image[7*6*6+5*6+2],image[7*6*6+5*6+3],image[7*6*6+5*6+4],image[7*6*6+5*6+5],image[8*6*6+1*6+1],image[8*6*6+1*6+2],image[8*6*6+1*6+3],image[8*6*6+1*6+4],image[8*6*6+1*6+5],image[8*6*6+2*6+1],image[8*6*6+2*6+2],image[8*6*6+2*6+3],image[8*6*6+2*6+4],image[8*6*6+2*6+5],image[8*6*6+3*6+1],image[8*6*6+3*6+2],image[8*6*6+3*6+3],image[8*6*6+3*6+4],image[8*6*6+3*6+5],image[8*6*6+4*6+1],image[8*6*6+4*6+2],image[8*6*6+4*6+3],image[8*6*6+4*6+4],image[8*6*6+4*6+5],image[8*6*6+5*6+1],image[8*6*6+5*6+2],image[8*6*6+5*6+3],image[8*6*6+5*6+4],image[8*6*6+5*6+5],image[9*6*6+1*6+1],image[9*6*6+1*6+2],image[9*6*6+1*6+3],image[9*6*6+1*6+4],image[9*6*6+1*6+5],image[9*6*6+2*6+1],image[9*6*6+2*6+2],image[9*6*6+2*6+3],image[9*6*6+2*6+4],image[9*6*6+2*6+5],image[9*6*6+3*6+1],image[9*6*6+3*6+2],image[9*6*6+3*6+3],image[9*6*6+3*6+4],image[9*6*6+3*6+5],image[9*6*6+4*6+1],image[9*6*6+4*6+2],image[9*6*6+4*6+3],image[9*6*6+4*6+4],image[9*6*6+4*6+5],image[9*6*6+5*6+1],image[9*6*6+5*6+2],image[9*6*6+5*6+3],image[9*6*6+5*6+4],image[9*6*6+5*6+5],image[10*6*6+1*6+1],image[10*6*6+1*6+2],image[10*6*6+1*6+3],image[10*6*6+1*6+4],image[10*6*6+1*6+5],image[10*6*6+2*6+1],image[10*6*6+2*6+2],image[10*6*6+2*6+3],image[10*6*6+2*6+4],image[10*6*6+2*6+5],image[10*6*6+3*6+1],image[10*6*6+3*6+2],image[10*6*6+3*6+3],image[10*6*6+3*6+4],image[10*6*6+3*6+5],image[10*6*6+4*6+1],image[10*6*6+4*6+2],image[10*6*6+4*6+3],image[10*6*6+4*6+4],image[10*6*6+4*6+5],image[10*6*6+5*6+1],image[10*6*6+5*6+2],image[10*6*6+5*6+3],image[10*6*6+5*6+4],image[10*6*6+5*6+5],image[11*6*6+1*6+1],image[11*6*6+1*6+2],image[11*6*6+1*6+3],image[11*6*6+1*6+4],image[11*6*6+1*6+5],image[11*6*6+2*6+1],image[11*6*6+2*6+2],image[11*6*6+2*6+3],image[11*6*6+2*6+4],image[11*6*6+2*6+5],image[11*6*6+3*6+1],image[11*6*6+3*6+2],image[11*6*6+3*6+3],image[11*6*6+3*6+4],image[11*6*6+3*6+5],image[11*6*6+4*6+1],image[11*6*6+4*6+2],image[11*6*6+4*6+3],image[11*6*6+4*6+4],image[11*6*6+4*6+5],image[11*6*6+5*6+1],image[11*6*6+5*6+2],image[11*6*6+5*6+3],image[11*6*6+5*6+4],image[11*6*6+5*6+5],image[12*6*6+1*6+1],image[12*6*6+1*6+2],image[12*6*6+1*6+3],image[12*6*6+1*6+4],image[12*6*6+1*6+5],image[12*6*6+2*6+1],image[12*6*6+2*6+2],image[12*6*6+2*6+3],image[12*6*6+2*6+4],image[12*6*6+2*6+5],image[12*6*6+3*6+1],image[12*6*6+3*6+2],image[12*6*6+3*6+3],image[12*6*6+3*6+4],image[12*6*6+3*6+5],image[12*6*6+4*6+1],image[12*6*6+4*6+2],image[12*6*6+4*6+3],image[12*6*6+4*6+4],image[12*6*6+4*6+5],image[12*6*6+5*6+1],image[12*6*6+5*6+2],image[12*6*6+5*6+3],image[12*6*6+5*6+4],image[12*6*6+5*6+5],image[13*6*6+1*6+1],image[13*6*6+1*6+2],image[13*6*6+1*6+3],image[13*6*6+1*6+4],image[13*6*6+1*6+5],image[13*6*6+2*6+1],image[13*6*6+2*6+2],image[13*6*6+2*6+3],image[13*6*6+2*6+4],image[13*6*6+2*6+5],image[13*6*6+3*6+1],image[13*6*6+3*6+2],image[13*6*6+3*6+3],image[13*6*6+3*6+4],image[13*6*6+3*6+5],image[13*6*6+4*6+1],image[13*6*6+4*6+2],image[13*6*6+4*6+3],image[13*6*6+4*6+4],image[13*6*6+4*6+5],image[13*6*6+5*6+1],image[13*6*6+5*6+2],image[13*6*6+5*6+3],image[13*6*6+5*6+4],image[13*6*6+5*6+5],image[14*6*6+1*6+1],image[14*6*6+1*6+2],image[14*6*6+1*6+3],image[14*6*6+1*6+4],image[14*6*6+1*6+5],image[14*6*6+2*6+1],image[14*6*6+2*6+2],image[14*6*6+2*6+3],image[14*6*6+2*6+4],image[14*6*6+2*6+5],image[14*6*6+3*6+1],image[14*6*6+3*6+2],image[14*6*6+3*6+3],image[14*6*6+3*6+4],image[14*6*6+3*6+5],image[14*6*6+4*6+1],image[14*6*6+4*6+2],image[14*6*6+4*6+3],image[14*6*6+4*6+4],image[14*6*6+4*6+5],image[14*6*6+5*6+1],image[14*6*6+5*6+2],image[14*6*6+5*6+3],image[14*6*6+5*6+4],image[14*6*6+5*6+5],image[15*6*6+1*6+1],image[15*6*6+1*6+2],image[15*6*6+1*6+3],image[15*6*6+1*6+4],image[15*6*6+1*6+5],image[15*6*6+2*6+1],image[15*6*6+2*6+2],image[15*6*6+2*6+3],image[15*6*6+2*6+4],image[15*6*6+2*6+5],image[15*6*6+3*6+1],image[15*6*6+3*6+2],image[15*6*6+3*6+3],image[15*6*6+3*6+4],image[15*6*6+3*6+5],image[15*6*6+4*6+1],image[15*6*6+4*6+2],image[15*6*6+4*6+3],image[15*6*6+4*6+4],image[15*6*6+4*6+5],image[15*6*6+5*6+1],image[15*6*6+5*6+2],image[15*6*6+5*6+3],image[15*6*6+5*6+4],image[15*6*6+5*6+5],image[16*6*6+1*6+1],image[16*6*6+1*6+2],image[16*6*6+1*6+3],image[16*6*6+1*6+4],image[16*6*6+1*6+5],image[16*6*6+2*6+1],image[16*6*6+2*6+2],image[16*6*6+2*6+3],image[16*6*6+2*6+4],image[16*6*6+2*6+5],image[16*6*6+3*6+1],image[16*6*6+3*6+2],image[16*6*6+3*6+3],image[16*6*6+3*6+4],image[16*6*6+3*6+5],image[16*6*6+4*6+1],image[16*6*6+4*6+2],image[16*6*6+4*6+3],image[16*6*6+4*6+4],image[16*6*6+4*6+5],image[16*6*6+5*6+1],image[16*6*6+5*6+2],image[16*6*6+5*6+3],image[16*6*6+5*6+4],image[16*6*6+5*6+5],image[17*6*6+1*6+1],image[17*6*6+1*6+2],image[17*6*6+1*6+3],image[17*6*6+1*6+4],image[17*6*6+1*6+5],image[17*6*6+2*6+1],image[17*6*6+2*6+2],image[17*6*6+2*6+3],image[17*6*6+2*6+4],image[17*6*6+2*6+5],image[17*6*6+3*6+1],image[17*6*6+3*6+2],image[17*6*6+3*6+3],image[17*6*6+3*6+4],image[17*6*6+3*6+5],image[17*6*6+4*6+1],image[17*6*6+4*6+2],image[17*6*6+4*6+3],image[17*6*6+4*6+4],image[17*6*6+4*6+5],image[17*6*6+5*6+1],image[17*6*6+5*6+2],image[17*6*6+5*6+3],image[17*6*6+5*6+4],image[17*6*6+5*6+5]};


logic [0:chan*5*5-1] kernel_slice;
assign kernel_slice = {kernels[0*25+0*5+0],kernels[0*25+0*5+1],kernels[0*25+0*5+2],kernels[0*25+0*5+3],kernels[0*25+0*5+4],kernels[0*25+1*5+0],kernels[0*25+1*5+1],kernels[0*25+1*5+2],kernels[0*25+1*5+3],kernels[0*25+1*5+4],kernels[0*25+2*5+0],kernels[0*25+2*5+1],kernels[0*25+2*5+2],kernels[0*25+2*5+3],kernels[0*25+2*5+4],kernels[0*25+3*5+0],kernels[0*25+3*5+1],kernels[0*25+3*5+2],kernels[0*25+3*5+3],kernels[0*25+3*5+4],kernels[0*25+4*5+0],kernels[0*25+4*5+1],kernels[0*25+4*5+2],kernels[0*25+4*5+3],kernels[0*25+4*5+4],kernels[1*25+0*5+0],kernels[1*25+0*5+1],kernels[1*25+0*5+2],kernels[1*25+0*5+3],kernels[1*25+0*5+4],kernels[1*25+1*5+0],kernels[1*25+1*5+1],kernels[1*25+1*5+2],kernels[1*25+1*5+3],kernels[1*25+1*5+4],kernels[1*25+2*5+0],kernels[1*25+2*5+1],kernels[1*25+2*5+2],kernels[1*25+2*5+3],kernels[1*25+2*5+4],kernels[1*25+3*5+0],kernels[1*25+3*5+1],kernels[1*25+3*5+2],kernels[1*25+3*5+3],kernels[1*25+3*5+4],kernels[1*25+4*5+0],kernels[1*25+4*5+1],kernels[1*25+4*5+2],kernels[1*25+4*5+3],kernels[1*25+4*5+4],kernels[2*25+0*5+0],kernels[2*25+0*5+1],kernels[2*25+0*5+2],kernels[2*25+0*5+3],kernels[2*25+0*5+4],kernels[2*25+1*5+0],kernels[2*25+1*5+1],kernels[2*25+1*5+2],kernels[2*25+1*5+3],kernels[2*25+1*5+4],kernels[2*25+2*5+0],kernels[2*25+2*5+1],kernels[2*25+2*5+2],kernels[2*25+2*5+3],kernels[2*25+2*5+4],kernels[2*25+3*5+0],kernels[2*25+3*5+1],kernels[2*25+3*5+2],kernels[2*25+3*5+3],kernels[2*25+3*5+4],kernels[2*25+4*5+0],kernels[2*25+4*5+1],kernels[2*25+4*5+2],kernels[2*25+4*5+3],kernels[2*25+4*5+4],kernels[3*25+0*5+0],kernels[3*25+0*5+1],kernels[3*25+0*5+2],kernels[3*25+0*5+3],kernels[3*25+0*5+4],kernels[3*25+1*5+0],kernels[3*25+1*5+1],kernels[3*25+1*5+2],kernels[3*25+1*5+3],kernels[3*25+1*5+4],kernels[3*25+2*5+0],kernels[3*25+2*5+1],kernels[3*25+2*5+2],kernels[3*25+2*5+3],kernels[3*25+2*5+4],kernels[3*25+3*5+0],kernels[3*25+3*5+1],kernels[3*25+3*5+2],kernels[3*25+3*5+3],kernels[3*25+3*5+4],kernels[3*25+4*5+0],kernels[3*25+4*5+1],kernels[3*25+4*5+2],kernels[3*25+4*5+3],kernels[3*25+4*5+4],kernels[4*25+0*5+0],kernels[4*25+0*5+1],kernels[4*25+0*5+2],kernels[4*25+0*5+3],kernels[4*25+0*5+4],kernels[4*25+1*5+0],kernels[4*25+1*5+1],kernels[4*25+1*5+2],kernels[4*25+1*5+3],kernels[4*25+1*5+4],kernels[4*25+2*5+0],kernels[4*25+2*5+1],kernels[4*25+2*5+2],kernels[4*25+2*5+3],kernels[4*25+2*5+4],kernels[4*25+3*5+0],kernels[4*25+3*5+1],kernels[4*25+3*5+2],kernels[4*25+3*5+3],kernels[4*25+3*5+4],kernels[4*25+4*5+0],kernels[4*25+4*5+1],kernels[4*25+4*5+2],kernels[4*25+4*5+3],kernels[4*25+4*5+4],kernels[5*25+0*5+0],kernels[5*25+0*5+1],kernels[5*25+0*5+2],kernels[5*25+0*5+3],kernels[5*25+0*5+4],kernels[5*25+1*5+0],kernels[5*25+1*5+1],kernels[5*25+1*5+2],kernels[5*25+1*5+3],kernels[5*25+1*5+4],kernels[5*25+2*5+0],kernels[5*25+2*5+1],kernels[5*25+2*5+2],kernels[5*25+2*5+3],kernels[5*25+2*5+4],kernels[5*25+3*5+0],kernels[5*25+3*5+1],kernels[5*25+3*5+2],kernels[5*25+3*5+3],kernels[5*25+3*5+4],kernels[5*25+4*5+0],kernels[5*25+4*5+1],kernels[5*25+4*5+2],kernels[5*25+4*5+3],kernels[5*25+4*5+4],kernels[6*25+0*5+0],kernels[6*25+0*5+1],kernels[6*25+0*5+2],kernels[6*25+0*5+3],kernels[6*25+0*5+4],kernels[6*25+1*5+0],kernels[6*25+1*5+1],kernels[6*25+1*5+2],kernels[6*25+1*5+3],kernels[6*25+1*5+4],kernels[6*25+2*5+0],kernels[6*25+2*5+1],kernels[6*25+2*5+2],kernels[6*25+2*5+3],kernels[6*25+2*5+4],kernels[6*25+3*5+0],kernels[6*25+3*5+1],kernels[6*25+3*5+2],kernels[6*25+3*5+3],kernels[6*25+3*5+4],kernels[6*25+4*5+0],kernels[6*25+4*5+1],kernels[6*25+4*5+2],kernels[6*25+4*5+3],kernels[6*25+4*5+4],kernels[7*25+0*5+0],kernels[7*25+0*5+1],kernels[7*25+0*5+2],kernels[7*25+0*5+3],kernels[7*25+0*5+4],kernels[7*25+1*5+0],kernels[7*25+1*5+1],kernels[7*25+1*5+2],kernels[7*25+1*5+3],kernels[7*25+1*5+4],kernels[7*25+2*5+0],kernels[7*25+2*5+1],kernels[7*25+2*5+2],kernels[7*25+2*5+3],kernels[7*25+2*5+4],kernels[7*25+3*5+0],kernels[7*25+3*5+1],kernels[7*25+3*5+2],kernels[7*25+3*5+3],kernels[7*25+3*5+4],kernels[7*25+4*5+0],kernels[7*25+4*5+1],kernels[7*25+4*5+2],kernels[7*25+4*5+3],kernels[7*25+4*5+4],kernels[8*25+0*5+0],kernels[8*25+0*5+1],kernels[8*25+0*5+2],kernels[8*25+0*5+3],kernels[8*25+0*5+4],kernels[8*25+1*5+0],kernels[8*25+1*5+1],kernels[8*25+1*5+2],kernels[8*25+1*5+3],kernels[8*25+1*5+4],kernels[8*25+2*5+0],kernels[8*25+2*5+1],kernels[8*25+2*5+2],kernels[8*25+2*5+3],kernels[8*25+2*5+4],kernels[8*25+3*5+0],kernels[8*25+3*5+1],kernels[8*25+3*5+2],kernels[8*25+3*5+3],kernels[8*25+3*5+4],kernels[8*25+4*5+0],kernels[8*25+4*5+1],kernels[8*25+4*5+2],kernels[8*25+4*5+3],kernels[8*25+4*5+4],kernels[9*25+0*5+0],kernels[9*25+0*5+1],kernels[9*25+0*5+2],kernels[9*25+0*5+3],kernels[9*25+0*5+4],kernels[9*25+1*5+0],kernels[9*25+1*5+1],kernels[9*25+1*5+2],kernels[9*25+1*5+3],kernels[9*25+1*5+4],kernels[9*25+2*5+0],kernels[9*25+2*5+1],kernels[9*25+2*5+2],kernels[9*25+2*5+3],kernels[9*25+2*5+4],kernels[9*25+3*5+0],kernels[9*25+3*5+1],kernels[9*25+3*5+2],kernels[9*25+3*5+3],kernels[9*25+3*5+4],kernels[9*25+4*5+0],kernels[9*25+4*5+1],kernels[9*25+4*5+2],kernels[9*25+4*5+3],kernels[9*25+4*5+4],kernels[10*25+0*5+0],kernels[10*25+0*5+1],kernels[10*25+0*5+2],kernels[10*25+0*5+3],kernels[10*25+0*5+4],kernels[10*25+1*5+0],kernels[10*25+1*5+1],kernels[10*25+1*5+2],kernels[10*25+1*5+3],kernels[10*25+1*5+4],kernels[10*25+2*5+0],kernels[10*25+2*5+1],kernels[10*25+2*5+2],kernels[10*25+2*5+3],kernels[10*25+2*5+4],kernels[10*25+3*5+0],kernels[10*25+3*5+1],kernels[10*25+3*5+2],kernels[10*25+3*5+3],kernels[10*25+3*5+4],kernels[10*25+4*5+0],kernels[10*25+4*5+1],kernels[10*25+4*5+2],kernels[10*25+4*5+3],kernels[10*25+4*5+4],kernels[11*25+0*5+0],kernels[11*25+0*5+1],kernels[11*25+0*5+2],kernels[11*25+0*5+3],kernels[11*25+0*5+4],kernels[11*25+1*5+0],kernels[11*25+1*5+1],kernels[11*25+1*5+2],kernels[11*25+1*5+3],kernels[11*25+1*5+4],kernels[11*25+2*5+0],kernels[11*25+2*5+1],kernels[11*25+2*5+2],kernels[11*25+2*5+3],kernels[11*25+2*5+4],kernels[11*25+3*5+0],kernels[11*25+3*5+1],kernels[11*25+3*5+2],kernels[11*25+3*5+3],kernels[11*25+3*5+4],kernels[11*25+4*5+0],kernels[11*25+4*5+1],kernels[11*25+4*5+2],kernels[11*25+4*5+3],kernels[11*25+4*5+4],kernels[12*25+0*5+0],kernels[12*25+0*5+1],kernels[12*25+0*5+2],kernels[12*25+0*5+3],kernels[12*25+0*5+4],kernels[12*25+1*5+0],kernels[12*25+1*5+1],kernels[12*25+1*5+2],kernels[12*25+1*5+3],kernels[12*25+1*5+4],kernels[12*25+2*5+0],kernels[12*25+2*5+1],kernels[12*25+2*5+2],kernels[12*25+2*5+3],kernels[12*25+2*5+4],kernels[12*25+3*5+0],kernels[12*25+3*5+1],kernels[12*25+3*5+2],kernels[12*25+3*5+3],kernels[12*25+3*5+4],kernels[12*25+4*5+0],kernels[12*25+4*5+1],kernels[12*25+4*5+2],kernels[12*25+4*5+3],kernels[12*25+4*5+4],kernels[13*25+0*5+0],kernels[13*25+0*5+1],kernels[13*25+0*5+2],kernels[13*25+0*5+3],kernels[13*25+0*5+4],kernels[13*25+1*5+0],kernels[13*25+1*5+1],kernels[13*25+1*5+2],kernels[13*25+1*5+3],kernels[13*25+1*5+4],kernels[13*25+2*5+0],kernels[13*25+2*5+1],kernels[13*25+2*5+2],kernels[13*25+2*5+3],kernels[13*25+2*5+4],kernels[13*25+3*5+0],kernels[13*25+3*5+1],kernels[13*25+3*5+2],kernels[13*25+3*5+3],kernels[13*25+3*5+4],kernels[13*25+4*5+0],kernels[13*25+4*5+1],kernels[13*25+4*5+2],kernels[13*25+4*5+3],kernels[13*25+4*5+4],kernels[14*25+0*5+0],kernels[14*25+0*5+1],kernels[14*25+0*5+2],kernels[14*25+0*5+3],kernels[14*25+0*5+4],kernels[14*25+1*5+0],kernels[14*25+1*5+1],kernels[14*25+1*5+2],kernels[14*25+1*5+3],kernels[14*25+1*5+4],kernels[14*25+2*5+0],kernels[14*25+2*5+1],kernels[14*25+2*5+2],kernels[14*25+2*5+3],kernels[14*25+2*5+4],kernels[14*25+3*5+0],kernels[14*25+3*5+1],kernels[14*25+3*5+2],kernels[14*25+3*5+3],kernels[14*25+3*5+4],kernels[14*25+4*5+0],kernels[14*25+4*5+1],kernels[14*25+4*5+2],kernels[14*25+4*5+3],kernels[14*25+4*5+4],kernels[15*25+0*5+0],kernels[15*25+0*5+1],kernels[15*25+0*5+2],kernels[15*25+0*5+3],kernels[15*25+0*5+4],kernels[15*25+1*5+0],kernels[15*25+1*5+1],kernels[15*25+1*5+2],kernels[15*25+1*5+3],kernels[15*25+1*5+4],kernels[15*25+2*5+0],kernels[15*25+2*5+1],kernels[15*25+2*5+2],kernels[15*25+2*5+3],kernels[15*25+2*5+4],kernels[15*25+3*5+0],kernels[15*25+3*5+1],kernels[15*25+3*5+2],kernels[15*25+3*5+3],kernels[15*25+3*5+4],kernels[15*25+4*5+0],kernels[15*25+4*5+1],kernels[15*25+4*5+2],kernels[15*25+4*5+3],kernels[15*25+4*5+4],kernels[16*25+0*5+0],kernels[16*25+0*5+1],kernels[16*25+0*5+2],kernels[16*25+0*5+3],kernels[16*25+0*5+4],kernels[16*25+1*5+0],kernels[16*25+1*5+1],kernels[16*25+1*5+2],kernels[16*25+1*5+3],kernels[16*25+1*5+4],kernels[16*25+2*5+0],kernels[16*25+2*5+1],kernels[16*25+2*5+2],kernels[16*25+2*5+3],kernels[16*25+2*5+4],kernels[16*25+3*5+0],kernels[16*25+3*5+1],kernels[16*25+3*5+2],kernels[16*25+3*5+3],kernels[16*25+3*5+4],kernels[16*25+4*5+0],kernels[16*25+4*5+1],kernels[16*25+4*5+2],kernels[16*25+4*5+3],kernels[16*25+4*5+4],kernels[17*25+0*5+0],kernels[17*25+0*5+1],kernels[17*25+0*5+2],kernels[17*25+0*5+3],kernels[17*25+0*5+4],kernels[17*25+1*5+0],kernels[17*25+1*5+1],kernels[17*25+1*5+2],kernels[17*25+1*5+3],kernels[17*25+1*5+4],kernels[17*25+2*5+0],kernels[17*25+2*5+1],kernels[17*25+2*5+2],kernels[17*25+2*5+3],kernels[17*25+2*5+4],kernels[17*25+3*5+0],kernels[17*25+3*5+1],kernels[17*25+3*5+2],kernels[17*25+3*5+3],kernels[17*25+3*5+4],kernels[17*25+4*5+0],kernels[17*25+4*5+1],kernels[17*25+4*5+2],kernels[17*25+4*5+3],kernels[17*25+4*5+4]};

logic [0:chan*5*5-1] xnor1, xnor2, xnor3, xnor4;
assign xnor1 = image_slice1 ~^ kernel_slice;
assign xnor2 = image_slice2 ~^ kernel_slice;
assign xnor3 = image_slice3 ~^ kernel_slice;
assign xnor4 = image_slice4 ~^ kernel_slice;

logic [bW-1:0] sum1;
logic [bW-1:0] sum2;
logic [bW-1:0] sum3;
logic [bW-1:0] sum4;

popadd450 p1 (.bits(xnor1), .cnt(sum1));
popadd450 p2 (.bits(xnor2), .cnt(sum2));
popadd450 p3 (.bits(xnor3), .cnt(sum3));
popadd450 p4 (.bits(xnor4), .cnt(sum4));

logic bin1, bin2, bin3, bin4;

assign bin1 = sum1 > offset;
assign bin2 = sum2 > offset;
assign bin3 = sum3 > offset;
assign bin4 = sum4 > offset;

assign pixel = bin1 | bin2 | bin3 | bin4;


endmodule
