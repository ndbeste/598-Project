module conv1(
    input  logic image           [0:27][0:27],
    input  logic kernels         [0:99][0: 4][0: 4],
    output logic conv_one_out    [0:19][0:23][0:23]
    );

logic       xor_out [0:99][0:23][0:23];
logic [2:0] sum_out [0:19][0:23][0:23];

convchan1 c_1_0 (.image, .kernel(kernels[0]), .out_fmap(xor_out[0]));
convchan1 c_1_1 (.image, .kernel(kernels[1]), .out_fmap(xor_out[1]));
convchan1 c_1_2 (.image, .kernel(kernels[2]), .out_fmap(xor_out[2]));
convchan1 c_1_3 (.image, .kernel(kernels[3]), .out_fmap(xor_out[3]));
convchan1 c_1_4 (.image, .kernel(kernels[4]), .out_fmap(xor_out[4]));
convchan1 c_1_5 (.image, .kernel(kernels[5]), .out_fmap(xor_out[5]));
convchan1 c_1_6 (.image, .kernel(kernels[6]), .out_fmap(xor_out[6]));
convchan1 c_1_7 (.image, .kernel(kernels[7]), .out_fmap(xor_out[7]));
convchan1 c_1_8 (.image, .kernel(kernels[8]), .out_fmap(xor_out[8]));
convchan1 c_1_9 (.image, .kernel(kernels[9]), .out_fmap(xor_out[9]));
convchan1 c_1_10 (.image, .kernel(kernels[10]), .out_fmap(xor_out[10]));
convchan1 c_1_11 (.image, .kernel(kernels[11]), .out_fmap(xor_out[11]));
convchan1 c_1_12 (.image, .kernel(kernels[12]), .out_fmap(xor_out[12]));
convchan1 c_1_13 (.image, .kernel(kernels[13]), .out_fmap(xor_out[13]));
convchan1 c_1_14 (.image, .kernel(kernels[14]), .out_fmap(xor_out[14]));
convchan1 c_1_15 (.image, .kernel(kernels[15]), .out_fmap(xor_out[15]));
convchan1 c_1_16 (.image, .kernel(kernels[16]), .out_fmap(xor_out[16]));
convchan1 c_1_17 (.image, .kernel(kernels[17]), .out_fmap(xor_out[17]));
convchan1 c_1_18 (.image, .kernel(kernels[18]), .out_fmap(xor_out[18]));
convchan1 c_1_19 (.image, .kernel(kernels[19]), .out_fmap(xor_out[19]));
convchan1 c_1_20 (.image, .kernel(kernels[20]), .out_fmap(xor_out[20]));
convchan1 c_1_21 (.image, .kernel(kernels[21]), .out_fmap(xor_out[21]));
convchan1 c_1_22 (.image, .kernel(kernels[22]), .out_fmap(xor_out[22]));
convchan1 c_1_23 (.image, .kernel(kernels[23]), .out_fmap(xor_out[23]));
convchan1 c_1_24 (.image, .kernel(kernels[24]), .out_fmap(xor_out[24]));
convchan1 c_1_25 (.image, .kernel(kernels[25]), .out_fmap(xor_out[25]));
convchan1 c_1_26 (.image, .kernel(kernels[26]), .out_fmap(xor_out[26]));
convchan1 c_1_27 (.image, .kernel(kernels[27]), .out_fmap(xor_out[27]));
convchan1 c_1_28 (.image, .kernel(kernels[28]), .out_fmap(xor_out[28]));
convchan1 c_1_29 (.image, .kernel(kernels[29]), .out_fmap(xor_out[29]));
convchan1 c_1_30 (.image, .kernel(kernels[30]), .out_fmap(xor_out[30]));
convchan1 c_1_31 (.image, .kernel(kernels[31]), .out_fmap(xor_out[31]));
convchan1 c_1_32 (.image, .kernel(kernels[32]), .out_fmap(xor_out[32]));
convchan1 c_1_33 (.image, .kernel(kernels[33]), .out_fmap(xor_out[33]));
convchan1 c_1_34 (.image, .kernel(kernels[34]), .out_fmap(xor_out[34]));
convchan1 c_1_35 (.image, .kernel(kernels[35]), .out_fmap(xor_out[35]));
convchan1 c_1_36 (.image, .kernel(kernels[36]), .out_fmap(xor_out[36]));
convchan1 c_1_37 (.image, .kernel(kernels[37]), .out_fmap(xor_out[37]));
convchan1 c_1_38 (.image, .kernel(kernels[38]), .out_fmap(xor_out[38]));
convchan1 c_1_39 (.image, .kernel(kernels[39]), .out_fmap(xor_out[39]));
convchan1 c_1_40 (.image, .kernel(kernels[40]), .out_fmap(xor_out[40]));
convchan1 c_1_41 (.image, .kernel(kernels[41]), .out_fmap(xor_out[41]));
convchan1 c_1_42 (.image, .kernel(kernels[42]), .out_fmap(xor_out[42]));
convchan1 c_1_43 (.image, .kernel(kernels[43]), .out_fmap(xor_out[43]));
convchan1 c_1_44 (.image, .kernel(kernels[44]), .out_fmap(xor_out[44]));
convchan1 c_1_45 (.image, .kernel(kernels[45]), .out_fmap(xor_out[45]));
convchan1 c_1_46 (.image, .kernel(kernels[46]), .out_fmap(xor_out[46]));
convchan1 c_1_47 (.image, .kernel(kernels[47]), .out_fmap(xor_out[47]));
convchan1 c_1_48 (.image, .kernel(kernels[48]), .out_fmap(xor_out[48]));
convchan1 c_1_49 (.image, .kernel(kernels[49]), .out_fmap(xor_out[49]));
convchan1 c_1_50 (.image, .kernel(kernels[50]), .out_fmap(xor_out[50]));
convchan1 c_1_51 (.image, .kernel(kernels[51]), .out_fmap(xor_out[51]));
convchan1 c_1_52 (.image, .kernel(kernels[52]), .out_fmap(xor_out[52]));
convchan1 c_1_53 (.image, .kernel(kernels[53]), .out_fmap(xor_out[53]));
convchan1 c_1_54 (.image, .kernel(kernels[54]), .out_fmap(xor_out[54]));
convchan1 c_1_55 (.image, .kernel(kernels[55]), .out_fmap(xor_out[55]));
convchan1 c_1_56 (.image, .kernel(kernels[56]), .out_fmap(xor_out[56]));
convchan1 c_1_57 (.image, .kernel(kernels[57]), .out_fmap(xor_out[57]));
convchan1 c_1_58 (.image, .kernel(kernels[58]), .out_fmap(xor_out[58]));
convchan1 c_1_59 (.image, .kernel(kernels[59]), .out_fmap(xor_out[59]));
convchan1 c_1_60 (.image, .kernel(kernels[60]), .out_fmap(xor_out[60]));
convchan1 c_1_61 (.image, .kernel(kernels[61]), .out_fmap(xor_out[61]));
convchan1 c_1_62 (.image, .kernel(kernels[62]), .out_fmap(xor_out[62]));
convchan1 c_1_63 (.image, .kernel(kernels[63]), .out_fmap(xor_out[63]));
convchan1 c_1_64 (.image, .kernel(kernels[64]), .out_fmap(xor_out[64]));
convchan1 c_1_65 (.image, .kernel(kernels[65]), .out_fmap(xor_out[65]));
convchan1 c_1_66 (.image, .kernel(kernels[66]), .out_fmap(xor_out[66]));
convchan1 c_1_67 (.image, .kernel(kernels[67]), .out_fmap(xor_out[67]));
convchan1 c_1_68 (.image, .kernel(kernels[68]), .out_fmap(xor_out[68]));
convchan1 c_1_69 (.image, .kernel(kernels[69]), .out_fmap(xor_out[69]));
convchan1 c_1_70 (.image, .kernel(kernels[70]), .out_fmap(xor_out[70]));
convchan1 c_1_71 (.image, .kernel(kernels[71]), .out_fmap(xor_out[71]));
convchan1 c_1_72 (.image, .kernel(kernels[72]), .out_fmap(xor_out[72]));
convchan1 c_1_73 (.image, .kernel(kernels[73]), .out_fmap(xor_out[73]));
convchan1 c_1_74 (.image, .kernel(kernels[74]), .out_fmap(xor_out[74]));
convchan1 c_1_75 (.image, .kernel(kernels[75]), .out_fmap(xor_out[75]));
convchan1 c_1_76 (.image, .kernel(kernels[76]), .out_fmap(xor_out[76]));
convchan1 c_1_77 (.image, .kernel(kernels[77]), .out_fmap(xor_out[77]));
convchan1 c_1_78 (.image, .kernel(kernels[78]), .out_fmap(xor_out[78]));
convchan1 c_1_79 (.image, .kernel(kernels[79]), .out_fmap(xor_out[79]));
convchan1 c_1_80 (.image, .kernel(kernels[80]), .out_fmap(xor_out[80]));
convchan1 c_1_81 (.image, .kernel(kernels[81]), .out_fmap(xor_out[81]));
convchan1 c_1_82 (.image, .kernel(kernels[82]), .out_fmap(xor_out[82]));
convchan1 c_1_83 (.image, .kernel(kernels[83]), .out_fmap(xor_out[83]));
convchan1 c_1_84 (.image, .kernel(kernels[84]), .out_fmap(xor_out[84]));
convchan1 c_1_85 (.image, .kernel(kernels[85]), .out_fmap(xor_out[85]));
convchan1 c_1_86 (.image, .kernel(kernels[86]), .out_fmap(xor_out[86]));
convchan1 c_1_87 (.image, .kernel(kernels[87]), .out_fmap(xor_out[87]));
convchan1 c_1_88 (.image, .kernel(kernels[88]), .out_fmap(xor_out[88]));
convchan1 c_1_89 (.image, .kernel(kernels[89]), .out_fmap(xor_out[89]));
convchan1 c_1_90 (.image, .kernel(kernels[90]), .out_fmap(xor_out[90]));
convchan1 c_1_91 (.image, .kernel(kernels[91]), .out_fmap(xor_out[91]));
convchan1 c_1_92 (.image, .kernel(kernels[92]), .out_fmap(xor_out[92]));
convchan1 c_1_93 (.image, .kernel(kernels[93]), .out_fmap(xor_out[93]));
convchan1 c_1_94 (.image, .kernel(kernels[94]), .out_fmap(xor_out[94]));
convchan1 c_1_95 (.image, .kernel(kernels[95]), .out_fmap(xor_out[95]));
convchan1 c_1_96 (.image, .kernel(kernels[96]), .out_fmap(xor_out[96]));
convchan1 c_1_97 (.image, .kernel(kernels[97]), .out_fmap(xor_out[97]));
convchan1 c_1_98 (.image, .kernel(kernels[98]), .out_fmap(xor_out[98]));
convchan1 c_1_99 (.image, .kernel(kernels[99]), .out_fmap(xor_out[99]));

assign sum_out[0][0][0] = xor_out[0][0][0] + xor_out[1][0][0] + xor_out[2][0][0] + xor_out[3][0][0] + xor_out[4][0][0];
assign sum_out[1][0][0] = xor_out[5][0][0] + xor_out[6][0][0] + xor_out[7][0][0] + xor_out[8][0][0] + xor_out[9][0][0];
assign sum_out[2][0][0] = xor_out[10][0][0] + xor_out[11][0][0] + xor_out[12][0][0] + xor_out[13][0][0] + xor_out[14][0][0];
assign sum_out[3][0][0] = xor_out[15][0][0] + xor_out[16][0][0] + xor_out[17][0][0] + xor_out[18][0][0] + xor_out[19][0][0];
assign sum_out[4][0][0] = xor_out[20][0][0] + xor_out[21][0][0] + xor_out[22][0][0] + xor_out[23][0][0] + xor_out[24][0][0];
assign sum_out[5][0][0] = xor_out[25][0][0] + xor_out[26][0][0] + xor_out[27][0][0] + xor_out[28][0][0] + xor_out[29][0][0];
assign sum_out[6][0][0] = xor_out[30][0][0] + xor_out[31][0][0] + xor_out[32][0][0] + xor_out[33][0][0] + xor_out[34][0][0];
assign sum_out[7][0][0] = xor_out[35][0][0] + xor_out[36][0][0] + xor_out[37][0][0] + xor_out[38][0][0] + xor_out[39][0][0];
assign sum_out[8][0][0] = xor_out[40][0][0] + xor_out[41][0][0] + xor_out[42][0][0] + xor_out[43][0][0] + xor_out[44][0][0];
assign sum_out[9][0][0] = xor_out[45][0][0] + xor_out[46][0][0] + xor_out[47][0][0] + xor_out[48][0][0] + xor_out[49][0][0];
assign sum_out[10][0][0] = xor_out[50][0][0] + xor_out[51][0][0] + xor_out[52][0][0] + xor_out[53][0][0] + xor_out[54][0][0];
assign sum_out[11][0][0] = xor_out[55][0][0] + xor_out[56][0][0] + xor_out[57][0][0] + xor_out[58][0][0] + xor_out[59][0][0];
assign sum_out[12][0][0] = xor_out[60][0][0] + xor_out[61][0][0] + xor_out[62][0][0] + xor_out[63][0][0] + xor_out[64][0][0];
assign sum_out[13][0][0] = xor_out[65][0][0] + xor_out[66][0][0] + xor_out[67][0][0] + xor_out[68][0][0] + xor_out[69][0][0];
assign sum_out[14][0][0] = xor_out[70][0][0] + xor_out[71][0][0] + xor_out[72][0][0] + xor_out[73][0][0] + xor_out[74][0][0];
assign sum_out[15][0][0] = xor_out[75][0][0] + xor_out[76][0][0] + xor_out[77][0][0] + xor_out[78][0][0] + xor_out[79][0][0];
assign sum_out[16][0][0] = xor_out[80][0][0] + xor_out[81][0][0] + xor_out[82][0][0] + xor_out[83][0][0] + xor_out[84][0][0];
assign sum_out[17][0][0] = xor_out[85][0][0] + xor_out[86][0][0] + xor_out[87][0][0] + xor_out[88][0][0] + xor_out[89][0][0];
assign sum_out[18][0][0] = xor_out[90][0][0] + xor_out[91][0][0] + xor_out[92][0][0] + xor_out[93][0][0] + xor_out[94][0][0];
assign sum_out[19][0][0] = xor_out[95][0][0] + xor_out[96][0][0] + xor_out[97][0][0] + xor_out[98][0][0] + xor_out[99][0][0];

assign sum_out[0][0][1] = xor_out[0][0][1] + xor_out[1][0][1] + xor_out[2][0][1] + xor_out[3][0][1] + xor_out[4][0][1];
assign sum_out[1][0][1] = xor_out[5][0][1] + xor_out[6][0][1] + xor_out[7][0][1] + xor_out[8][0][1] + xor_out[9][0][1];
assign sum_out[2][0][1] = xor_out[10][0][1] + xor_out[11][0][1] + xor_out[12][0][1] + xor_out[13][0][1] + xor_out[14][0][1];
assign sum_out[3][0][1] = xor_out[15][0][1] + xor_out[16][0][1] + xor_out[17][0][1] + xor_out[18][0][1] + xor_out[19][0][1];
assign sum_out[4][0][1] = xor_out[20][0][1] + xor_out[21][0][1] + xor_out[22][0][1] + xor_out[23][0][1] + xor_out[24][0][1];
assign sum_out[5][0][1] = xor_out[25][0][1] + xor_out[26][0][1] + xor_out[27][0][1] + xor_out[28][0][1] + xor_out[29][0][1];
assign sum_out[6][0][1] = xor_out[30][0][1] + xor_out[31][0][1] + xor_out[32][0][1] + xor_out[33][0][1] + xor_out[34][0][1];
assign sum_out[7][0][1] = xor_out[35][0][1] + xor_out[36][0][1] + xor_out[37][0][1] + xor_out[38][0][1] + xor_out[39][0][1];
assign sum_out[8][0][1] = xor_out[40][0][1] + xor_out[41][0][1] + xor_out[42][0][1] + xor_out[43][0][1] + xor_out[44][0][1];
assign sum_out[9][0][1] = xor_out[45][0][1] + xor_out[46][0][1] + xor_out[47][0][1] + xor_out[48][0][1] + xor_out[49][0][1];
assign sum_out[10][0][1] = xor_out[50][0][1] + xor_out[51][0][1] + xor_out[52][0][1] + xor_out[53][0][1] + xor_out[54][0][1];
assign sum_out[11][0][1] = xor_out[55][0][1] + xor_out[56][0][1] + xor_out[57][0][1] + xor_out[58][0][1] + xor_out[59][0][1];
assign sum_out[12][0][1] = xor_out[60][0][1] + xor_out[61][0][1] + xor_out[62][0][1] + xor_out[63][0][1] + xor_out[64][0][1];
assign sum_out[13][0][1] = xor_out[65][0][1] + xor_out[66][0][1] + xor_out[67][0][1] + xor_out[68][0][1] + xor_out[69][0][1];
assign sum_out[14][0][1] = xor_out[70][0][1] + xor_out[71][0][1] + xor_out[72][0][1] + xor_out[73][0][1] + xor_out[74][0][1];
assign sum_out[15][0][1] = xor_out[75][0][1] + xor_out[76][0][1] + xor_out[77][0][1] + xor_out[78][0][1] + xor_out[79][0][1];
assign sum_out[16][0][1] = xor_out[80][0][1] + xor_out[81][0][1] + xor_out[82][0][1] + xor_out[83][0][1] + xor_out[84][0][1];
assign sum_out[17][0][1] = xor_out[85][0][1] + xor_out[86][0][1] + xor_out[87][0][1] + xor_out[88][0][1] + xor_out[89][0][1];
assign sum_out[18][0][1] = xor_out[90][0][1] + xor_out[91][0][1] + xor_out[92][0][1] + xor_out[93][0][1] + xor_out[94][0][1];
assign sum_out[19][0][1] = xor_out[95][0][1] + xor_out[96][0][1] + xor_out[97][0][1] + xor_out[98][0][1] + xor_out[99][0][1];

assign sum_out[0][0][2] = xor_out[0][0][2] + xor_out[1][0][2] + xor_out[2][0][2] + xor_out[3][0][2] + xor_out[4][0][2];
assign sum_out[1][0][2] = xor_out[5][0][2] + xor_out[6][0][2] + xor_out[7][0][2] + xor_out[8][0][2] + xor_out[9][0][2];
assign sum_out[2][0][2] = xor_out[10][0][2] + xor_out[11][0][2] + xor_out[12][0][2] + xor_out[13][0][2] + xor_out[14][0][2];
assign sum_out[3][0][2] = xor_out[15][0][2] + xor_out[16][0][2] + xor_out[17][0][2] + xor_out[18][0][2] + xor_out[19][0][2];
assign sum_out[4][0][2] = xor_out[20][0][2] + xor_out[21][0][2] + xor_out[22][0][2] + xor_out[23][0][2] + xor_out[24][0][2];
assign sum_out[5][0][2] = xor_out[25][0][2] + xor_out[26][0][2] + xor_out[27][0][2] + xor_out[28][0][2] + xor_out[29][0][2];
assign sum_out[6][0][2] = xor_out[30][0][2] + xor_out[31][0][2] + xor_out[32][0][2] + xor_out[33][0][2] + xor_out[34][0][2];
assign sum_out[7][0][2] = xor_out[35][0][2] + xor_out[36][0][2] + xor_out[37][0][2] + xor_out[38][0][2] + xor_out[39][0][2];
assign sum_out[8][0][2] = xor_out[40][0][2] + xor_out[41][0][2] + xor_out[42][0][2] + xor_out[43][0][2] + xor_out[44][0][2];
assign sum_out[9][0][2] = xor_out[45][0][2] + xor_out[46][0][2] + xor_out[47][0][2] + xor_out[48][0][2] + xor_out[49][0][2];
assign sum_out[10][0][2] = xor_out[50][0][2] + xor_out[51][0][2] + xor_out[52][0][2] + xor_out[53][0][2] + xor_out[54][0][2];
assign sum_out[11][0][2] = xor_out[55][0][2] + xor_out[56][0][2] + xor_out[57][0][2] + xor_out[58][0][2] + xor_out[59][0][2];
assign sum_out[12][0][2] = xor_out[60][0][2] + xor_out[61][0][2] + xor_out[62][0][2] + xor_out[63][0][2] + xor_out[64][0][2];
assign sum_out[13][0][2] = xor_out[65][0][2] + xor_out[66][0][2] + xor_out[67][0][2] + xor_out[68][0][2] + xor_out[69][0][2];
assign sum_out[14][0][2] = xor_out[70][0][2] + xor_out[71][0][2] + xor_out[72][0][2] + xor_out[73][0][2] + xor_out[74][0][2];
assign sum_out[15][0][2] = xor_out[75][0][2] + xor_out[76][0][2] + xor_out[77][0][2] + xor_out[78][0][2] + xor_out[79][0][2];
assign sum_out[16][0][2] = xor_out[80][0][2] + xor_out[81][0][2] + xor_out[82][0][2] + xor_out[83][0][2] + xor_out[84][0][2];
assign sum_out[17][0][2] = xor_out[85][0][2] + xor_out[86][0][2] + xor_out[87][0][2] + xor_out[88][0][2] + xor_out[89][0][2];
assign sum_out[18][0][2] = xor_out[90][0][2] + xor_out[91][0][2] + xor_out[92][0][2] + xor_out[93][0][2] + xor_out[94][0][2];
assign sum_out[19][0][2] = xor_out[95][0][2] + xor_out[96][0][2] + xor_out[97][0][2] + xor_out[98][0][2] + xor_out[99][0][2];

assign sum_out[0][0][3] = xor_out[0][0][3] + xor_out[1][0][3] + xor_out[2][0][3] + xor_out[3][0][3] + xor_out[4][0][3];
assign sum_out[1][0][3] = xor_out[5][0][3] + xor_out[6][0][3] + xor_out[7][0][3] + xor_out[8][0][3] + xor_out[9][0][3];
assign sum_out[2][0][3] = xor_out[10][0][3] + xor_out[11][0][3] + xor_out[12][0][3] + xor_out[13][0][3] + xor_out[14][0][3];
assign sum_out[3][0][3] = xor_out[15][0][3] + xor_out[16][0][3] + xor_out[17][0][3] + xor_out[18][0][3] + xor_out[19][0][3];
assign sum_out[4][0][3] = xor_out[20][0][3] + xor_out[21][0][3] + xor_out[22][0][3] + xor_out[23][0][3] + xor_out[24][0][3];
assign sum_out[5][0][3] = xor_out[25][0][3] + xor_out[26][0][3] + xor_out[27][0][3] + xor_out[28][0][3] + xor_out[29][0][3];
assign sum_out[6][0][3] = xor_out[30][0][3] + xor_out[31][0][3] + xor_out[32][0][3] + xor_out[33][0][3] + xor_out[34][0][3];
assign sum_out[7][0][3] = xor_out[35][0][3] + xor_out[36][0][3] + xor_out[37][0][3] + xor_out[38][0][3] + xor_out[39][0][3];
assign sum_out[8][0][3] = xor_out[40][0][3] + xor_out[41][0][3] + xor_out[42][0][3] + xor_out[43][0][3] + xor_out[44][0][3];
assign sum_out[9][0][3] = xor_out[45][0][3] + xor_out[46][0][3] + xor_out[47][0][3] + xor_out[48][0][3] + xor_out[49][0][3];
assign sum_out[10][0][3] = xor_out[50][0][3] + xor_out[51][0][3] + xor_out[52][0][3] + xor_out[53][0][3] + xor_out[54][0][3];
assign sum_out[11][0][3] = xor_out[55][0][3] + xor_out[56][0][3] + xor_out[57][0][3] + xor_out[58][0][3] + xor_out[59][0][3];
assign sum_out[12][0][3] = xor_out[60][0][3] + xor_out[61][0][3] + xor_out[62][0][3] + xor_out[63][0][3] + xor_out[64][0][3];
assign sum_out[13][0][3] = xor_out[65][0][3] + xor_out[66][0][3] + xor_out[67][0][3] + xor_out[68][0][3] + xor_out[69][0][3];
assign sum_out[14][0][3] = xor_out[70][0][3] + xor_out[71][0][3] + xor_out[72][0][3] + xor_out[73][0][3] + xor_out[74][0][3];
assign sum_out[15][0][3] = xor_out[75][0][3] + xor_out[76][0][3] + xor_out[77][0][3] + xor_out[78][0][3] + xor_out[79][0][3];
assign sum_out[16][0][3] = xor_out[80][0][3] + xor_out[81][0][3] + xor_out[82][0][3] + xor_out[83][0][3] + xor_out[84][0][3];
assign sum_out[17][0][3] = xor_out[85][0][3] + xor_out[86][0][3] + xor_out[87][0][3] + xor_out[88][0][3] + xor_out[89][0][3];
assign sum_out[18][0][3] = xor_out[90][0][3] + xor_out[91][0][3] + xor_out[92][0][3] + xor_out[93][0][3] + xor_out[94][0][3];
assign sum_out[19][0][3] = xor_out[95][0][3] + xor_out[96][0][3] + xor_out[97][0][3] + xor_out[98][0][3] + xor_out[99][0][3];

assign sum_out[0][0][4] = xor_out[0][0][4] + xor_out[1][0][4] + xor_out[2][0][4] + xor_out[3][0][4] + xor_out[4][0][4];
assign sum_out[1][0][4] = xor_out[5][0][4] + xor_out[6][0][4] + xor_out[7][0][4] + xor_out[8][0][4] + xor_out[9][0][4];
assign sum_out[2][0][4] = xor_out[10][0][4] + xor_out[11][0][4] + xor_out[12][0][4] + xor_out[13][0][4] + xor_out[14][0][4];
assign sum_out[3][0][4] = xor_out[15][0][4] + xor_out[16][0][4] + xor_out[17][0][4] + xor_out[18][0][4] + xor_out[19][0][4];
assign sum_out[4][0][4] = xor_out[20][0][4] + xor_out[21][0][4] + xor_out[22][0][4] + xor_out[23][0][4] + xor_out[24][0][4];
assign sum_out[5][0][4] = xor_out[25][0][4] + xor_out[26][0][4] + xor_out[27][0][4] + xor_out[28][0][4] + xor_out[29][0][4];
assign sum_out[6][0][4] = xor_out[30][0][4] + xor_out[31][0][4] + xor_out[32][0][4] + xor_out[33][0][4] + xor_out[34][0][4];
assign sum_out[7][0][4] = xor_out[35][0][4] + xor_out[36][0][4] + xor_out[37][0][4] + xor_out[38][0][4] + xor_out[39][0][4];
assign sum_out[8][0][4] = xor_out[40][0][4] + xor_out[41][0][4] + xor_out[42][0][4] + xor_out[43][0][4] + xor_out[44][0][4];
assign sum_out[9][0][4] = xor_out[45][0][4] + xor_out[46][0][4] + xor_out[47][0][4] + xor_out[48][0][4] + xor_out[49][0][4];
assign sum_out[10][0][4] = xor_out[50][0][4] + xor_out[51][0][4] + xor_out[52][0][4] + xor_out[53][0][4] + xor_out[54][0][4];
assign sum_out[11][0][4] = xor_out[55][0][4] + xor_out[56][0][4] + xor_out[57][0][4] + xor_out[58][0][4] + xor_out[59][0][4];
assign sum_out[12][0][4] = xor_out[60][0][4] + xor_out[61][0][4] + xor_out[62][0][4] + xor_out[63][0][4] + xor_out[64][0][4];
assign sum_out[13][0][4] = xor_out[65][0][4] + xor_out[66][0][4] + xor_out[67][0][4] + xor_out[68][0][4] + xor_out[69][0][4];
assign sum_out[14][0][4] = xor_out[70][0][4] + xor_out[71][0][4] + xor_out[72][0][4] + xor_out[73][0][4] + xor_out[74][0][4];
assign sum_out[15][0][4] = xor_out[75][0][4] + xor_out[76][0][4] + xor_out[77][0][4] + xor_out[78][0][4] + xor_out[79][0][4];
assign sum_out[16][0][4] = xor_out[80][0][4] + xor_out[81][0][4] + xor_out[82][0][4] + xor_out[83][0][4] + xor_out[84][0][4];
assign sum_out[17][0][4] = xor_out[85][0][4] + xor_out[86][0][4] + xor_out[87][0][4] + xor_out[88][0][4] + xor_out[89][0][4];
assign sum_out[18][0][4] = xor_out[90][0][4] + xor_out[91][0][4] + xor_out[92][0][4] + xor_out[93][0][4] + xor_out[94][0][4];
assign sum_out[19][0][4] = xor_out[95][0][4] + xor_out[96][0][4] + xor_out[97][0][4] + xor_out[98][0][4] + xor_out[99][0][4];

assign sum_out[0][0][5] = xor_out[0][0][5] + xor_out[1][0][5] + xor_out[2][0][5] + xor_out[3][0][5] + xor_out[4][0][5];
assign sum_out[1][0][5] = xor_out[5][0][5] + xor_out[6][0][5] + xor_out[7][0][5] + xor_out[8][0][5] + xor_out[9][0][5];
assign sum_out[2][0][5] = xor_out[10][0][5] + xor_out[11][0][5] + xor_out[12][0][5] + xor_out[13][0][5] + xor_out[14][0][5];
assign sum_out[3][0][5] = xor_out[15][0][5] + xor_out[16][0][5] + xor_out[17][0][5] + xor_out[18][0][5] + xor_out[19][0][5];
assign sum_out[4][0][5] = xor_out[20][0][5] + xor_out[21][0][5] + xor_out[22][0][5] + xor_out[23][0][5] + xor_out[24][0][5];
assign sum_out[5][0][5] = xor_out[25][0][5] + xor_out[26][0][5] + xor_out[27][0][5] + xor_out[28][0][5] + xor_out[29][0][5];
assign sum_out[6][0][5] = xor_out[30][0][5] + xor_out[31][0][5] + xor_out[32][0][5] + xor_out[33][0][5] + xor_out[34][0][5];
assign sum_out[7][0][5] = xor_out[35][0][5] + xor_out[36][0][5] + xor_out[37][0][5] + xor_out[38][0][5] + xor_out[39][0][5];
assign sum_out[8][0][5] = xor_out[40][0][5] + xor_out[41][0][5] + xor_out[42][0][5] + xor_out[43][0][5] + xor_out[44][0][5];
assign sum_out[9][0][5] = xor_out[45][0][5] + xor_out[46][0][5] + xor_out[47][0][5] + xor_out[48][0][5] + xor_out[49][0][5];
assign sum_out[10][0][5] = xor_out[50][0][5] + xor_out[51][0][5] + xor_out[52][0][5] + xor_out[53][0][5] + xor_out[54][0][5];
assign sum_out[11][0][5] = xor_out[55][0][5] + xor_out[56][0][5] + xor_out[57][0][5] + xor_out[58][0][5] + xor_out[59][0][5];
assign sum_out[12][0][5] = xor_out[60][0][5] + xor_out[61][0][5] + xor_out[62][0][5] + xor_out[63][0][5] + xor_out[64][0][5];
assign sum_out[13][0][5] = xor_out[65][0][5] + xor_out[66][0][5] + xor_out[67][0][5] + xor_out[68][0][5] + xor_out[69][0][5];
assign sum_out[14][0][5] = xor_out[70][0][5] + xor_out[71][0][5] + xor_out[72][0][5] + xor_out[73][0][5] + xor_out[74][0][5];
assign sum_out[15][0][5] = xor_out[75][0][5] + xor_out[76][0][5] + xor_out[77][0][5] + xor_out[78][0][5] + xor_out[79][0][5];
assign sum_out[16][0][5] = xor_out[80][0][5] + xor_out[81][0][5] + xor_out[82][0][5] + xor_out[83][0][5] + xor_out[84][0][5];
assign sum_out[17][0][5] = xor_out[85][0][5] + xor_out[86][0][5] + xor_out[87][0][5] + xor_out[88][0][5] + xor_out[89][0][5];
assign sum_out[18][0][5] = xor_out[90][0][5] + xor_out[91][0][5] + xor_out[92][0][5] + xor_out[93][0][5] + xor_out[94][0][5];
assign sum_out[19][0][5] = xor_out[95][0][5] + xor_out[96][0][5] + xor_out[97][0][5] + xor_out[98][0][5] + xor_out[99][0][5];

assign sum_out[0][0][6] = xor_out[0][0][6] + xor_out[1][0][6] + xor_out[2][0][6] + xor_out[3][0][6] + xor_out[4][0][6];
assign sum_out[1][0][6] = xor_out[5][0][6] + xor_out[6][0][6] + xor_out[7][0][6] + xor_out[8][0][6] + xor_out[9][0][6];
assign sum_out[2][0][6] = xor_out[10][0][6] + xor_out[11][0][6] + xor_out[12][0][6] + xor_out[13][0][6] + xor_out[14][0][6];
assign sum_out[3][0][6] = xor_out[15][0][6] + xor_out[16][0][6] + xor_out[17][0][6] + xor_out[18][0][6] + xor_out[19][0][6];
assign sum_out[4][0][6] = xor_out[20][0][6] + xor_out[21][0][6] + xor_out[22][0][6] + xor_out[23][0][6] + xor_out[24][0][6];
assign sum_out[5][0][6] = xor_out[25][0][6] + xor_out[26][0][6] + xor_out[27][0][6] + xor_out[28][0][6] + xor_out[29][0][6];
assign sum_out[6][0][6] = xor_out[30][0][6] + xor_out[31][0][6] + xor_out[32][0][6] + xor_out[33][0][6] + xor_out[34][0][6];
assign sum_out[7][0][6] = xor_out[35][0][6] + xor_out[36][0][6] + xor_out[37][0][6] + xor_out[38][0][6] + xor_out[39][0][6];
assign sum_out[8][0][6] = xor_out[40][0][6] + xor_out[41][0][6] + xor_out[42][0][6] + xor_out[43][0][6] + xor_out[44][0][6];
assign sum_out[9][0][6] = xor_out[45][0][6] + xor_out[46][0][6] + xor_out[47][0][6] + xor_out[48][0][6] + xor_out[49][0][6];
assign sum_out[10][0][6] = xor_out[50][0][6] + xor_out[51][0][6] + xor_out[52][0][6] + xor_out[53][0][6] + xor_out[54][0][6];
assign sum_out[11][0][6] = xor_out[55][0][6] + xor_out[56][0][6] + xor_out[57][0][6] + xor_out[58][0][6] + xor_out[59][0][6];
assign sum_out[12][0][6] = xor_out[60][0][6] + xor_out[61][0][6] + xor_out[62][0][6] + xor_out[63][0][6] + xor_out[64][0][6];
assign sum_out[13][0][6] = xor_out[65][0][6] + xor_out[66][0][6] + xor_out[67][0][6] + xor_out[68][0][6] + xor_out[69][0][6];
assign sum_out[14][0][6] = xor_out[70][0][6] + xor_out[71][0][6] + xor_out[72][0][6] + xor_out[73][0][6] + xor_out[74][0][6];
assign sum_out[15][0][6] = xor_out[75][0][6] + xor_out[76][0][6] + xor_out[77][0][6] + xor_out[78][0][6] + xor_out[79][0][6];
assign sum_out[16][0][6] = xor_out[80][0][6] + xor_out[81][0][6] + xor_out[82][0][6] + xor_out[83][0][6] + xor_out[84][0][6];
assign sum_out[17][0][6] = xor_out[85][0][6] + xor_out[86][0][6] + xor_out[87][0][6] + xor_out[88][0][6] + xor_out[89][0][6];
assign sum_out[18][0][6] = xor_out[90][0][6] + xor_out[91][0][6] + xor_out[92][0][6] + xor_out[93][0][6] + xor_out[94][0][6];
assign sum_out[19][0][6] = xor_out[95][0][6] + xor_out[96][0][6] + xor_out[97][0][6] + xor_out[98][0][6] + xor_out[99][0][6];

assign sum_out[0][0][7] = xor_out[0][0][7] + xor_out[1][0][7] + xor_out[2][0][7] + xor_out[3][0][7] + xor_out[4][0][7];
assign sum_out[1][0][7] = xor_out[5][0][7] + xor_out[6][0][7] + xor_out[7][0][7] + xor_out[8][0][7] + xor_out[9][0][7];
assign sum_out[2][0][7] = xor_out[10][0][7] + xor_out[11][0][7] + xor_out[12][0][7] + xor_out[13][0][7] + xor_out[14][0][7];
assign sum_out[3][0][7] = xor_out[15][0][7] + xor_out[16][0][7] + xor_out[17][0][7] + xor_out[18][0][7] + xor_out[19][0][7];
assign sum_out[4][0][7] = xor_out[20][0][7] + xor_out[21][0][7] + xor_out[22][0][7] + xor_out[23][0][7] + xor_out[24][0][7];
assign sum_out[5][0][7] = xor_out[25][0][7] + xor_out[26][0][7] + xor_out[27][0][7] + xor_out[28][0][7] + xor_out[29][0][7];
assign sum_out[6][0][7] = xor_out[30][0][7] + xor_out[31][0][7] + xor_out[32][0][7] + xor_out[33][0][7] + xor_out[34][0][7];
assign sum_out[7][0][7] = xor_out[35][0][7] + xor_out[36][0][7] + xor_out[37][0][7] + xor_out[38][0][7] + xor_out[39][0][7];
assign sum_out[8][0][7] = xor_out[40][0][7] + xor_out[41][0][7] + xor_out[42][0][7] + xor_out[43][0][7] + xor_out[44][0][7];
assign sum_out[9][0][7] = xor_out[45][0][7] + xor_out[46][0][7] + xor_out[47][0][7] + xor_out[48][0][7] + xor_out[49][0][7];
assign sum_out[10][0][7] = xor_out[50][0][7] + xor_out[51][0][7] + xor_out[52][0][7] + xor_out[53][0][7] + xor_out[54][0][7];
assign sum_out[11][0][7] = xor_out[55][0][7] + xor_out[56][0][7] + xor_out[57][0][7] + xor_out[58][0][7] + xor_out[59][0][7];
assign sum_out[12][0][7] = xor_out[60][0][7] + xor_out[61][0][7] + xor_out[62][0][7] + xor_out[63][0][7] + xor_out[64][0][7];
assign sum_out[13][0][7] = xor_out[65][0][7] + xor_out[66][0][7] + xor_out[67][0][7] + xor_out[68][0][7] + xor_out[69][0][7];
assign sum_out[14][0][7] = xor_out[70][0][7] + xor_out[71][0][7] + xor_out[72][0][7] + xor_out[73][0][7] + xor_out[74][0][7];
assign sum_out[15][0][7] = xor_out[75][0][7] + xor_out[76][0][7] + xor_out[77][0][7] + xor_out[78][0][7] + xor_out[79][0][7];
assign sum_out[16][0][7] = xor_out[80][0][7] + xor_out[81][0][7] + xor_out[82][0][7] + xor_out[83][0][7] + xor_out[84][0][7];
assign sum_out[17][0][7] = xor_out[85][0][7] + xor_out[86][0][7] + xor_out[87][0][7] + xor_out[88][0][7] + xor_out[89][0][7];
assign sum_out[18][0][7] = xor_out[90][0][7] + xor_out[91][0][7] + xor_out[92][0][7] + xor_out[93][0][7] + xor_out[94][0][7];
assign sum_out[19][0][7] = xor_out[95][0][7] + xor_out[96][0][7] + xor_out[97][0][7] + xor_out[98][0][7] + xor_out[99][0][7];

assign sum_out[0][0][8] = xor_out[0][0][8] + xor_out[1][0][8] + xor_out[2][0][8] + xor_out[3][0][8] + xor_out[4][0][8];
assign sum_out[1][0][8] = xor_out[5][0][8] + xor_out[6][0][8] + xor_out[7][0][8] + xor_out[8][0][8] + xor_out[9][0][8];
assign sum_out[2][0][8] = xor_out[10][0][8] + xor_out[11][0][8] + xor_out[12][0][8] + xor_out[13][0][8] + xor_out[14][0][8];
assign sum_out[3][0][8] = xor_out[15][0][8] + xor_out[16][0][8] + xor_out[17][0][8] + xor_out[18][0][8] + xor_out[19][0][8];
assign sum_out[4][0][8] = xor_out[20][0][8] + xor_out[21][0][8] + xor_out[22][0][8] + xor_out[23][0][8] + xor_out[24][0][8];
assign sum_out[5][0][8] = xor_out[25][0][8] + xor_out[26][0][8] + xor_out[27][0][8] + xor_out[28][0][8] + xor_out[29][0][8];
assign sum_out[6][0][8] = xor_out[30][0][8] + xor_out[31][0][8] + xor_out[32][0][8] + xor_out[33][0][8] + xor_out[34][0][8];
assign sum_out[7][0][8] = xor_out[35][0][8] + xor_out[36][0][8] + xor_out[37][0][8] + xor_out[38][0][8] + xor_out[39][0][8];
assign sum_out[8][0][8] = xor_out[40][0][8] + xor_out[41][0][8] + xor_out[42][0][8] + xor_out[43][0][8] + xor_out[44][0][8];
assign sum_out[9][0][8] = xor_out[45][0][8] + xor_out[46][0][8] + xor_out[47][0][8] + xor_out[48][0][8] + xor_out[49][0][8];
assign sum_out[10][0][8] = xor_out[50][0][8] + xor_out[51][0][8] + xor_out[52][0][8] + xor_out[53][0][8] + xor_out[54][0][8];
assign sum_out[11][0][8] = xor_out[55][0][8] + xor_out[56][0][8] + xor_out[57][0][8] + xor_out[58][0][8] + xor_out[59][0][8];
assign sum_out[12][0][8] = xor_out[60][0][8] + xor_out[61][0][8] + xor_out[62][0][8] + xor_out[63][0][8] + xor_out[64][0][8];
assign sum_out[13][0][8] = xor_out[65][0][8] + xor_out[66][0][8] + xor_out[67][0][8] + xor_out[68][0][8] + xor_out[69][0][8];
assign sum_out[14][0][8] = xor_out[70][0][8] + xor_out[71][0][8] + xor_out[72][0][8] + xor_out[73][0][8] + xor_out[74][0][8];
assign sum_out[15][0][8] = xor_out[75][0][8] + xor_out[76][0][8] + xor_out[77][0][8] + xor_out[78][0][8] + xor_out[79][0][8];
assign sum_out[16][0][8] = xor_out[80][0][8] + xor_out[81][0][8] + xor_out[82][0][8] + xor_out[83][0][8] + xor_out[84][0][8];
assign sum_out[17][0][8] = xor_out[85][0][8] + xor_out[86][0][8] + xor_out[87][0][8] + xor_out[88][0][8] + xor_out[89][0][8];
assign sum_out[18][0][8] = xor_out[90][0][8] + xor_out[91][0][8] + xor_out[92][0][8] + xor_out[93][0][8] + xor_out[94][0][8];
assign sum_out[19][0][8] = xor_out[95][0][8] + xor_out[96][0][8] + xor_out[97][0][8] + xor_out[98][0][8] + xor_out[99][0][8];

assign sum_out[0][0][9] = xor_out[0][0][9] + xor_out[1][0][9] + xor_out[2][0][9] + xor_out[3][0][9] + xor_out[4][0][9];
assign sum_out[1][0][9] = xor_out[5][0][9] + xor_out[6][0][9] + xor_out[7][0][9] + xor_out[8][0][9] + xor_out[9][0][9];
assign sum_out[2][0][9] = xor_out[10][0][9] + xor_out[11][0][9] + xor_out[12][0][9] + xor_out[13][0][9] + xor_out[14][0][9];
assign sum_out[3][0][9] = xor_out[15][0][9] + xor_out[16][0][9] + xor_out[17][0][9] + xor_out[18][0][9] + xor_out[19][0][9];
assign sum_out[4][0][9] = xor_out[20][0][9] + xor_out[21][0][9] + xor_out[22][0][9] + xor_out[23][0][9] + xor_out[24][0][9];
assign sum_out[5][0][9] = xor_out[25][0][9] + xor_out[26][0][9] + xor_out[27][0][9] + xor_out[28][0][9] + xor_out[29][0][9];
assign sum_out[6][0][9] = xor_out[30][0][9] + xor_out[31][0][9] + xor_out[32][0][9] + xor_out[33][0][9] + xor_out[34][0][9];
assign sum_out[7][0][9] = xor_out[35][0][9] + xor_out[36][0][9] + xor_out[37][0][9] + xor_out[38][0][9] + xor_out[39][0][9];
assign sum_out[8][0][9] = xor_out[40][0][9] + xor_out[41][0][9] + xor_out[42][0][9] + xor_out[43][0][9] + xor_out[44][0][9];
assign sum_out[9][0][9] = xor_out[45][0][9] + xor_out[46][0][9] + xor_out[47][0][9] + xor_out[48][0][9] + xor_out[49][0][9];
assign sum_out[10][0][9] = xor_out[50][0][9] + xor_out[51][0][9] + xor_out[52][0][9] + xor_out[53][0][9] + xor_out[54][0][9];
assign sum_out[11][0][9] = xor_out[55][0][9] + xor_out[56][0][9] + xor_out[57][0][9] + xor_out[58][0][9] + xor_out[59][0][9];
assign sum_out[12][0][9] = xor_out[60][0][9] + xor_out[61][0][9] + xor_out[62][0][9] + xor_out[63][0][9] + xor_out[64][0][9];
assign sum_out[13][0][9] = xor_out[65][0][9] + xor_out[66][0][9] + xor_out[67][0][9] + xor_out[68][0][9] + xor_out[69][0][9];
assign sum_out[14][0][9] = xor_out[70][0][9] + xor_out[71][0][9] + xor_out[72][0][9] + xor_out[73][0][9] + xor_out[74][0][9];
assign sum_out[15][0][9] = xor_out[75][0][9] + xor_out[76][0][9] + xor_out[77][0][9] + xor_out[78][0][9] + xor_out[79][0][9];
assign sum_out[16][0][9] = xor_out[80][0][9] + xor_out[81][0][9] + xor_out[82][0][9] + xor_out[83][0][9] + xor_out[84][0][9];
assign sum_out[17][0][9] = xor_out[85][0][9] + xor_out[86][0][9] + xor_out[87][0][9] + xor_out[88][0][9] + xor_out[89][0][9];
assign sum_out[18][0][9] = xor_out[90][0][9] + xor_out[91][0][9] + xor_out[92][0][9] + xor_out[93][0][9] + xor_out[94][0][9];
assign sum_out[19][0][9] = xor_out[95][0][9] + xor_out[96][0][9] + xor_out[97][0][9] + xor_out[98][0][9] + xor_out[99][0][9];

assign sum_out[0][0][10] = xor_out[0][0][10] + xor_out[1][0][10] + xor_out[2][0][10] + xor_out[3][0][10] + xor_out[4][0][10];
assign sum_out[1][0][10] = xor_out[5][0][10] + xor_out[6][0][10] + xor_out[7][0][10] + xor_out[8][0][10] + xor_out[9][0][10];
assign sum_out[2][0][10] = xor_out[10][0][10] + xor_out[11][0][10] + xor_out[12][0][10] + xor_out[13][0][10] + xor_out[14][0][10];
assign sum_out[3][0][10] = xor_out[15][0][10] + xor_out[16][0][10] + xor_out[17][0][10] + xor_out[18][0][10] + xor_out[19][0][10];
assign sum_out[4][0][10] = xor_out[20][0][10] + xor_out[21][0][10] + xor_out[22][0][10] + xor_out[23][0][10] + xor_out[24][0][10];
assign sum_out[5][0][10] = xor_out[25][0][10] + xor_out[26][0][10] + xor_out[27][0][10] + xor_out[28][0][10] + xor_out[29][0][10];
assign sum_out[6][0][10] = xor_out[30][0][10] + xor_out[31][0][10] + xor_out[32][0][10] + xor_out[33][0][10] + xor_out[34][0][10];
assign sum_out[7][0][10] = xor_out[35][0][10] + xor_out[36][0][10] + xor_out[37][0][10] + xor_out[38][0][10] + xor_out[39][0][10];
assign sum_out[8][0][10] = xor_out[40][0][10] + xor_out[41][0][10] + xor_out[42][0][10] + xor_out[43][0][10] + xor_out[44][0][10];
assign sum_out[9][0][10] = xor_out[45][0][10] + xor_out[46][0][10] + xor_out[47][0][10] + xor_out[48][0][10] + xor_out[49][0][10];
assign sum_out[10][0][10] = xor_out[50][0][10] + xor_out[51][0][10] + xor_out[52][0][10] + xor_out[53][0][10] + xor_out[54][0][10];
assign sum_out[11][0][10] = xor_out[55][0][10] + xor_out[56][0][10] + xor_out[57][0][10] + xor_out[58][0][10] + xor_out[59][0][10];
assign sum_out[12][0][10] = xor_out[60][0][10] + xor_out[61][0][10] + xor_out[62][0][10] + xor_out[63][0][10] + xor_out[64][0][10];
assign sum_out[13][0][10] = xor_out[65][0][10] + xor_out[66][0][10] + xor_out[67][0][10] + xor_out[68][0][10] + xor_out[69][0][10];
assign sum_out[14][0][10] = xor_out[70][0][10] + xor_out[71][0][10] + xor_out[72][0][10] + xor_out[73][0][10] + xor_out[74][0][10];
assign sum_out[15][0][10] = xor_out[75][0][10] + xor_out[76][0][10] + xor_out[77][0][10] + xor_out[78][0][10] + xor_out[79][0][10];
assign sum_out[16][0][10] = xor_out[80][0][10] + xor_out[81][0][10] + xor_out[82][0][10] + xor_out[83][0][10] + xor_out[84][0][10];
assign sum_out[17][0][10] = xor_out[85][0][10] + xor_out[86][0][10] + xor_out[87][0][10] + xor_out[88][0][10] + xor_out[89][0][10];
assign sum_out[18][0][10] = xor_out[90][0][10] + xor_out[91][0][10] + xor_out[92][0][10] + xor_out[93][0][10] + xor_out[94][0][10];
assign sum_out[19][0][10] = xor_out[95][0][10] + xor_out[96][0][10] + xor_out[97][0][10] + xor_out[98][0][10] + xor_out[99][0][10];

assign sum_out[0][0][11] = xor_out[0][0][11] + xor_out[1][0][11] + xor_out[2][0][11] + xor_out[3][0][11] + xor_out[4][0][11];
assign sum_out[1][0][11] = xor_out[5][0][11] + xor_out[6][0][11] + xor_out[7][0][11] + xor_out[8][0][11] + xor_out[9][0][11];
assign sum_out[2][0][11] = xor_out[10][0][11] + xor_out[11][0][11] + xor_out[12][0][11] + xor_out[13][0][11] + xor_out[14][0][11];
assign sum_out[3][0][11] = xor_out[15][0][11] + xor_out[16][0][11] + xor_out[17][0][11] + xor_out[18][0][11] + xor_out[19][0][11];
assign sum_out[4][0][11] = xor_out[20][0][11] + xor_out[21][0][11] + xor_out[22][0][11] + xor_out[23][0][11] + xor_out[24][0][11];
assign sum_out[5][0][11] = xor_out[25][0][11] + xor_out[26][0][11] + xor_out[27][0][11] + xor_out[28][0][11] + xor_out[29][0][11];
assign sum_out[6][0][11] = xor_out[30][0][11] + xor_out[31][0][11] + xor_out[32][0][11] + xor_out[33][0][11] + xor_out[34][0][11];
assign sum_out[7][0][11] = xor_out[35][0][11] + xor_out[36][0][11] + xor_out[37][0][11] + xor_out[38][0][11] + xor_out[39][0][11];
assign sum_out[8][0][11] = xor_out[40][0][11] + xor_out[41][0][11] + xor_out[42][0][11] + xor_out[43][0][11] + xor_out[44][0][11];
assign sum_out[9][0][11] = xor_out[45][0][11] + xor_out[46][0][11] + xor_out[47][0][11] + xor_out[48][0][11] + xor_out[49][0][11];
assign sum_out[10][0][11] = xor_out[50][0][11] + xor_out[51][0][11] + xor_out[52][0][11] + xor_out[53][0][11] + xor_out[54][0][11];
assign sum_out[11][0][11] = xor_out[55][0][11] + xor_out[56][0][11] + xor_out[57][0][11] + xor_out[58][0][11] + xor_out[59][0][11];
assign sum_out[12][0][11] = xor_out[60][0][11] + xor_out[61][0][11] + xor_out[62][0][11] + xor_out[63][0][11] + xor_out[64][0][11];
assign sum_out[13][0][11] = xor_out[65][0][11] + xor_out[66][0][11] + xor_out[67][0][11] + xor_out[68][0][11] + xor_out[69][0][11];
assign sum_out[14][0][11] = xor_out[70][0][11] + xor_out[71][0][11] + xor_out[72][0][11] + xor_out[73][0][11] + xor_out[74][0][11];
assign sum_out[15][0][11] = xor_out[75][0][11] + xor_out[76][0][11] + xor_out[77][0][11] + xor_out[78][0][11] + xor_out[79][0][11];
assign sum_out[16][0][11] = xor_out[80][0][11] + xor_out[81][0][11] + xor_out[82][0][11] + xor_out[83][0][11] + xor_out[84][0][11];
assign sum_out[17][0][11] = xor_out[85][0][11] + xor_out[86][0][11] + xor_out[87][0][11] + xor_out[88][0][11] + xor_out[89][0][11];
assign sum_out[18][0][11] = xor_out[90][0][11] + xor_out[91][0][11] + xor_out[92][0][11] + xor_out[93][0][11] + xor_out[94][0][11];
assign sum_out[19][0][11] = xor_out[95][0][11] + xor_out[96][0][11] + xor_out[97][0][11] + xor_out[98][0][11] + xor_out[99][0][11];

assign sum_out[0][0][12] = xor_out[0][0][12] + xor_out[1][0][12] + xor_out[2][0][12] + xor_out[3][0][12] + xor_out[4][0][12];
assign sum_out[1][0][12] = xor_out[5][0][12] + xor_out[6][0][12] + xor_out[7][0][12] + xor_out[8][0][12] + xor_out[9][0][12];
assign sum_out[2][0][12] = xor_out[10][0][12] + xor_out[11][0][12] + xor_out[12][0][12] + xor_out[13][0][12] + xor_out[14][0][12];
assign sum_out[3][0][12] = xor_out[15][0][12] + xor_out[16][0][12] + xor_out[17][0][12] + xor_out[18][0][12] + xor_out[19][0][12];
assign sum_out[4][0][12] = xor_out[20][0][12] + xor_out[21][0][12] + xor_out[22][0][12] + xor_out[23][0][12] + xor_out[24][0][12];
assign sum_out[5][0][12] = xor_out[25][0][12] + xor_out[26][0][12] + xor_out[27][0][12] + xor_out[28][0][12] + xor_out[29][0][12];
assign sum_out[6][0][12] = xor_out[30][0][12] + xor_out[31][0][12] + xor_out[32][0][12] + xor_out[33][0][12] + xor_out[34][0][12];
assign sum_out[7][0][12] = xor_out[35][0][12] + xor_out[36][0][12] + xor_out[37][0][12] + xor_out[38][0][12] + xor_out[39][0][12];
assign sum_out[8][0][12] = xor_out[40][0][12] + xor_out[41][0][12] + xor_out[42][0][12] + xor_out[43][0][12] + xor_out[44][0][12];
assign sum_out[9][0][12] = xor_out[45][0][12] + xor_out[46][0][12] + xor_out[47][0][12] + xor_out[48][0][12] + xor_out[49][0][12];
assign sum_out[10][0][12] = xor_out[50][0][12] + xor_out[51][0][12] + xor_out[52][0][12] + xor_out[53][0][12] + xor_out[54][0][12];
assign sum_out[11][0][12] = xor_out[55][0][12] + xor_out[56][0][12] + xor_out[57][0][12] + xor_out[58][0][12] + xor_out[59][0][12];
assign sum_out[12][0][12] = xor_out[60][0][12] + xor_out[61][0][12] + xor_out[62][0][12] + xor_out[63][0][12] + xor_out[64][0][12];
assign sum_out[13][0][12] = xor_out[65][0][12] + xor_out[66][0][12] + xor_out[67][0][12] + xor_out[68][0][12] + xor_out[69][0][12];
assign sum_out[14][0][12] = xor_out[70][0][12] + xor_out[71][0][12] + xor_out[72][0][12] + xor_out[73][0][12] + xor_out[74][0][12];
assign sum_out[15][0][12] = xor_out[75][0][12] + xor_out[76][0][12] + xor_out[77][0][12] + xor_out[78][0][12] + xor_out[79][0][12];
assign sum_out[16][0][12] = xor_out[80][0][12] + xor_out[81][0][12] + xor_out[82][0][12] + xor_out[83][0][12] + xor_out[84][0][12];
assign sum_out[17][0][12] = xor_out[85][0][12] + xor_out[86][0][12] + xor_out[87][0][12] + xor_out[88][0][12] + xor_out[89][0][12];
assign sum_out[18][0][12] = xor_out[90][0][12] + xor_out[91][0][12] + xor_out[92][0][12] + xor_out[93][0][12] + xor_out[94][0][12];
assign sum_out[19][0][12] = xor_out[95][0][12] + xor_out[96][0][12] + xor_out[97][0][12] + xor_out[98][0][12] + xor_out[99][0][12];

assign sum_out[0][0][13] = xor_out[0][0][13] + xor_out[1][0][13] + xor_out[2][0][13] + xor_out[3][0][13] + xor_out[4][0][13];
assign sum_out[1][0][13] = xor_out[5][0][13] + xor_out[6][0][13] + xor_out[7][0][13] + xor_out[8][0][13] + xor_out[9][0][13];
assign sum_out[2][0][13] = xor_out[10][0][13] + xor_out[11][0][13] + xor_out[12][0][13] + xor_out[13][0][13] + xor_out[14][0][13];
assign sum_out[3][0][13] = xor_out[15][0][13] + xor_out[16][0][13] + xor_out[17][0][13] + xor_out[18][0][13] + xor_out[19][0][13];
assign sum_out[4][0][13] = xor_out[20][0][13] + xor_out[21][0][13] + xor_out[22][0][13] + xor_out[23][0][13] + xor_out[24][0][13];
assign sum_out[5][0][13] = xor_out[25][0][13] + xor_out[26][0][13] + xor_out[27][0][13] + xor_out[28][0][13] + xor_out[29][0][13];
assign sum_out[6][0][13] = xor_out[30][0][13] + xor_out[31][0][13] + xor_out[32][0][13] + xor_out[33][0][13] + xor_out[34][0][13];
assign sum_out[7][0][13] = xor_out[35][0][13] + xor_out[36][0][13] + xor_out[37][0][13] + xor_out[38][0][13] + xor_out[39][0][13];
assign sum_out[8][0][13] = xor_out[40][0][13] + xor_out[41][0][13] + xor_out[42][0][13] + xor_out[43][0][13] + xor_out[44][0][13];
assign sum_out[9][0][13] = xor_out[45][0][13] + xor_out[46][0][13] + xor_out[47][0][13] + xor_out[48][0][13] + xor_out[49][0][13];
assign sum_out[10][0][13] = xor_out[50][0][13] + xor_out[51][0][13] + xor_out[52][0][13] + xor_out[53][0][13] + xor_out[54][0][13];
assign sum_out[11][0][13] = xor_out[55][0][13] + xor_out[56][0][13] + xor_out[57][0][13] + xor_out[58][0][13] + xor_out[59][0][13];
assign sum_out[12][0][13] = xor_out[60][0][13] + xor_out[61][0][13] + xor_out[62][0][13] + xor_out[63][0][13] + xor_out[64][0][13];
assign sum_out[13][0][13] = xor_out[65][0][13] + xor_out[66][0][13] + xor_out[67][0][13] + xor_out[68][0][13] + xor_out[69][0][13];
assign sum_out[14][0][13] = xor_out[70][0][13] + xor_out[71][0][13] + xor_out[72][0][13] + xor_out[73][0][13] + xor_out[74][0][13];
assign sum_out[15][0][13] = xor_out[75][0][13] + xor_out[76][0][13] + xor_out[77][0][13] + xor_out[78][0][13] + xor_out[79][0][13];
assign sum_out[16][0][13] = xor_out[80][0][13] + xor_out[81][0][13] + xor_out[82][0][13] + xor_out[83][0][13] + xor_out[84][0][13];
assign sum_out[17][0][13] = xor_out[85][0][13] + xor_out[86][0][13] + xor_out[87][0][13] + xor_out[88][0][13] + xor_out[89][0][13];
assign sum_out[18][0][13] = xor_out[90][0][13] + xor_out[91][0][13] + xor_out[92][0][13] + xor_out[93][0][13] + xor_out[94][0][13];
assign sum_out[19][0][13] = xor_out[95][0][13] + xor_out[96][0][13] + xor_out[97][0][13] + xor_out[98][0][13] + xor_out[99][0][13];

assign sum_out[0][0][14] = xor_out[0][0][14] + xor_out[1][0][14] + xor_out[2][0][14] + xor_out[3][0][14] + xor_out[4][0][14];
assign sum_out[1][0][14] = xor_out[5][0][14] + xor_out[6][0][14] + xor_out[7][0][14] + xor_out[8][0][14] + xor_out[9][0][14];
assign sum_out[2][0][14] = xor_out[10][0][14] + xor_out[11][0][14] + xor_out[12][0][14] + xor_out[13][0][14] + xor_out[14][0][14];
assign sum_out[3][0][14] = xor_out[15][0][14] + xor_out[16][0][14] + xor_out[17][0][14] + xor_out[18][0][14] + xor_out[19][0][14];
assign sum_out[4][0][14] = xor_out[20][0][14] + xor_out[21][0][14] + xor_out[22][0][14] + xor_out[23][0][14] + xor_out[24][0][14];
assign sum_out[5][0][14] = xor_out[25][0][14] + xor_out[26][0][14] + xor_out[27][0][14] + xor_out[28][0][14] + xor_out[29][0][14];
assign sum_out[6][0][14] = xor_out[30][0][14] + xor_out[31][0][14] + xor_out[32][0][14] + xor_out[33][0][14] + xor_out[34][0][14];
assign sum_out[7][0][14] = xor_out[35][0][14] + xor_out[36][0][14] + xor_out[37][0][14] + xor_out[38][0][14] + xor_out[39][0][14];
assign sum_out[8][0][14] = xor_out[40][0][14] + xor_out[41][0][14] + xor_out[42][0][14] + xor_out[43][0][14] + xor_out[44][0][14];
assign sum_out[9][0][14] = xor_out[45][0][14] + xor_out[46][0][14] + xor_out[47][0][14] + xor_out[48][0][14] + xor_out[49][0][14];
assign sum_out[10][0][14] = xor_out[50][0][14] + xor_out[51][0][14] + xor_out[52][0][14] + xor_out[53][0][14] + xor_out[54][0][14];
assign sum_out[11][0][14] = xor_out[55][0][14] + xor_out[56][0][14] + xor_out[57][0][14] + xor_out[58][0][14] + xor_out[59][0][14];
assign sum_out[12][0][14] = xor_out[60][0][14] + xor_out[61][0][14] + xor_out[62][0][14] + xor_out[63][0][14] + xor_out[64][0][14];
assign sum_out[13][0][14] = xor_out[65][0][14] + xor_out[66][0][14] + xor_out[67][0][14] + xor_out[68][0][14] + xor_out[69][0][14];
assign sum_out[14][0][14] = xor_out[70][0][14] + xor_out[71][0][14] + xor_out[72][0][14] + xor_out[73][0][14] + xor_out[74][0][14];
assign sum_out[15][0][14] = xor_out[75][0][14] + xor_out[76][0][14] + xor_out[77][0][14] + xor_out[78][0][14] + xor_out[79][0][14];
assign sum_out[16][0][14] = xor_out[80][0][14] + xor_out[81][0][14] + xor_out[82][0][14] + xor_out[83][0][14] + xor_out[84][0][14];
assign sum_out[17][0][14] = xor_out[85][0][14] + xor_out[86][0][14] + xor_out[87][0][14] + xor_out[88][0][14] + xor_out[89][0][14];
assign sum_out[18][0][14] = xor_out[90][0][14] + xor_out[91][0][14] + xor_out[92][0][14] + xor_out[93][0][14] + xor_out[94][0][14];
assign sum_out[19][0][14] = xor_out[95][0][14] + xor_out[96][0][14] + xor_out[97][0][14] + xor_out[98][0][14] + xor_out[99][0][14];

assign sum_out[0][0][15] = xor_out[0][0][15] + xor_out[1][0][15] + xor_out[2][0][15] + xor_out[3][0][15] + xor_out[4][0][15];
assign sum_out[1][0][15] = xor_out[5][0][15] + xor_out[6][0][15] + xor_out[7][0][15] + xor_out[8][0][15] + xor_out[9][0][15];
assign sum_out[2][0][15] = xor_out[10][0][15] + xor_out[11][0][15] + xor_out[12][0][15] + xor_out[13][0][15] + xor_out[14][0][15];
assign sum_out[3][0][15] = xor_out[15][0][15] + xor_out[16][0][15] + xor_out[17][0][15] + xor_out[18][0][15] + xor_out[19][0][15];
assign sum_out[4][0][15] = xor_out[20][0][15] + xor_out[21][0][15] + xor_out[22][0][15] + xor_out[23][0][15] + xor_out[24][0][15];
assign sum_out[5][0][15] = xor_out[25][0][15] + xor_out[26][0][15] + xor_out[27][0][15] + xor_out[28][0][15] + xor_out[29][0][15];
assign sum_out[6][0][15] = xor_out[30][0][15] + xor_out[31][0][15] + xor_out[32][0][15] + xor_out[33][0][15] + xor_out[34][0][15];
assign sum_out[7][0][15] = xor_out[35][0][15] + xor_out[36][0][15] + xor_out[37][0][15] + xor_out[38][0][15] + xor_out[39][0][15];
assign sum_out[8][0][15] = xor_out[40][0][15] + xor_out[41][0][15] + xor_out[42][0][15] + xor_out[43][0][15] + xor_out[44][0][15];
assign sum_out[9][0][15] = xor_out[45][0][15] + xor_out[46][0][15] + xor_out[47][0][15] + xor_out[48][0][15] + xor_out[49][0][15];
assign sum_out[10][0][15] = xor_out[50][0][15] + xor_out[51][0][15] + xor_out[52][0][15] + xor_out[53][0][15] + xor_out[54][0][15];
assign sum_out[11][0][15] = xor_out[55][0][15] + xor_out[56][0][15] + xor_out[57][0][15] + xor_out[58][0][15] + xor_out[59][0][15];
assign sum_out[12][0][15] = xor_out[60][0][15] + xor_out[61][0][15] + xor_out[62][0][15] + xor_out[63][0][15] + xor_out[64][0][15];
assign sum_out[13][0][15] = xor_out[65][0][15] + xor_out[66][0][15] + xor_out[67][0][15] + xor_out[68][0][15] + xor_out[69][0][15];
assign sum_out[14][0][15] = xor_out[70][0][15] + xor_out[71][0][15] + xor_out[72][0][15] + xor_out[73][0][15] + xor_out[74][0][15];
assign sum_out[15][0][15] = xor_out[75][0][15] + xor_out[76][0][15] + xor_out[77][0][15] + xor_out[78][0][15] + xor_out[79][0][15];
assign sum_out[16][0][15] = xor_out[80][0][15] + xor_out[81][0][15] + xor_out[82][0][15] + xor_out[83][0][15] + xor_out[84][0][15];
assign sum_out[17][0][15] = xor_out[85][0][15] + xor_out[86][0][15] + xor_out[87][0][15] + xor_out[88][0][15] + xor_out[89][0][15];
assign sum_out[18][0][15] = xor_out[90][0][15] + xor_out[91][0][15] + xor_out[92][0][15] + xor_out[93][0][15] + xor_out[94][0][15];
assign sum_out[19][0][15] = xor_out[95][0][15] + xor_out[96][0][15] + xor_out[97][0][15] + xor_out[98][0][15] + xor_out[99][0][15];

assign sum_out[0][0][16] = xor_out[0][0][16] + xor_out[1][0][16] + xor_out[2][0][16] + xor_out[3][0][16] + xor_out[4][0][16];
assign sum_out[1][0][16] = xor_out[5][0][16] + xor_out[6][0][16] + xor_out[7][0][16] + xor_out[8][0][16] + xor_out[9][0][16];
assign sum_out[2][0][16] = xor_out[10][0][16] + xor_out[11][0][16] + xor_out[12][0][16] + xor_out[13][0][16] + xor_out[14][0][16];
assign sum_out[3][0][16] = xor_out[15][0][16] + xor_out[16][0][16] + xor_out[17][0][16] + xor_out[18][0][16] + xor_out[19][0][16];
assign sum_out[4][0][16] = xor_out[20][0][16] + xor_out[21][0][16] + xor_out[22][0][16] + xor_out[23][0][16] + xor_out[24][0][16];
assign sum_out[5][0][16] = xor_out[25][0][16] + xor_out[26][0][16] + xor_out[27][0][16] + xor_out[28][0][16] + xor_out[29][0][16];
assign sum_out[6][0][16] = xor_out[30][0][16] + xor_out[31][0][16] + xor_out[32][0][16] + xor_out[33][0][16] + xor_out[34][0][16];
assign sum_out[7][0][16] = xor_out[35][0][16] + xor_out[36][0][16] + xor_out[37][0][16] + xor_out[38][0][16] + xor_out[39][0][16];
assign sum_out[8][0][16] = xor_out[40][0][16] + xor_out[41][0][16] + xor_out[42][0][16] + xor_out[43][0][16] + xor_out[44][0][16];
assign sum_out[9][0][16] = xor_out[45][0][16] + xor_out[46][0][16] + xor_out[47][0][16] + xor_out[48][0][16] + xor_out[49][0][16];
assign sum_out[10][0][16] = xor_out[50][0][16] + xor_out[51][0][16] + xor_out[52][0][16] + xor_out[53][0][16] + xor_out[54][0][16];
assign sum_out[11][0][16] = xor_out[55][0][16] + xor_out[56][0][16] + xor_out[57][0][16] + xor_out[58][0][16] + xor_out[59][0][16];
assign sum_out[12][0][16] = xor_out[60][0][16] + xor_out[61][0][16] + xor_out[62][0][16] + xor_out[63][0][16] + xor_out[64][0][16];
assign sum_out[13][0][16] = xor_out[65][0][16] + xor_out[66][0][16] + xor_out[67][0][16] + xor_out[68][0][16] + xor_out[69][0][16];
assign sum_out[14][0][16] = xor_out[70][0][16] + xor_out[71][0][16] + xor_out[72][0][16] + xor_out[73][0][16] + xor_out[74][0][16];
assign sum_out[15][0][16] = xor_out[75][0][16] + xor_out[76][0][16] + xor_out[77][0][16] + xor_out[78][0][16] + xor_out[79][0][16];
assign sum_out[16][0][16] = xor_out[80][0][16] + xor_out[81][0][16] + xor_out[82][0][16] + xor_out[83][0][16] + xor_out[84][0][16];
assign sum_out[17][0][16] = xor_out[85][0][16] + xor_out[86][0][16] + xor_out[87][0][16] + xor_out[88][0][16] + xor_out[89][0][16];
assign sum_out[18][0][16] = xor_out[90][0][16] + xor_out[91][0][16] + xor_out[92][0][16] + xor_out[93][0][16] + xor_out[94][0][16];
assign sum_out[19][0][16] = xor_out[95][0][16] + xor_out[96][0][16] + xor_out[97][0][16] + xor_out[98][0][16] + xor_out[99][0][16];

assign sum_out[0][0][17] = xor_out[0][0][17] + xor_out[1][0][17] + xor_out[2][0][17] + xor_out[3][0][17] + xor_out[4][0][17];
assign sum_out[1][0][17] = xor_out[5][0][17] + xor_out[6][0][17] + xor_out[7][0][17] + xor_out[8][0][17] + xor_out[9][0][17];
assign sum_out[2][0][17] = xor_out[10][0][17] + xor_out[11][0][17] + xor_out[12][0][17] + xor_out[13][0][17] + xor_out[14][0][17];
assign sum_out[3][0][17] = xor_out[15][0][17] + xor_out[16][0][17] + xor_out[17][0][17] + xor_out[18][0][17] + xor_out[19][0][17];
assign sum_out[4][0][17] = xor_out[20][0][17] + xor_out[21][0][17] + xor_out[22][0][17] + xor_out[23][0][17] + xor_out[24][0][17];
assign sum_out[5][0][17] = xor_out[25][0][17] + xor_out[26][0][17] + xor_out[27][0][17] + xor_out[28][0][17] + xor_out[29][0][17];
assign sum_out[6][0][17] = xor_out[30][0][17] + xor_out[31][0][17] + xor_out[32][0][17] + xor_out[33][0][17] + xor_out[34][0][17];
assign sum_out[7][0][17] = xor_out[35][0][17] + xor_out[36][0][17] + xor_out[37][0][17] + xor_out[38][0][17] + xor_out[39][0][17];
assign sum_out[8][0][17] = xor_out[40][0][17] + xor_out[41][0][17] + xor_out[42][0][17] + xor_out[43][0][17] + xor_out[44][0][17];
assign sum_out[9][0][17] = xor_out[45][0][17] + xor_out[46][0][17] + xor_out[47][0][17] + xor_out[48][0][17] + xor_out[49][0][17];
assign sum_out[10][0][17] = xor_out[50][0][17] + xor_out[51][0][17] + xor_out[52][0][17] + xor_out[53][0][17] + xor_out[54][0][17];
assign sum_out[11][0][17] = xor_out[55][0][17] + xor_out[56][0][17] + xor_out[57][0][17] + xor_out[58][0][17] + xor_out[59][0][17];
assign sum_out[12][0][17] = xor_out[60][0][17] + xor_out[61][0][17] + xor_out[62][0][17] + xor_out[63][0][17] + xor_out[64][0][17];
assign sum_out[13][0][17] = xor_out[65][0][17] + xor_out[66][0][17] + xor_out[67][0][17] + xor_out[68][0][17] + xor_out[69][0][17];
assign sum_out[14][0][17] = xor_out[70][0][17] + xor_out[71][0][17] + xor_out[72][0][17] + xor_out[73][0][17] + xor_out[74][0][17];
assign sum_out[15][0][17] = xor_out[75][0][17] + xor_out[76][0][17] + xor_out[77][0][17] + xor_out[78][0][17] + xor_out[79][0][17];
assign sum_out[16][0][17] = xor_out[80][0][17] + xor_out[81][0][17] + xor_out[82][0][17] + xor_out[83][0][17] + xor_out[84][0][17];
assign sum_out[17][0][17] = xor_out[85][0][17] + xor_out[86][0][17] + xor_out[87][0][17] + xor_out[88][0][17] + xor_out[89][0][17];
assign sum_out[18][0][17] = xor_out[90][0][17] + xor_out[91][0][17] + xor_out[92][0][17] + xor_out[93][0][17] + xor_out[94][0][17];
assign sum_out[19][0][17] = xor_out[95][0][17] + xor_out[96][0][17] + xor_out[97][0][17] + xor_out[98][0][17] + xor_out[99][0][17];

assign sum_out[0][0][18] = xor_out[0][0][18] + xor_out[1][0][18] + xor_out[2][0][18] + xor_out[3][0][18] + xor_out[4][0][18];
assign sum_out[1][0][18] = xor_out[5][0][18] + xor_out[6][0][18] + xor_out[7][0][18] + xor_out[8][0][18] + xor_out[9][0][18];
assign sum_out[2][0][18] = xor_out[10][0][18] + xor_out[11][0][18] + xor_out[12][0][18] + xor_out[13][0][18] + xor_out[14][0][18];
assign sum_out[3][0][18] = xor_out[15][0][18] + xor_out[16][0][18] + xor_out[17][0][18] + xor_out[18][0][18] + xor_out[19][0][18];
assign sum_out[4][0][18] = xor_out[20][0][18] + xor_out[21][0][18] + xor_out[22][0][18] + xor_out[23][0][18] + xor_out[24][0][18];
assign sum_out[5][0][18] = xor_out[25][0][18] + xor_out[26][0][18] + xor_out[27][0][18] + xor_out[28][0][18] + xor_out[29][0][18];
assign sum_out[6][0][18] = xor_out[30][0][18] + xor_out[31][0][18] + xor_out[32][0][18] + xor_out[33][0][18] + xor_out[34][0][18];
assign sum_out[7][0][18] = xor_out[35][0][18] + xor_out[36][0][18] + xor_out[37][0][18] + xor_out[38][0][18] + xor_out[39][0][18];
assign sum_out[8][0][18] = xor_out[40][0][18] + xor_out[41][0][18] + xor_out[42][0][18] + xor_out[43][0][18] + xor_out[44][0][18];
assign sum_out[9][0][18] = xor_out[45][0][18] + xor_out[46][0][18] + xor_out[47][0][18] + xor_out[48][0][18] + xor_out[49][0][18];
assign sum_out[10][0][18] = xor_out[50][0][18] + xor_out[51][0][18] + xor_out[52][0][18] + xor_out[53][0][18] + xor_out[54][0][18];
assign sum_out[11][0][18] = xor_out[55][0][18] + xor_out[56][0][18] + xor_out[57][0][18] + xor_out[58][0][18] + xor_out[59][0][18];
assign sum_out[12][0][18] = xor_out[60][0][18] + xor_out[61][0][18] + xor_out[62][0][18] + xor_out[63][0][18] + xor_out[64][0][18];
assign sum_out[13][0][18] = xor_out[65][0][18] + xor_out[66][0][18] + xor_out[67][0][18] + xor_out[68][0][18] + xor_out[69][0][18];
assign sum_out[14][0][18] = xor_out[70][0][18] + xor_out[71][0][18] + xor_out[72][0][18] + xor_out[73][0][18] + xor_out[74][0][18];
assign sum_out[15][0][18] = xor_out[75][0][18] + xor_out[76][0][18] + xor_out[77][0][18] + xor_out[78][0][18] + xor_out[79][0][18];
assign sum_out[16][0][18] = xor_out[80][0][18] + xor_out[81][0][18] + xor_out[82][0][18] + xor_out[83][0][18] + xor_out[84][0][18];
assign sum_out[17][0][18] = xor_out[85][0][18] + xor_out[86][0][18] + xor_out[87][0][18] + xor_out[88][0][18] + xor_out[89][0][18];
assign sum_out[18][0][18] = xor_out[90][0][18] + xor_out[91][0][18] + xor_out[92][0][18] + xor_out[93][0][18] + xor_out[94][0][18];
assign sum_out[19][0][18] = xor_out[95][0][18] + xor_out[96][0][18] + xor_out[97][0][18] + xor_out[98][0][18] + xor_out[99][0][18];

assign sum_out[0][0][19] = xor_out[0][0][19] + xor_out[1][0][19] + xor_out[2][0][19] + xor_out[3][0][19] + xor_out[4][0][19];
assign sum_out[1][0][19] = xor_out[5][0][19] + xor_out[6][0][19] + xor_out[7][0][19] + xor_out[8][0][19] + xor_out[9][0][19];
assign sum_out[2][0][19] = xor_out[10][0][19] + xor_out[11][0][19] + xor_out[12][0][19] + xor_out[13][0][19] + xor_out[14][0][19];
assign sum_out[3][0][19] = xor_out[15][0][19] + xor_out[16][0][19] + xor_out[17][0][19] + xor_out[18][0][19] + xor_out[19][0][19];
assign sum_out[4][0][19] = xor_out[20][0][19] + xor_out[21][0][19] + xor_out[22][0][19] + xor_out[23][0][19] + xor_out[24][0][19];
assign sum_out[5][0][19] = xor_out[25][0][19] + xor_out[26][0][19] + xor_out[27][0][19] + xor_out[28][0][19] + xor_out[29][0][19];
assign sum_out[6][0][19] = xor_out[30][0][19] + xor_out[31][0][19] + xor_out[32][0][19] + xor_out[33][0][19] + xor_out[34][0][19];
assign sum_out[7][0][19] = xor_out[35][0][19] + xor_out[36][0][19] + xor_out[37][0][19] + xor_out[38][0][19] + xor_out[39][0][19];
assign sum_out[8][0][19] = xor_out[40][0][19] + xor_out[41][0][19] + xor_out[42][0][19] + xor_out[43][0][19] + xor_out[44][0][19];
assign sum_out[9][0][19] = xor_out[45][0][19] + xor_out[46][0][19] + xor_out[47][0][19] + xor_out[48][0][19] + xor_out[49][0][19];
assign sum_out[10][0][19] = xor_out[50][0][19] + xor_out[51][0][19] + xor_out[52][0][19] + xor_out[53][0][19] + xor_out[54][0][19];
assign sum_out[11][0][19] = xor_out[55][0][19] + xor_out[56][0][19] + xor_out[57][0][19] + xor_out[58][0][19] + xor_out[59][0][19];
assign sum_out[12][0][19] = xor_out[60][0][19] + xor_out[61][0][19] + xor_out[62][0][19] + xor_out[63][0][19] + xor_out[64][0][19];
assign sum_out[13][0][19] = xor_out[65][0][19] + xor_out[66][0][19] + xor_out[67][0][19] + xor_out[68][0][19] + xor_out[69][0][19];
assign sum_out[14][0][19] = xor_out[70][0][19] + xor_out[71][0][19] + xor_out[72][0][19] + xor_out[73][0][19] + xor_out[74][0][19];
assign sum_out[15][0][19] = xor_out[75][0][19] + xor_out[76][0][19] + xor_out[77][0][19] + xor_out[78][0][19] + xor_out[79][0][19];
assign sum_out[16][0][19] = xor_out[80][0][19] + xor_out[81][0][19] + xor_out[82][0][19] + xor_out[83][0][19] + xor_out[84][0][19];
assign sum_out[17][0][19] = xor_out[85][0][19] + xor_out[86][0][19] + xor_out[87][0][19] + xor_out[88][0][19] + xor_out[89][0][19];
assign sum_out[18][0][19] = xor_out[90][0][19] + xor_out[91][0][19] + xor_out[92][0][19] + xor_out[93][0][19] + xor_out[94][0][19];
assign sum_out[19][0][19] = xor_out[95][0][19] + xor_out[96][0][19] + xor_out[97][0][19] + xor_out[98][0][19] + xor_out[99][0][19];

assign sum_out[0][0][20] = xor_out[0][0][20] + xor_out[1][0][20] + xor_out[2][0][20] + xor_out[3][0][20] + xor_out[4][0][20];
assign sum_out[1][0][20] = xor_out[5][0][20] + xor_out[6][0][20] + xor_out[7][0][20] + xor_out[8][0][20] + xor_out[9][0][20];
assign sum_out[2][0][20] = xor_out[10][0][20] + xor_out[11][0][20] + xor_out[12][0][20] + xor_out[13][0][20] + xor_out[14][0][20];
assign sum_out[3][0][20] = xor_out[15][0][20] + xor_out[16][0][20] + xor_out[17][0][20] + xor_out[18][0][20] + xor_out[19][0][20];
assign sum_out[4][0][20] = xor_out[20][0][20] + xor_out[21][0][20] + xor_out[22][0][20] + xor_out[23][0][20] + xor_out[24][0][20];
assign sum_out[5][0][20] = xor_out[25][0][20] + xor_out[26][0][20] + xor_out[27][0][20] + xor_out[28][0][20] + xor_out[29][0][20];
assign sum_out[6][0][20] = xor_out[30][0][20] + xor_out[31][0][20] + xor_out[32][0][20] + xor_out[33][0][20] + xor_out[34][0][20];
assign sum_out[7][0][20] = xor_out[35][0][20] + xor_out[36][0][20] + xor_out[37][0][20] + xor_out[38][0][20] + xor_out[39][0][20];
assign sum_out[8][0][20] = xor_out[40][0][20] + xor_out[41][0][20] + xor_out[42][0][20] + xor_out[43][0][20] + xor_out[44][0][20];
assign sum_out[9][0][20] = xor_out[45][0][20] + xor_out[46][0][20] + xor_out[47][0][20] + xor_out[48][0][20] + xor_out[49][0][20];
assign sum_out[10][0][20] = xor_out[50][0][20] + xor_out[51][0][20] + xor_out[52][0][20] + xor_out[53][0][20] + xor_out[54][0][20];
assign sum_out[11][0][20] = xor_out[55][0][20] + xor_out[56][0][20] + xor_out[57][0][20] + xor_out[58][0][20] + xor_out[59][0][20];
assign sum_out[12][0][20] = xor_out[60][0][20] + xor_out[61][0][20] + xor_out[62][0][20] + xor_out[63][0][20] + xor_out[64][0][20];
assign sum_out[13][0][20] = xor_out[65][0][20] + xor_out[66][0][20] + xor_out[67][0][20] + xor_out[68][0][20] + xor_out[69][0][20];
assign sum_out[14][0][20] = xor_out[70][0][20] + xor_out[71][0][20] + xor_out[72][0][20] + xor_out[73][0][20] + xor_out[74][0][20];
assign sum_out[15][0][20] = xor_out[75][0][20] + xor_out[76][0][20] + xor_out[77][0][20] + xor_out[78][0][20] + xor_out[79][0][20];
assign sum_out[16][0][20] = xor_out[80][0][20] + xor_out[81][0][20] + xor_out[82][0][20] + xor_out[83][0][20] + xor_out[84][0][20];
assign sum_out[17][0][20] = xor_out[85][0][20] + xor_out[86][0][20] + xor_out[87][0][20] + xor_out[88][0][20] + xor_out[89][0][20];
assign sum_out[18][0][20] = xor_out[90][0][20] + xor_out[91][0][20] + xor_out[92][0][20] + xor_out[93][0][20] + xor_out[94][0][20];
assign sum_out[19][0][20] = xor_out[95][0][20] + xor_out[96][0][20] + xor_out[97][0][20] + xor_out[98][0][20] + xor_out[99][0][20];

assign sum_out[0][0][21] = xor_out[0][0][21] + xor_out[1][0][21] + xor_out[2][0][21] + xor_out[3][0][21] + xor_out[4][0][21];
assign sum_out[1][0][21] = xor_out[5][0][21] + xor_out[6][0][21] + xor_out[7][0][21] + xor_out[8][0][21] + xor_out[9][0][21];
assign sum_out[2][0][21] = xor_out[10][0][21] + xor_out[11][0][21] + xor_out[12][0][21] + xor_out[13][0][21] + xor_out[14][0][21];
assign sum_out[3][0][21] = xor_out[15][0][21] + xor_out[16][0][21] + xor_out[17][0][21] + xor_out[18][0][21] + xor_out[19][0][21];
assign sum_out[4][0][21] = xor_out[20][0][21] + xor_out[21][0][21] + xor_out[22][0][21] + xor_out[23][0][21] + xor_out[24][0][21];
assign sum_out[5][0][21] = xor_out[25][0][21] + xor_out[26][0][21] + xor_out[27][0][21] + xor_out[28][0][21] + xor_out[29][0][21];
assign sum_out[6][0][21] = xor_out[30][0][21] + xor_out[31][0][21] + xor_out[32][0][21] + xor_out[33][0][21] + xor_out[34][0][21];
assign sum_out[7][0][21] = xor_out[35][0][21] + xor_out[36][0][21] + xor_out[37][0][21] + xor_out[38][0][21] + xor_out[39][0][21];
assign sum_out[8][0][21] = xor_out[40][0][21] + xor_out[41][0][21] + xor_out[42][0][21] + xor_out[43][0][21] + xor_out[44][0][21];
assign sum_out[9][0][21] = xor_out[45][0][21] + xor_out[46][0][21] + xor_out[47][0][21] + xor_out[48][0][21] + xor_out[49][0][21];
assign sum_out[10][0][21] = xor_out[50][0][21] + xor_out[51][0][21] + xor_out[52][0][21] + xor_out[53][0][21] + xor_out[54][0][21];
assign sum_out[11][0][21] = xor_out[55][0][21] + xor_out[56][0][21] + xor_out[57][0][21] + xor_out[58][0][21] + xor_out[59][0][21];
assign sum_out[12][0][21] = xor_out[60][0][21] + xor_out[61][0][21] + xor_out[62][0][21] + xor_out[63][0][21] + xor_out[64][0][21];
assign sum_out[13][0][21] = xor_out[65][0][21] + xor_out[66][0][21] + xor_out[67][0][21] + xor_out[68][0][21] + xor_out[69][0][21];
assign sum_out[14][0][21] = xor_out[70][0][21] + xor_out[71][0][21] + xor_out[72][0][21] + xor_out[73][0][21] + xor_out[74][0][21];
assign sum_out[15][0][21] = xor_out[75][0][21] + xor_out[76][0][21] + xor_out[77][0][21] + xor_out[78][0][21] + xor_out[79][0][21];
assign sum_out[16][0][21] = xor_out[80][0][21] + xor_out[81][0][21] + xor_out[82][0][21] + xor_out[83][0][21] + xor_out[84][0][21];
assign sum_out[17][0][21] = xor_out[85][0][21] + xor_out[86][0][21] + xor_out[87][0][21] + xor_out[88][0][21] + xor_out[89][0][21];
assign sum_out[18][0][21] = xor_out[90][0][21] + xor_out[91][0][21] + xor_out[92][0][21] + xor_out[93][0][21] + xor_out[94][0][21];
assign sum_out[19][0][21] = xor_out[95][0][21] + xor_out[96][0][21] + xor_out[97][0][21] + xor_out[98][0][21] + xor_out[99][0][21];

assign sum_out[0][0][22] = xor_out[0][0][22] + xor_out[1][0][22] + xor_out[2][0][22] + xor_out[3][0][22] + xor_out[4][0][22];
assign sum_out[1][0][22] = xor_out[5][0][22] + xor_out[6][0][22] + xor_out[7][0][22] + xor_out[8][0][22] + xor_out[9][0][22];
assign sum_out[2][0][22] = xor_out[10][0][22] + xor_out[11][0][22] + xor_out[12][0][22] + xor_out[13][0][22] + xor_out[14][0][22];
assign sum_out[3][0][22] = xor_out[15][0][22] + xor_out[16][0][22] + xor_out[17][0][22] + xor_out[18][0][22] + xor_out[19][0][22];
assign sum_out[4][0][22] = xor_out[20][0][22] + xor_out[21][0][22] + xor_out[22][0][22] + xor_out[23][0][22] + xor_out[24][0][22];
assign sum_out[5][0][22] = xor_out[25][0][22] + xor_out[26][0][22] + xor_out[27][0][22] + xor_out[28][0][22] + xor_out[29][0][22];
assign sum_out[6][0][22] = xor_out[30][0][22] + xor_out[31][0][22] + xor_out[32][0][22] + xor_out[33][0][22] + xor_out[34][0][22];
assign sum_out[7][0][22] = xor_out[35][0][22] + xor_out[36][0][22] + xor_out[37][0][22] + xor_out[38][0][22] + xor_out[39][0][22];
assign sum_out[8][0][22] = xor_out[40][0][22] + xor_out[41][0][22] + xor_out[42][0][22] + xor_out[43][0][22] + xor_out[44][0][22];
assign sum_out[9][0][22] = xor_out[45][0][22] + xor_out[46][0][22] + xor_out[47][0][22] + xor_out[48][0][22] + xor_out[49][0][22];
assign sum_out[10][0][22] = xor_out[50][0][22] + xor_out[51][0][22] + xor_out[52][0][22] + xor_out[53][0][22] + xor_out[54][0][22];
assign sum_out[11][0][22] = xor_out[55][0][22] + xor_out[56][0][22] + xor_out[57][0][22] + xor_out[58][0][22] + xor_out[59][0][22];
assign sum_out[12][0][22] = xor_out[60][0][22] + xor_out[61][0][22] + xor_out[62][0][22] + xor_out[63][0][22] + xor_out[64][0][22];
assign sum_out[13][0][22] = xor_out[65][0][22] + xor_out[66][0][22] + xor_out[67][0][22] + xor_out[68][0][22] + xor_out[69][0][22];
assign sum_out[14][0][22] = xor_out[70][0][22] + xor_out[71][0][22] + xor_out[72][0][22] + xor_out[73][0][22] + xor_out[74][0][22];
assign sum_out[15][0][22] = xor_out[75][0][22] + xor_out[76][0][22] + xor_out[77][0][22] + xor_out[78][0][22] + xor_out[79][0][22];
assign sum_out[16][0][22] = xor_out[80][0][22] + xor_out[81][0][22] + xor_out[82][0][22] + xor_out[83][0][22] + xor_out[84][0][22];
assign sum_out[17][0][22] = xor_out[85][0][22] + xor_out[86][0][22] + xor_out[87][0][22] + xor_out[88][0][22] + xor_out[89][0][22];
assign sum_out[18][0][22] = xor_out[90][0][22] + xor_out[91][0][22] + xor_out[92][0][22] + xor_out[93][0][22] + xor_out[94][0][22];
assign sum_out[19][0][22] = xor_out[95][0][22] + xor_out[96][0][22] + xor_out[97][0][22] + xor_out[98][0][22] + xor_out[99][0][22];

assign sum_out[0][0][23] = xor_out[0][0][23] + xor_out[1][0][23] + xor_out[2][0][23] + xor_out[3][0][23] + xor_out[4][0][23];
assign sum_out[1][0][23] = xor_out[5][0][23] + xor_out[6][0][23] + xor_out[7][0][23] + xor_out[8][0][23] + xor_out[9][0][23];
assign sum_out[2][0][23] = xor_out[10][0][23] + xor_out[11][0][23] + xor_out[12][0][23] + xor_out[13][0][23] + xor_out[14][0][23];
assign sum_out[3][0][23] = xor_out[15][0][23] + xor_out[16][0][23] + xor_out[17][0][23] + xor_out[18][0][23] + xor_out[19][0][23];
assign sum_out[4][0][23] = xor_out[20][0][23] + xor_out[21][0][23] + xor_out[22][0][23] + xor_out[23][0][23] + xor_out[24][0][23];
assign sum_out[5][0][23] = xor_out[25][0][23] + xor_out[26][0][23] + xor_out[27][0][23] + xor_out[28][0][23] + xor_out[29][0][23];
assign sum_out[6][0][23] = xor_out[30][0][23] + xor_out[31][0][23] + xor_out[32][0][23] + xor_out[33][0][23] + xor_out[34][0][23];
assign sum_out[7][0][23] = xor_out[35][0][23] + xor_out[36][0][23] + xor_out[37][0][23] + xor_out[38][0][23] + xor_out[39][0][23];
assign sum_out[8][0][23] = xor_out[40][0][23] + xor_out[41][0][23] + xor_out[42][0][23] + xor_out[43][0][23] + xor_out[44][0][23];
assign sum_out[9][0][23] = xor_out[45][0][23] + xor_out[46][0][23] + xor_out[47][0][23] + xor_out[48][0][23] + xor_out[49][0][23];
assign sum_out[10][0][23] = xor_out[50][0][23] + xor_out[51][0][23] + xor_out[52][0][23] + xor_out[53][0][23] + xor_out[54][0][23];
assign sum_out[11][0][23] = xor_out[55][0][23] + xor_out[56][0][23] + xor_out[57][0][23] + xor_out[58][0][23] + xor_out[59][0][23];
assign sum_out[12][0][23] = xor_out[60][0][23] + xor_out[61][0][23] + xor_out[62][0][23] + xor_out[63][0][23] + xor_out[64][0][23];
assign sum_out[13][0][23] = xor_out[65][0][23] + xor_out[66][0][23] + xor_out[67][0][23] + xor_out[68][0][23] + xor_out[69][0][23];
assign sum_out[14][0][23] = xor_out[70][0][23] + xor_out[71][0][23] + xor_out[72][0][23] + xor_out[73][0][23] + xor_out[74][0][23];
assign sum_out[15][0][23] = xor_out[75][0][23] + xor_out[76][0][23] + xor_out[77][0][23] + xor_out[78][0][23] + xor_out[79][0][23];
assign sum_out[16][0][23] = xor_out[80][0][23] + xor_out[81][0][23] + xor_out[82][0][23] + xor_out[83][0][23] + xor_out[84][0][23];
assign sum_out[17][0][23] = xor_out[85][0][23] + xor_out[86][0][23] + xor_out[87][0][23] + xor_out[88][0][23] + xor_out[89][0][23];
assign sum_out[18][0][23] = xor_out[90][0][23] + xor_out[91][0][23] + xor_out[92][0][23] + xor_out[93][0][23] + xor_out[94][0][23];
assign sum_out[19][0][23] = xor_out[95][0][23] + xor_out[96][0][23] + xor_out[97][0][23] + xor_out[98][0][23] + xor_out[99][0][23];

assign sum_out[0][1][0] = xor_out[0][1][0] + xor_out[1][1][0] + xor_out[2][1][0] + xor_out[3][1][0] + xor_out[4][1][0];
assign sum_out[1][1][0] = xor_out[5][1][0] + xor_out[6][1][0] + xor_out[7][1][0] + xor_out[8][1][0] + xor_out[9][1][0];
assign sum_out[2][1][0] = xor_out[10][1][0] + xor_out[11][1][0] + xor_out[12][1][0] + xor_out[13][1][0] + xor_out[14][1][0];
assign sum_out[3][1][0] = xor_out[15][1][0] + xor_out[16][1][0] + xor_out[17][1][0] + xor_out[18][1][0] + xor_out[19][1][0];
assign sum_out[4][1][0] = xor_out[20][1][0] + xor_out[21][1][0] + xor_out[22][1][0] + xor_out[23][1][0] + xor_out[24][1][0];
assign sum_out[5][1][0] = xor_out[25][1][0] + xor_out[26][1][0] + xor_out[27][1][0] + xor_out[28][1][0] + xor_out[29][1][0];
assign sum_out[6][1][0] = xor_out[30][1][0] + xor_out[31][1][0] + xor_out[32][1][0] + xor_out[33][1][0] + xor_out[34][1][0];
assign sum_out[7][1][0] = xor_out[35][1][0] + xor_out[36][1][0] + xor_out[37][1][0] + xor_out[38][1][0] + xor_out[39][1][0];
assign sum_out[8][1][0] = xor_out[40][1][0] + xor_out[41][1][0] + xor_out[42][1][0] + xor_out[43][1][0] + xor_out[44][1][0];
assign sum_out[9][1][0] = xor_out[45][1][0] + xor_out[46][1][0] + xor_out[47][1][0] + xor_out[48][1][0] + xor_out[49][1][0];
assign sum_out[10][1][0] = xor_out[50][1][0] + xor_out[51][1][0] + xor_out[52][1][0] + xor_out[53][1][0] + xor_out[54][1][0];
assign sum_out[11][1][0] = xor_out[55][1][0] + xor_out[56][1][0] + xor_out[57][1][0] + xor_out[58][1][0] + xor_out[59][1][0];
assign sum_out[12][1][0] = xor_out[60][1][0] + xor_out[61][1][0] + xor_out[62][1][0] + xor_out[63][1][0] + xor_out[64][1][0];
assign sum_out[13][1][0] = xor_out[65][1][0] + xor_out[66][1][0] + xor_out[67][1][0] + xor_out[68][1][0] + xor_out[69][1][0];
assign sum_out[14][1][0] = xor_out[70][1][0] + xor_out[71][1][0] + xor_out[72][1][0] + xor_out[73][1][0] + xor_out[74][1][0];
assign sum_out[15][1][0] = xor_out[75][1][0] + xor_out[76][1][0] + xor_out[77][1][0] + xor_out[78][1][0] + xor_out[79][1][0];
assign sum_out[16][1][0] = xor_out[80][1][0] + xor_out[81][1][0] + xor_out[82][1][0] + xor_out[83][1][0] + xor_out[84][1][0];
assign sum_out[17][1][0] = xor_out[85][1][0] + xor_out[86][1][0] + xor_out[87][1][0] + xor_out[88][1][0] + xor_out[89][1][0];
assign sum_out[18][1][0] = xor_out[90][1][0] + xor_out[91][1][0] + xor_out[92][1][0] + xor_out[93][1][0] + xor_out[94][1][0];
assign sum_out[19][1][0] = xor_out[95][1][0] + xor_out[96][1][0] + xor_out[97][1][0] + xor_out[98][1][0] + xor_out[99][1][0];

assign sum_out[0][1][1] = xor_out[0][1][1] + xor_out[1][1][1] + xor_out[2][1][1] + xor_out[3][1][1] + xor_out[4][1][1];
assign sum_out[1][1][1] = xor_out[5][1][1] + xor_out[6][1][1] + xor_out[7][1][1] + xor_out[8][1][1] + xor_out[9][1][1];
assign sum_out[2][1][1] = xor_out[10][1][1] + xor_out[11][1][1] + xor_out[12][1][1] + xor_out[13][1][1] + xor_out[14][1][1];
assign sum_out[3][1][1] = xor_out[15][1][1] + xor_out[16][1][1] + xor_out[17][1][1] + xor_out[18][1][1] + xor_out[19][1][1];
assign sum_out[4][1][1] = xor_out[20][1][1] + xor_out[21][1][1] + xor_out[22][1][1] + xor_out[23][1][1] + xor_out[24][1][1];
assign sum_out[5][1][1] = xor_out[25][1][1] + xor_out[26][1][1] + xor_out[27][1][1] + xor_out[28][1][1] + xor_out[29][1][1];
assign sum_out[6][1][1] = xor_out[30][1][1] + xor_out[31][1][1] + xor_out[32][1][1] + xor_out[33][1][1] + xor_out[34][1][1];
assign sum_out[7][1][1] = xor_out[35][1][1] + xor_out[36][1][1] + xor_out[37][1][1] + xor_out[38][1][1] + xor_out[39][1][1];
assign sum_out[8][1][1] = xor_out[40][1][1] + xor_out[41][1][1] + xor_out[42][1][1] + xor_out[43][1][1] + xor_out[44][1][1];
assign sum_out[9][1][1] = xor_out[45][1][1] + xor_out[46][1][1] + xor_out[47][1][1] + xor_out[48][1][1] + xor_out[49][1][1];
assign sum_out[10][1][1] = xor_out[50][1][1] + xor_out[51][1][1] + xor_out[52][1][1] + xor_out[53][1][1] + xor_out[54][1][1];
assign sum_out[11][1][1] = xor_out[55][1][1] + xor_out[56][1][1] + xor_out[57][1][1] + xor_out[58][1][1] + xor_out[59][1][1];
assign sum_out[12][1][1] = xor_out[60][1][1] + xor_out[61][1][1] + xor_out[62][1][1] + xor_out[63][1][1] + xor_out[64][1][1];
assign sum_out[13][1][1] = xor_out[65][1][1] + xor_out[66][1][1] + xor_out[67][1][1] + xor_out[68][1][1] + xor_out[69][1][1];
assign sum_out[14][1][1] = xor_out[70][1][1] + xor_out[71][1][1] + xor_out[72][1][1] + xor_out[73][1][1] + xor_out[74][1][1];
assign sum_out[15][1][1] = xor_out[75][1][1] + xor_out[76][1][1] + xor_out[77][1][1] + xor_out[78][1][1] + xor_out[79][1][1];
assign sum_out[16][1][1] = xor_out[80][1][1] + xor_out[81][1][1] + xor_out[82][1][1] + xor_out[83][1][1] + xor_out[84][1][1];
assign sum_out[17][1][1] = xor_out[85][1][1] + xor_out[86][1][1] + xor_out[87][1][1] + xor_out[88][1][1] + xor_out[89][1][1];
assign sum_out[18][1][1] = xor_out[90][1][1] + xor_out[91][1][1] + xor_out[92][1][1] + xor_out[93][1][1] + xor_out[94][1][1];
assign sum_out[19][1][1] = xor_out[95][1][1] + xor_out[96][1][1] + xor_out[97][1][1] + xor_out[98][1][1] + xor_out[99][1][1];

assign sum_out[0][1][2] = xor_out[0][1][2] + xor_out[1][1][2] + xor_out[2][1][2] + xor_out[3][1][2] + xor_out[4][1][2];
assign sum_out[1][1][2] = xor_out[5][1][2] + xor_out[6][1][2] + xor_out[7][1][2] + xor_out[8][1][2] + xor_out[9][1][2];
assign sum_out[2][1][2] = xor_out[10][1][2] + xor_out[11][1][2] + xor_out[12][1][2] + xor_out[13][1][2] + xor_out[14][1][2];
assign sum_out[3][1][2] = xor_out[15][1][2] + xor_out[16][1][2] + xor_out[17][1][2] + xor_out[18][1][2] + xor_out[19][1][2];
assign sum_out[4][1][2] = xor_out[20][1][2] + xor_out[21][1][2] + xor_out[22][1][2] + xor_out[23][1][2] + xor_out[24][1][2];
assign sum_out[5][1][2] = xor_out[25][1][2] + xor_out[26][1][2] + xor_out[27][1][2] + xor_out[28][1][2] + xor_out[29][1][2];
assign sum_out[6][1][2] = xor_out[30][1][2] + xor_out[31][1][2] + xor_out[32][1][2] + xor_out[33][1][2] + xor_out[34][1][2];
assign sum_out[7][1][2] = xor_out[35][1][2] + xor_out[36][1][2] + xor_out[37][1][2] + xor_out[38][1][2] + xor_out[39][1][2];
assign sum_out[8][1][2] = xor_out[40][1][2] + xor_out[41][1][2] + xor_out[42][1][2] + xor_out[43][1][2] + xor_out[44][1][2];
assign sum_out[9][1][2] = xor_out[45][1][2] + xor_out[46][1][2] + xor_out[47][1][2] + xor_out[48][1][2] + xor_out[49][1][2];
assign sum_out[10][1][2] = xor_out[50][1][2] + xor_out[51][1][2] + xor_out[52][1][2] + xor_out[53][1][2] + xor_out[54][1][2];
assign sum_out[11][1][2] = xor_out[55][1][2] + xor_out[56][1][2] + xor_out[57][1][2] + xor_out[58][1][2] + xor_out[59][1][2];
assign sum_out[12][1][2] = xor_out[60][1][2] + xor_out[61][1][2] + xor_out[62][1][2] + xor_out[63][1][2] + xor_out[64][1][2];
assign sum_out[13][1][2] = xor_out[65][1][2] + xor_out[66][1][2] + xor_out[67][1][2] + xor_out[68][1][2] + xor_out[69][1][2];
assign sum_out[14][1][2] = xor_out[70][1][2] + xor_out[71][1][2] + xor_out[72][1][2] + xor_out[73][1][2] + xor_out[74][1][2];
assign sum_out[15][1][2] = xor_out[75][1][2] + xor_out[76][1][2] + xor_out[77][1][2] + xor_out[78][1][2] + xor_out[79][1][2];
assign sum_out[16][1][2] = xor_out[80][1][2] + xor_out[81][1][2] + xor_out[82][1][2] + xor_out[83][1][2] + xor_out[84][1][2];
assign sum_out[17][1][2] = xor_out[85][1][2] + xor_out[86][1][2] + xor_out[87][1][2] + xor_out[88][1][2] + xor_out[89][1][2];
assign sum_out[18][1][2] = xor_out[90][1][2] + xor_out[91][1][2] + xor_out[92][1][2] + xor_out[93][1][2] + xor_out[94][1][2];
assign sum_out[19][1][2] = xor_out[95][1][2] + xor_out[96][1][2] + xor_out[97][1][2] + xor_out[98][1][2] + xor_out[99][1][2];

assign sum_out[0][1][3] = xor_out[0][1][3] + xor_out[1][1][3] + xor_out[2][1][3] + xor_out[3][1][3] + xor_out[4][1][3];
assign sum_out[1][1][3] = xor_out[5][1][3] + xor_out[6][1][3] + xor_out[7][1][3] + xor_out[8][1][3] + xor_out[9][1][3];
assign sum_out[2][1][3] = xor_out[10][1][3] + xor_out[11][1][3] + xor_out[12][1][3] + xor_out[13][1][3] + xor_out[14][1][3];
assign sum_out[3][1][3] = xor_out[15][1][3] + xor_out[16][1][3] + xor_out[17][1][3] + xor_out[18][1][3] + xor_out[19][1][3];
assign sum_out[4][1][3] = xor_out[20][1][3] + xor_out[21][1][3] + xor_out[22][1][3] + xor_out[23][1][3] + xor_out[24][1][3];
assign sum_out[5][1][3] = xor_out[25][1][3] + xor_out[26][1][3] + xor_out[27][1][3] + xor_out[28][1][3] + xor_out[29][1][3];
assign sum_out[6][1][3] = xor_out[30][1][3] + xor_out[31][1][3] + xor_out[32][1][3] + xor_out[33][1][3] + xor_out[34][1][3];
assign sum_out[7][1][3] = xor_out[35][1][3] + xor_out[36][1][3] + xor_out[37][1][3] + xor_out[38][1][3] + xor_out[39][1][3];
assign sum_out[8][1][3] = xor_out[40][1][3] + xor_out[41][1][3] + xor_out[42][1][3] + xor_out[43][1][3] + xor_out[44][1][3];
assign sum_out[9][1][3] = xor_out[45][1][3] + xor_out[46][1][3] + xor_out[47][1][3] + xor_out[48][1][3] + xor_out[49][1][3];
assign sum_out[10][1][3] = xor_out[50][1][3] + xor_out[51][1][3] + xor_out[52][1][3] + xor_out[53][1][3] + xor_out[54][1][3];
assign sum_out[11][1][3] = xor_out[55][1][3] + xor_out[56][1][3] + xor_out[57][1][3] + xor_out[58][1][3] + xor_out[59][1][3];
assign sum_out[12][1][3] = xor_out[60][1][3] + xor_out[61][1][3] + xor_out[62][1][3] + xor_out[63][1][3] + xor_out[64][1][3];
assign sum_out[13][1][3] = xor_out[65][1][3] + xor_out[66][1][3] + xor_out[67][1][3] + xor_out[68][1][3] + xor_out[69][1][3];
assign sum_out[14][1][3] = xor_out[70][1][3] + xor_out[71][1][3] + xor_out[72][1][3] + xor_out[73][1][3] + xor_out[74][1][3];
assign sum_out[15][1][3] = xor_out[75][1][3] + xor_out[76][1][3] + xor_out[77][1][3] + xor_out[78][1][3] + xor_out[79][1][3];
assign sum_out[16][1][3] = xor_out[80][1][3] + xor_out[81][1][3] + xor_out[82][1][3] + xor_out[83][1][3] + xor_out[84][1][3];
assign sum_out[17][1][3] = xor_out[85][1][3] + xor_out[86][1][3] + xor_out[87][1][3] + xor_out[88][1][3] + xor_out[89][1][3];
assign sum_out[18][1][3] = xor_out[90][1][3] + xor_out[91][1][3] + xor_out[92][1][3] + xor_out[93][1][3] + xor_out[94][1][3];
assign sum_out[19][1][3] = xor_out[95][1][3] + xor_out[96][1][3] + xor_out[97][1][3] + xor_out[98][1][3] + xor_out[99][1][3];

assign sum_out[0][1][4] = xor_out[0][1][4] + xor_out[1][1][4] + xor_out[2][1][4] + xor_out[3][1][4] + xor_out[4][1][4];
assign sum_out[1][1][4] = xor_out[5][1][4] + xor_out[6][1][4] + xor_out[7][1][4] + xor_out[8][1][4] + xor_out[9][1][4];
assign sum_out[2][1][4] = xor_out[10][1][4] + xor_out[11][1][4] + xor_out[12][1][4] + xor_out[13][1][4] + xor_out[14][1][4];
assign sum_out[3][1][4] = xor_out[15][1][4] + xor_out[16][1][4] + xor_out[17][1][4] + xor_out[18][1][4] + xor_out[19][1][4];
assign sum_out[4][1][4] = xor_out[20][1][4] + xor_out[21][1][4] + xor_out[22][1][4] + xor_out[23][1][4] + xor_out[24][1][4];
assign sum_out[5][1][4] = xor_out[25][1][4] + xor_out[26][1][4] + xor_out[27][1][4] + xor_out[28][1][4] + xor_out[29][1][4];
assign sum_out[6][1][4] = xor_out[30][1][4] + xor_out[31][1][4] + xor_out[32][1][4] + xor_out[33][1][4] + xor_out[34][1][4];
assign sum_out[7][1][4] = xor_out[35][1][4] + xor_out[36][1][4] + xor_out[37][1][4] + xor_out[38][1][4] + xor_out[39][1][4];
assign sum_out[8][1][4] = xor_out[40][1][4] + xor_out[41][1][4] + xor_out[42][1][4] + xor_out[43][1][4] + xor_out[44][1][4];
assign sum_out[9][1][4] = xor_out[45][1][4] + xor_out[46][1][4] + xor_out[47][1][4] + xor_out[48][1][4] + xor_out[49][1][4];
assign sum_out[10][1][4] = xor_out[50][1][4] + xor_out[51][1][4] + xor_out[52][1][4] + xor_out[53][1][4] + xor_out[54][1][4];
assign sum_out[11][1][4] = xor_out[55][1][4] + xor_out[56][1][4] + xor_out[57][1][4] + xor_out[58][1][4] + xor_out[59][1][4];
assign sum_out[12][1][4] = xor_out[60][1][4] + xor_out[61][1][4] + xor_out[62][1][4] + xor_out[63][1][4] + xor_out[64][1][4];
assign sum_out[13][1][4] = xor_out[65][1][4] + xor_out[66][1][4] + xor_out[67][1][4] + xor_out[68][1][4] + xor_out[69][1][4];
assign sum_out[14][1][4] = xor_out[70][1][4] + xor_out[71][1][4] + xor_out[72][1][4] + xor_out[73][1][4] + xor_out[74][1][4];
assign sum_out[15][1][4] = xor_out[75][1][4] + xor_out[76][1][4] + xor_out[77][1][4] + xor_out[78][1][4] + xor_out[79][1][4];
assign sum_out[16][1][4] = xor_out[80][1][4] + xor_out[81][1][4] + xor_out[82][1][4] + xor_out[83][1][4] + xor_out[84][1][4];
assign sum_out[17][1][4] = xor_out[85][1][4] + xor_out[86][1][4] + xor_out[87][1][4] + xor_out[88][1][4] + xor_out[89][1][4];
assign sum_out[18][1][4] = xor_out[90][1][4] + xor_out[91][1][4] + xor_out[92][1][4] + xor_out[93][1][4] + xor_out[94][1][4];
assign sum_out[19][1][4] = xor_out[95][1][4] + xor_out[96][1][4] + xor_out[97][1][4] + xor_out[98][1][4] + xor_out[99][1][4];

assign sum_out[0][1][5] = xor_out[0][1][5] + xor_out[1][1][5] + xor_out[2][1][5] + xor_out[3][1][5] + xor_out[4][1][5];
assign sum_out[1][1][5] = xor_out[5][1][5] + xor_out[6][1][5] + xor_out[7][1][5] + xor_out[8][1][5] + xor_out[9][1][5];
assign sum_out[2][1][5] = xor_out[10][1][5] + xor_out[11][1][5] + xor_out[12][1][5] + xor_out[13][1][5] + xor_out[14][1][5];
assign sum_out[3][1][5] = xor_out[15][1][5] + xor_out[16][1][5] + xor_out[17][1][5] + xor_out[18][1][5] + xor_out[19][1][5];
assign sum_out[4][1][5] = xor_out[20][1][5] + xor_out[21][1][5] + xor_out[22][1][5] + xor_out[23][1][5] + xor_out[24][1][5];
assign sum_out[5][1][5] = xor_out[25][1][5] + xor_out[26][1][5] + xor_out[27][1][5] + xor_out[28][1][5] + xor_out[29][1][5];
assign sum_out[6][1][5] = xor_out[30][1][5] + xor_out[31][1][5] + xor_out[32][1][5] + xor_out[33][1][5] + xor_out[34][1][5];
assign sum_out[7][1][5] = xor_out[35][1][5] + xor_out[36][1][5] + xor_out[37][1][5] + xor_out[38][1][5] + xor_out[39][1][5];
assign sum_out[8][1][5] = xor_out[40][1][5] + xor_out[41][1][5] + xor_out[42][1][5] + xor_out[43][1][5] + xor_out[44][1][5];
assign sum_out[9][1][5] = xor_out[45][1][5] + xor_out[46][1][5] + xor_out[47][1][5] + xor_out[48][1][5] + xor_out[49][1][5];
assign sum_out[10][1][5] = xor_out[50][1][5] + xor_out[51][1][5] + xor_out[52][1][5] + xor_out[53][1][5] + xor_out[54][1][5];
assign sum_out[11][1][5] = xor_out[55][1][5] + xor_out[56][1][5] + xor_out[57][1][5] + xor_out[58][1][5] + xor_out[59][1][5];
assign sum_out[12][1][5] = xor_out[60][1][5] + xor_out[61][1][5] + xor_out[62][1][5] + xor_out[63][1][5] + xor_out[64][1][5];
assign sum_out[13][1][5] = xor_out[65][1][5] + xor_out[66][1][5] + xor_out[67][1][5] + xor_out[68][1][5] + xor_out[69][1][5];
assign sum_out[14][1][5] = xor_out[70][1][5] + xor_out[71][1][5] + xor_out[72][1][5] + xor_out[73][1][5] + xor_out[74][1][5];
assign sum_out[15][1][5] = xor_out[75][1][5] + xor_out[76][1][5] + xor_out[77][1][5] + xor_out[78][1][5] + xor_out[79][1][5];
assign sum_out[16][1][5] = xor_out[80][1][5] + xor_out[81][1][5] + xor_out[82][1][5] + xor_out[83][1][5] + xor_out[84][1][5];
assign sum_out[17][1][5] = xor_out[85][1][5] + xor_out[86][1][5] + xor_out[87][1][5] + xor_out[88][1][5] + xor_out[89][1][5];
assign sum_out[18][1][5] = xor_out[90][1][5] + xor_out[91][1][5] + xor_out[92][1][5] + xor_out[93][1][5] + xor_out[94][1][5];
assign sum_out[19][1][5] = xor_out[95][1][5] + xor_out[96][1][5] + xor_out[97][1][5] + xor_out[98][1][5] + xor_out[99][1][5];

assign sum_out[0][1][6] = xor_out[0][1][6] + xor_out[1][1][6] + xor_out[2][1][6] + xor_out[3][1][6] + xor_out[4][1][6];
assign sum_out[1][1][6] = xor_out[5][1][6] + xor_out[6][1][6] + xor_out[7][1][6] + xor_out[8][1][6] + xor_out[9][1][6];
assign sum_out[2][1][6] = xor_out[10][1][6] + xor_out[11][1][6] + xor_out[12][1][6] + xor_out[13][1][6] + xor_out[14][1][6];
assign sum_out[3][1][6] = xor_out[15][1][6] + xor_out[16][1][6] + xor_out[17][1][6] + xor_out[18][1][6] + xor_out[19][1][6];
assign sum_out[4][1][6] = xor_out[20][1][6] + xor_out[21][1][6] + xor_out[22][1][6] + xor_out[23][1][6] + xor_out[24][1][6];
assign sum_out[5][1][6] = xor_out[25][1][6] + xor_out[26][1][6] + xor_out[27][1][6] + xor_out[28][1][6] + xor_out[29][1][6];
assign sum_out[6][1][6] = xor_out[30][1][6] + xor_out[31][1][6] + xor_out[32][1][6] + xor_out[33][1][6] + xor_out[34][1][6];
assign sum_out[7][1][6] = xor_out[35][1][6] + xor_out[36][1][6] + xor_out[37][1][6] + xor_out[38][1][6] + xor_out[39][1][6];
assign sum_out[8][1][6] = xor_out[40][1][6] + xor_out[41][1][6] + xor_out[42][1][6] + xor_out[43][1][6] + xor_out[44][1][6];
assign sum_out[9][1][6] = xor_out[45][1][6] + xor_out[46][1][6] + xor_out[47][1][6] + xor_out[48][1][6] + xor_out[49][1][6];
assign sum_out[10][1][6] = xor_out[50][1][6] + xor_out[51][1][6] + xor_out[52][1][6] + xor_out[53][1][6] + xor_out[54][1][6];
assign sum_out[11][1][6] = xor_out[55][1][6] + xor_out[56][1][6] + xor_out[57][1][6] + xor_out[58][1][6] + xor_out[59][1][6];
assign sum_out[12][1][6] = xor_out[60][1][6] + xor_out[61][1][6] + xor_out[62][1][6] + xor_out[63][1][6] + xor_out[64][1][6];
assign sum_out[13][1][6] = xor_out[65][1][6] + xor_out[66][1][6] + xor_out[67][1][6] + xor_out[68][1][6] + xor_out[69][1][6];
assign sum_out[14][1][6] = xor_out[70][1][6] + xor_out[71][1][6] + xor_out[72][1][6] + xor_out[73][1][6] + xor_out[74][1][6];
assign sum_out[15][1][6] = xor_out[75][1][6] + xor_out[76][1][6] + xor_out[77][1][6] + xor_out[78][1][6] + xor_out[79][1][6];
assign sum_out[16][1][6] = xor_out[80][1][6] + xor_out[81][1][6] + xor_out[82][1][6] + xor_out[83][1][6] + xor_out[84][1][6];
assign sum_out[17][1][6] = xor_out[85][1][6] + xor_out[86][1][6] + xor_out[87][1][6] + xor_out[88][1][6] + xor_out[89][1][6];
assign sum_out[18][1][6] = xor_out[90][1][6] + xor_out[91][1][6] + xor_out[92][1][6] + xor_out[93][1][6] + xor_out[94][1][6];
assign sum_out[19][1][6] = xor_out[95][1][6] + xor_out[96][1][6] + xor_out[97][1][6] + xor_out[98][1][6] + xor_out[99][1][6];

assign sum_out[0][1][7] = xor_out[0][1][7] + xor_out[1][1][7] + xor_out[2][1][7] + xor_out[3][1][7] + xor_out[4][1][7];
assign sum_out[1][1][7] = xor_out[5][1][7] + xor_out[6][1][7] + xor_out[7][1][7] + xor_out[8][1][7] + xor_out[9][1][7];
assign sum_out[2][1][7] = xor_out[10][1][7] + xor_out[11][1][7] + xor_out[12][1][7] + xor_out[13][1][7] + xor_out[14][1][7];
assign sum_out[3][1][7] = xor_out[15][1][7] + xor_out[16][1][7] + xor_out[17][1][7] + xor_out[18][1][7] + xor_out[19][1][7];
assign sum_out[4][1][7] = xor_out[20][1][7] + xor_out[21][1][7] + xor_out[22][1][7] + xor_out[23][1][7] + xor_out[24][1][7];
assign sum_out[5][1][7] = xor_out[25][1][7] + xor_out[26][1][7] + xor_out[27][1][7] + xor_out[28][1][7] + xor_out[29][1][7];
assign sum_out[6][1][7] = xor_out[30][1][7] + xor_out[31][1][7] + xor_out[32][1][7] + xor_out[33][1][7] + xor_out[34][1][7];
assign sum_out[7][1][7] = xor_out[35][1][7] + xor_out[36][1][7] + xor_out[37][1][7] + xor_out[38][1][7] + xor_out[39][1][7];
assign sum_out[8][1][7] = xor_out[40][1][7] + xor_out[41][1][7] + xor_out[42][1][7] + xor_out[43][1][7] + xor_out[44][1][7];
assign sum_out[9][1][7] = xor_out[45][1][7] + xor_out[46][1][7] + xor_out[47][1][7] + xor_out[48][1][7] + xor_out[49][1][7];
assign sum_out[10][1][7] = xor_out[50][1][7] + xor_out[51][1][7] + xor_out[52][1][7] + xor_out[53][1][7] + xor_out[54][1][7];
assign sum_out[11][1][7] = xor_out[55][1][7] + xor_out[56][1][7] + xor_out[57][1][7] + xor_out[58][1][7] + xor_out[59][1][7];
assign sum_out[12][1][7] = xor_out[60][1][7] + xor_out[61][1][7] + xor_out[62][1][7] + xor_out[63][1][7] + xor_out[64][1][7];
assign sum_out[13][1][7] = xor_out[65][1][7] + xor_out[66][1][7] + xor_out[67][1][7] + xor_out[68][1][7] + xor_out[69][1][7];
assign sum_out[14][1][7] = xor_out[70][1][7] + xor_out[71][1][7] + xor_out[72][1][7] + xor_out[73][1][7] + xor_out[74][1][7];
assign sum_out[15][1][7] = xor_out[75][1][7] + xor_out[76][1][7] + xor_out[77][1][7] + xor_out[78][1][7] + xor_out[79][1][7];
assign sum_out[16][1][7] = xor_out[80][1][7] + xor_out[81][1][7] + xor_out[82][1][7] + xor_out[83][1][7] + xor_out[84][1][7];
assign sum_out[17][1][7] = xor_out[85][1][7] + xor_out[86][1][7] + xor_out[87][1][7] + xor_out[88][1][7] + xor_out[89][1][7];
assign sum_out[18][1][7] = xor_out[90][1][7] + xor_out[91][1][7] + xor_out[92][1][7] + xor_out[93][1][7] + xor_out[94][1][7];
assign sum_out[19][1][7] = xor_out[95][1][7] + xor_out[96][1][7] + xor_out[97][1][7] + xor_out[98][1][7] + xor_out[99][1][7];

assign sum_out[0][1][8] = xor_out[0][1][8] + xor_out[1][1][8] + xor_out[2][1][8] + xor_out[3][1][8] + xor_out[4][1][8];
assign sum_out[1][1][8] = xor_out[5][1][8] + xor_out[6][1][8] + xor_out[7][1][8] + xor_out[8][1][8] + xor_out[9][1][8];
assign sum_out[2][1][8] = xor_out[10][1][8] + xor_out[11][1][8] + xor_out[12][1][8] + xor_out[13][1][8] + xor_out[14][1][8];
assign sum_out[3][1][8] = xor_out[15][1][8] + xor_out[16][1][8] + xor_out[17][1][8] + xor_out[18][1][8] + xor_out[19][1][8];
assign sum_out[4][1][8] = xor_out[20][1][8] + xor_out[21][1][8] + xor_out[22][1][8] + xor_out[23][1][8] + xor_out[24][1][8];
assign sum_out[5][1][8] = xor_out[25][1][8] + xor_out[26][1][8] + xor_out[27][1][8] + xor_out[28][1][8] + xor_out[29][1][8];
assign sum_out[6][1][8] = xor_out[30][1][8] + xor_out[31][1][8] + xor_out[32][1][8] + xor_out[33][1][8] + xor_out[34][1][8];
assign sum_out[7][1][8] = xor_out[35][1][8] + xor_out[36][1][8] + xor_out[37][1][8] + xor_out[38][1][8] + xor_out[39][1][8];
assign sum_out[8][1][8] = xor_out[40][1][8] + xor_out[41][1][8] + xor_out[42][1][8] + xor_out[43][1][8] + xor_out[44][1][8];
assign sum_out[9][1][8] = xor_out[45][1][8] + xor_out[46][1][8] + xor_out[47][1][8] + xor_out[48][1][8] + xor_out[49][1][8];
assign sum_out[10][1][8] = xor_out[50][1][8] + xor_out[51][1][8] + xor_out[52][1][8] + xor_out[53][1][8] + xor_out[54][1][8];
assign sum_out[11][1][8] = xor_out[55][1][8] + xor_out[56][1][8] + xor_out[57][1][8] + xor_out[58][1][8] + xor_out[59][1][8];
assign sum_out[12][1][8] = xor_out[60][1][8] + xor_out[61][1][8] + xor_out[62][1][8] + xor_out[63][1][8] + xor_out[64][1][8];
assign sum_out[13][1][8] = xor_out[65][1][8] + xor_out[66][1][8] + xor_out[67][1][8] + xor_out[68][1][8] + xor_out[69][1][8];
assign sum_out[14][1][8] = xor_out[70][1][8] + xor_out[71][1][8] + xor_out[72][1][8] + xor_out[73][1][8] + xor_out[74][1][8];
assign sum_out[15][1][8] = xor_out[75][1][8] + xor_out[76][1][8] + xor_out[77][1][8] + xor_out[78][1][8] + xor_out[79][1][8];
assign sum_out[16][1][8] = xor_out[80][1][8] + xor_out[81][1][8] + xor_out[82][1][8] + xor_out[83][1][8] + xor_out[84][1][8];
assign sum_out[17][1][8] = xor_out[85][1][8] + xor_out[86][1][8] + xor_out[87][1][8] + xor_out[88][1][8] + xor_out[89][1][8];
assign sum_out[18][1][8] = xor_out[90][1][8] + xor_out[91][1][8] + xor_out[92][1][8] + xor_out[93][1][8] + xor_out[94][1][8];
assign sum_out[19][1][8] = xor_out[95][1][8] + xor_out[96][1][8] + xor_out[97][1][8] + xor_out[98][1][8] + xor_out[99][1][8];

assign sum_out[0][1][9] = xor_out[0][1][9] + xor_out[1][1][9] + xor_out[2][1][9] + xor_out[3][1][9] + xor_out[4][1][9];
assign sum_out[1][1][9] = xor_out[5][1][9] + xor_out[6][1][9] + xor_out[7][1][9] + xor_out[8][1][9] + xor_out[9][1][9];
assign sum_out[2][1][9] = xor_out[10][1][9] + xor_out[11][1][9] + xor_out[12][1][9] + xor_out[13][1][9] + xor_out[14][1][9];
assign sum_out[3][1][9] = xor_out[15][1][9] + xor_out[16][1][9] + xor_out[17][1][9] + xor_out[18][1][9] + xor_out[19][1][9];
assign sum_out[4][1][9] = xor_out[20][1][9] + xor_out[21][1][9] + xor_out[22][1][9] + xor_out[23][1][9] + xor_out[24][1][9];
assign sum_out[5][1][9] = xor_out[25][1][9] + xor_out[26][1][9] + xor_out[27][1][9] + xor_out[28][1][9] + xor_out[29][1][9];
assign sum_out[6][1][9] = xor_out[30][1][9] + xor_out[31][1][9] + xor_out[32][1][9] + xor_out[33][1][9] + xor_out[34][1][9];
assign sum_out[7][1][9] = xor_out[35][1][9] + xor_out[36][1][9] + xor_out[37][1][9] + xor_out[38][1][9] + xor_out[39][1][9];
assign sum_out[8][1][9] = xor_out[40][1][9] + xor_out[41][1][9] + xor_out[42][1][9] + xor_out[43][1][9] + xor_out[44][1][9];
assign sum_out[9][1][9] = xor_out[45][1][9] + xor_out[46][1][9] + xor_out[47][1][9] + xor_out[48][1][9] + xor_out[49][1][9];
assign sum_out[10][1][9] = xor_out[50][1][9] + xor_out[51][1][9] + xor_out[52][1][9] + xor_out[53][1][9] + xor_out[54][1][9];
assign sum_out[11][1][9] = xor_out[55][1][9] + xor_out[56][1][9] + xor_out[57][1][9] + xor_out[58][1][9] + xor_out[59][1][9];
assign sum_out[12][1][9] = xor_out[60][1][9] + xor_out[61][1][9] + xor_out[62][1][9] + xor_out[63][1][9] + xor_out[64][1][9];
assign sum_out[13][1][9] = xor_out[65][1][9] + xor_out[66][1][9] + xor_out[67][1][9] + xor_out[68][1][9] + xor_out[69][1][9];
assign sum_out[14][1][9] = xor_out[70][1][9] + xor_out[71][1][9] + xor_out[72][1][9] + xor_out[73][1][9] + xor_out[74][1][9];
assign sum_out[15][1][9] = xor_out[75][1][9] + xor_out[76][1][9] + xor_out[77][1][9] + xor_out[78][1][9] + xor_out[79][1][9];
assign sum_out[16][1][9] = xor_out[80][1][9] + xor_out[81][1][9] + xor_out[82][1][9] + xor_out[83][1][9] + xor_out[84][1][9];
assign sum_out[17][1][9] = xor_out[85][1][9] + xor_out[86][1][9] + xor_out[87][1][9] + xor_out[88][1][9] + xor_out[89][1][9];
assign sum_out[18][1][9] = xor_out[90][1][9] + xor_out[91][1][9] + xor_out[92][1][9] + xor_out[93][1][9] + xor_out[94][1][9];
assign sum_out[19][1][9] = xor_out[95][1][9] + xor_out[96][1][9] + xor_out[97][1][9] + xor_out[98][1][9] + xor_out[99][1][9];

assign sum_out[0][1][10] = xor_out[0][1][10] + xor_out[1][1][10] + xor_out[2][1][10] + xor_out[3][1][10] + xor_out[4][1][10];
assign sum_out[1][1][10] = xor_out[5][1][10] + xor_out[6][1][10] + xor_out[7][1][10] + xor_out[8][1][10] + xor_out[9][1][10];
assign sum_out[2][1][10] = xor_out[10][1][10] + xor_out[11][1][10] + xor_out[12][1][10] + xor_out[13][1][10] + xor_out[14][1][10];
assign sum_out[3][1][10] = xor_out[15][1][10] + xor_out[16][1][10] + xor_out[17][1][10] + xor_out[18][1][10] + xor_out[19][1][10];
assign sum_out[4][1][10] = xor_out[20][1][10] + xor_out[21][1][10] + xor_out[22][1][10] + xor_out[23][1][10] + xor_out[24][1][10];
assign sum_out[5][1][10] = xor_out[25][1][10] + xor_out[26][1][10] + xor_out[27][1][10] + xor_out[28][1][10] + xor_out[29][1][10];
assign sum_out[6][1][10] = xor_out[30][1][10] + xor_out[31][1][10] + xor_out[32][1][10] + xor_out[33][1][10] + xor_out[34][1][10];
assign sum_out[7][1][10] = xor_out[35][1][10] + xor_out[36][1][10] + xor_out[37][1][10] + xor_out[38][1][10] + xor_out[39][1][10];
assign sum_out[8][1][10] = xor_out[40][1][10] + xor_out[41][1][10] + xor_out[42][1][10] + xor_out[43][1][10] + xor_out[44][1][10];
assign sum_out[9][1][10] = xor_out[45][1][10] + xor_out[46][1][10] + xor_out[47][1][10] + xor_out[48][1][10] + xor_out[49][1][10];
assign sum_out[10][1][10] = xor_out[50][1][10] + xor_out[51][1][10] + xor_out[52][1][10] + xor_out[53][1][10] + xor_out[54][1][10];
assign sum_out[11][1][10] = xor_out[55][1][10] + xor_out[56][1][10] + xor_out[57][1][10] + xor_out[58][1][10] + xor_out[59][1][10];
assign sum_out[12][1][10] = xor_out[60][1][10] + xor_out[61][1][10] + xor_out[62][1][10] + xor_out[63][1][10] + xor_out[64][1][10];
assign sum_out[13][1][10] = xor_out[65][1][10] + xor_out[66][1][10] + xor_out[67][1][10] + xor_out[68][1][10] + xor_out[69][1][10];
assign sum_out[14][1][10] = xor_out[70][1][10] + xor_out[71][1][10] + xor_out[72][1][10] + xor_out[73][1][10] + xor_out[74][1][10];
assign sum_out[15][1][10] = xor_out[75][1][10] + xor_out[76][1][10] + xor_out[77][1][10] + xor_out[78][1][10] + xor_out[79][1][10];
assign sum_out[16][1][10] = xor_out[80][1][10] + xor_out[81][1][10] + xor_out[82][1][10] + xor_out[83][1][10] + xor_out[84][1][10];
assign sum_out[17][1][10] = xor_out[85][1][10] + xor_out[86][1][10] + xor_out[87][1][10] + xor_out[88][1][10] + xor_out[89][1][10];
assign sum_out[18][1][10] = xor_out[90][1][10] + xor_out[91][1][10] + xor_out[92][1][10] + xor_out[93][1][10] + xor_out[94][1][10];
assign sum_out[19][1][10] = xor_out[95][1][10] + xor_out[96][1][10] + xor_out[97][1][10] + xor_out[98][1][10] + xor_out[99][1][10];

assign sum_out[0][1][11] = xor_out[0][1][11] + xor_out[1][1][11] + xor_out[2][1][11] + xor_out[3][1][11] + xor_out[4][1][11];
assign sum_out[1][1][11] = xor_out[5][1][11] + xor_out[6][1][11] + xor_out[7][1][11] + xor_out[8][1][11] + xor_out[9][1][11];
assign sum_out[2][1][11] = xor_out[10][1][11] + xor_out[11][1][11] + xor_out[12][1][11] + xor_out[13][1][11] + xor_out[14][1][11];
assign sum_out[3][1][11] = xor_out[15][1][11] + xor_out[16][1][11] + xor_out[17][1][11] + xor_out[18][1][11] + xor_out[19][1][11];
assign sum_out[4][1][11] = xor_out[20][1][11] + xor_out[21][1][11] + xor_out[22][1][11] + xor_out[23][1][11] + xor_out[24][1][11];
assign sum_out[5][1][11] = xor_out[25][1][11] + xor_out[26][1][11] + xor_out[27][1][11] + xor_out[28][1][11] + xor_out[29][1][11];
assign sum_out[6][1][11] = xor_out[30][1][11] + xor_out[31][1][11] + xor_out[32][1][11] + xor_out[33][1][11] + xor_out[34][1][11];
assign sum_out[7][1][11] = xor_out[35][1][11] + xor_out[36][1][11] + xor_out[37][1][11] + xor_out[38][1][11] + xor_out[39][1][11];
assign sum_out[8][1][11] = xor_out[40][1][11] + xor_out[41][1][11] + xor_out[42][1][11] + xor_out[43][1][11] + xor_out[44][1][11];
assign sum_out[9][1][11] = xor_out[45][1][11] + xor_out[46][1][11] + xor_out[47][1][11] + xor_out[48][1][11] + xor_out[49][1][11];
assign sum_out[10][1][11] = xor_out[50][1][11] + xor_out[51][1][11] + xor_out[52][1][11] + xor_out[53][1][11] + xor_out[54][1][11];
assign sum_out[11][1][11] = xor_out[55][1][11] + xor_out[56][1][11] + xor_out[57][1][11] + xor_out[58][1][11] + xor_out[59][1][11];
assign sum_out[12][1][11] = xor_out[60][1][11] + xor_out[61][1][11] + xor_out[62][1][11] + xor_out[63][1][11] + xor_out[64][1][11];
assign sum_out[13][1][11] = xor_out[65][1][11] + xor_out[66][1][11] + xor_out[67][1][11] + xor_out[68][1][11] + xor_out[69][1][11];
assign sum_out[14][1][11] = xor_out[70][1][11] + xor_out[71][1][11] + xor_out[72][1][11] + xor_out[73][1][11] + xor_out[74][1][11];
assign sum_out[15][1][11] = xor_out[75][1][11] + xor_out[76][1][11] + xor_out[77][1][11] + xor_out[78][1][11] + xor_out[79][1][11];
assign sum_out[16][1][11] = xor_out[80][1][11] + xor_out[81][1][11] + xor_out[82][1][11] + xor_out[83][1][11] + xor_out[84][1][11];
assign sum_out[17][1][11] = xor_out[85][1][11] + xor_out[86][1][11] + xor_out[87][1][11] + xor_out[88][1][11] + xor_out[89][1][11];
assign sum_out[18][1][11] = xor_out[90][1][11] + xor_out[91][1][11] + xor_out[92][1][11] + xor_out[93][1][11] + xor_out[94][1][11];
assign sum_out[19][1][11] = xor_out[95][1][11] + xor_out[96][1][11] + xor_out[97][1][11] + xor_out[98][1][11] + xor_out[99][1][11];

assign sum_out[0][1][12] = xor_out[0][1][12] + xor_out[1][1][12] + xor_out[2][1][12] + xor_out[3][1][12] + xor_out[4][1][12];
assign sum_out[1][1][12] = xor_out[5][1][12] + xor_out[6][1][12] + xor_out[7][1][12] + xor_out[8][1][12] + xor_out[9][1][12];
assign sum_out[2][1][12] = xor_out[10][1][12] + xor_out[11][1][12] + xor_out[12][1][12] + xor_out[13][1][12] + xor_out[14][1][12];
assign sum_out[3][1][12] = xor_out[15][1][12] + xor_out[16][1][12] + xor_out[17][1][12] + xor_out[18][1][12] + xor_out[19][1][12];
assign sum_out[4][1][12] = xor_out[20][1][12] + xor_out[21][1][12] + xor_out[22][1][12] + xor_out[23][1][12] + xor_out[24][1][12];
assign sum_out[5][1][12] = xor_out[25][1][12] + xor_out[26][1][12] + xor_out[27][1][12] + xor_out[28][1][12] + xor_out[29][1][12];
assign sum_out[6][1][12] = xor_out[30][1][12] + xor_out[31][1][12] + xor_out[32][1][12] + xor_out[33][1][12] + xor_out[34][1][12];
assign sum_out[7][1][12] = xor_out[35][1][12] + xor_out[36][1][12] + xor_out[37][1][12] + xor_out[38][1][12] + xor_out[39][1][12];
assign sum_out[8][1][12] = xor_out[40][1][12] + xor_out[41][1][12] + xor_out[42][1][12] + xor_out[43][1][12] + xor_out[44][1][12];
assign sum_out[9][1][12] = xor_out[45][1][12] + xor_out[46][1][12] + xor_out[47][1][12] + xor_out[48][1][12] + xor_out[49][1][12];
assign sum_out[10][1][12] = xor_out[50][1][12] + xor_out[51][1][12] + xor_out[52][1][12] + xor_out[53][1][12] + xor_out[54][1][12];
assign sum_out[11][1][12] = xor_out[55][1][12] + xor_out[56][1][12] + xor_out[57][1][12] + xor_out[58][1][12] + xor_out[59][1][12];
assign sum_out[12][1][12] = xor_out[60][1][12] + xor_out[61][1][12] + xor_out[62][1][12] + xor_out[63][1][12] + xor_out[64][1][12];
assign sum_out[13][1][12] = xor_out[65][1][12] + xor_out[66][1][12] + xor_out[67][1][12] + xor_out[68][1][12] + xor_out[69][1][12];
assign sum_out[14][1][12] = xor_out[70][1][12] + xor_out[71][1][12] + xor_out[72][1][12] + xor_out[73][1][12] + xor_out[74][1][12];
assign sum_out[15][1][12] = xor_out[75][1][12] + xor_out[76][1][12] + xor_out[77][1][12] + xor_out[78][1][12] + xor_out[79][1][12];
assign sum_out[16][1][12] = xor_out[80][1][12] + xor_out[81][1][12] + xor_out[82][1][12] + xor_out[83][1][12] + xor_out[84][1][12];
assign sum_out[17][1][12] = xor_out[85][1][12] + xor_out[86][1][12] + xor_out[87][1][12] + xor_out[88][1][12] + xor_out[89][1][12];
assign sum_out[18][1][12] = xor_out[90][1][12] + xor_out[91][1][12] + xor_out[92][1][12] + xor_out[93][1][12] + xor_out[94][1][12];
assign sum_out[19][1][12] = xor_out[95][1][12] + xor_out[96][1][12] + xor_out[97][1][12] + xor_out[98][1][12] + xor_out[99][1][12];

assign sum_out[0][1][13] = xor_out[0][1][13] + xor_out[1][1][13] + xor_out[2][1][13] + xor_out[3][1][13] + xor_out[4][1][13];
assign sum_out[1][1][13] = xor_out[5][1][13] + xor_out[6][1][13] + xor_out[7][1][13] + xor_out[8][1][13] + xor_out[9][1][13];
assign sum_out[2][1][13] = xor_out[10][1][13] + xor_out[11][1][13] + xor_out[12][1][13] + xor_out[13][1][13] + xor_out[14][1][13];
assign sum_out[3][1][13] = xor_out[15][1][13] + xor_out[16][1][13] + xor_out[17][1][13] + xor_out[18][1][13] + xor_out[19][1][13];
assign sum_out[4][1][13] = xor_out[20][1][13] + xor_out[21][1][13] + xor_out[22][1][13] + xor_out[23][1][13] + xor_out[24][1][13];
assign sum_out[5][1][13] = xor_out[25][1][13] + xor_out[26][1][13] + xor_out[27][1][13] + xor_out[28][1][13] + xor_out[29][1][13];
assign sum_out[6][1][13] = xor_out[30][1][13] + xor_out[31][1][13] + xor_out[32][1][13] + xor_out[33][1][13] + xor_out[34][1][13];
assign sum_out[7][1][13] = xor_out[35][1][13] + xor_out[36][1][13] + xor_out[37][1][13] + xor_out[38][1][13] + xor_out[39][1][13];
assign sum_out[8][1][13] = xor_out[40][1][13] + xor_out[41][1][13] + xor_out[42][1][13] + xor_out[43][1][13] + xor_out[44][1][13];
assign sum_out[9][1][13] = xor_out[45][1][13] + xor_out[46][1][13] + xor_out[47][1][13] + xor_out[48][1][13] + xor_out[49][1][13];
assign sum_out[10][1][13] = xor_out[50][1][13] + xor_out[51][1][13] + xor_out[52][1][13] + xor_out[53][1][13] + xor_out[54][1][13];
assign sum_out[11][1][13] = xor_out[55][1][13] + xor_out[56][1][13] + xor_out[57][1][13] + xor_out[58][1][13] + xor_out[59][1][13];
assign sum_out[12][1][13] = xor_out[60][1][13] + xor_out[61][1][13] + xor_out[62][1][13] + xor_out[63][1][13] + xor_out[64][1][13];
assign sum_out[13][1][13] = xor_out[65][1][13] + xor_out[66][1][13] + xor_out[67][1][13] + xor_out[68][1][13] + xor_out[69][1][13];
assign sum_out[14][1][13] = xor_out[70][1][13] + xor_out[71][1][13] + xor_out[72][1][13] + xor_out[73][1][13] + xor_out[74][1][13];
assign sum_out[15][1][13] = xor_out[75][1][13] + xor_out[76][1][13] + xor_out[77][1][13] + xor_out[78][1][13] + xor_out[79][1][13];
assign sum_out[16][1][13] = xor_out[80][1][13] + xor_out[81][1][13] + xor_out[82][1][13] + xor_out[83][1][13] + xor_out[84][1][13];
assign sum_out[17][1][13] = xor_out[85][1][13] + xor_out[86][1][13] + xor_out[87][1][13] + xor_out[88][1][13] + xor_out[89][1][13];
assign sum_out[18][1][13] = xor_out[90][1][13] + xor_out[91][1][13] + xor_out[92][1][13] + xor_out[93][1][13] + xor_out[94][1][13];
assign sum_out[19][1][13] = xor_out[95][1][13] + xor_out[96][1][13] + xor_out[97][1][13] + xor_out[98][1][13] + xor_out[99][1][13];

assign sum_out[0][1][14] = xor_out[0][1][14] + xor_out[1][1][14] + xor_out[2][1][14] + xor_out[3][1][14] + xor_out[4][1][14];
assign sum_out[1][1][14] = xor_out[5][1][14] + xor_out[6][1][14] + xor_out[7][1][14] + xor_out[8][1][14] + xor_out[9][1][14];
assign sum_out[2][1][14] = xor_out[10][1][14] + xor_out[11][1][14] + xor_out[12][1][14] + xor_out[13][1][14] + xor_out[14][1][14];
assign sum_out[3][1][14] = xor_out[15][1][14] + xor_out[16][1][14] + xor_out[17][1][14] + xor_out[18][1][14] + xor_out[19][1][14];
assign sum_out[4][1][14] = xor_out[20][1][14] + xor_out[21][1][14] + xor_out[22][1][14] + xor_out[23][1][14] + xor_out[24][1][14];
assign sum_out[5][1][14] = xor_out[25][1][14] + xor_out[26][1][14] + xor_out[27][1][14] + xor_out[28][1][14] + xor_out[29][1][14];
assign sum_out[6][1][14] = xor_out[30][1][14] + xor_out[31][1][14] + xor_out[32][1][14] + xor_out[33][1][14] + xor_out[34][1][14];
assign sum_out[7][1][14] = xor_out[35][1][14] + xor_out[36][1][14] + xor_out[37][1][14] + xor_out[38][1][14] + xor_out[39][1][14];
assign sum_out[8][1][14] = xor_out[40][1][14] + xor_out[41][1][14] + xor_out[42][1][14] + xor_out[43][1][14] + xor_out[44][1][14];
assign sum_out[9][1][14] = xor_out[45][1][14] + xor_out[46][1][14] + xor_out[47][1][14] + xor_out[48][1][14] + xor_out[49][1][14];
assign sum_out[10][1][14] = xor_out[50][1][14] + xor_out[51][1][14] + xor_out[52][1][14] + xor_out[53][1][14] + xor_out[54][1][14];
assign sum_out[11][1][14] = xor_out[55][1][14] + xor_out[56][1][14] + xor_out[57][1][14] + xor_out[58][1][14] + xor_out[59][1][14];
assign sum_out[12][1][14] = xor_out[60][1][14] + xor_out[61][1][14] + xor_out[62][1][14] + xor_out[63][1][14] + xor_out[64][1][14];
assign sum_out[13][1][14] = xor_out[65][1][14] + xor_out[66][1][14] + xor_out[67][1][14] + xor_out[68][1][14] + xor_out[69][1][14];
assign sum_out[14][1][14] = xor_out[70][1][14] + xor_out[71][1][14] + xor_out[72][1][14] + xor_out[73][1][14] + xor_out[74][1][14];
assign sum_out[15][1][14] = xor_out[75][1][14] + xor_out[76][1][14] + xor_out[77][1][14] + xor_out[78][1][14] + xor_out[79][1][14];
assign sum_out[16][1][14] = xor_out[80][1][14] + xor_out[81][1][14] + xor_out[82][1][14] + xor_out[83][1][14] + xor_out[84][1][14];
assign sum_out[17][1][14] = xor_out[85][1][14] + xor_out[86][1][14] + xor_out[87][1][14] + xor_out[88][1][14] + xor_out[89][1][14];
assign sum_out[18][1][14] = xor_out[90][1][14] + xor_out[91][1][14] + xor_out[92][1][14] + xor_out[93][1][14] + xor_out[94][1][14];
assign sum_out[19][1][14] = xor_out[95][1][14] + xor_out[96][1][14] + xor_out[97][1][14] + xor_out[98][1][14] + xor_out[99][1][14];

assign sum_out[0][1][15] = xor_out[0][1][15] + xor_out[1][1][15] + xor_out[2][1][15] + xor_out[3][1][15] + xor_out[4][1][15];
assign sum_out[1][1][15] = xor_out[5][1][15] + xor_out[6][1][15] + xor_out[7][1][15] + xor_out[8][1][15] + xor_out[9][1][15];
assign sum_out[2][1][15] = xor_out[10][1][15] + xor_out[11][1][15] + xor_out[12][1][15] + xor_out[13][1][15] + xor_out[14][1][15];
assign sum_out[3][1][15] = xor_out[15][1][15] + xor_out[16][1][15] + xor_out[17][1][15] + xor_out[18][1][15] + xor_out[19][1][15];
assign sum_out[4][1][15] = xor_out[20][1][15] + xor_out[21][1][15] + xor_out[22][1][15] + xor_out[23][1][15] + xor_out[24][1][15];
assign sum_out[5][1][15] = xor_out[25][1][15] + xor_out[26][1][15] + xor_out[27][1][15] + xor_out[28][1][15] + xor_out[29][1][15];
assign sum_out[6][1][15] = xor_out[30][1][15] + xor_out[31][1][15] + xor_out[32][1][15] + xor_out[33][1][15] + xor_out[34][1][15];
assign sum_out[7][1][15] = xor_out[35][1][15] + xor_out[36][1][15] + xor_out[37][1][15] + xor_out[38][1][15] + xor_out[39][1][15];
assign sum_out[8][1][15] = xor_out[40][1][15] + xor_out[41][1][15] + xor_out[42][1][15] + xor_out[43][1][15] + xor_out[44][1][15];
assign sum_out[9][1][15] = xor_out[45][1][15] + xor_out[46][1][15] + xor_out[47][1][15] + xor_out[48][1][15] + xor_out[49][1][15];
assign sum_out[10][1][15] = xor_out[50][1][15] + xor_out[51][1][15] + xor_out[52][1][15] + xor_out[53][1][15] + xor_out[54][1][15];
assign sum_out[11][1][15] = xor_out[55][1][15] + xor_out[56][1][15] + xor_out[57][1][15] + xor_out[58][1][15] + xor_out[59][1][15];
assign sum_out[12][1][15] = xor_out[60][1][15] + xor_out[61][1][15] + xor_out[62][1][15] + xor_out[63][1][15] + xor_out[64][1][15];
assign sum_out[13][1][15] = xor_out[65][1][15] + xor_out[66][1][15] + xor_out[67][1][15] + xor_out[68][1][15] + xor_out[69][1][15];
assign sum_out[14][1][15] = xor_out[70][1][15] + xor_out[71][1][15] + xor_out[72][1][15] + xor_out[73][1][15] + xor_out[74][1][15];
assign sum_out[15][1][15] = xor_out[75][1][15] + xor_out[76][1][15] + xor_out[77][1][15] + xor_out[78][1][15] + xor_out[79][1][15];
assign sum_out[16][1][15] = xor_out[80][1][15] + xor_out[81][1][15] + xor_out[82][1][15] + xor_out[83][1][15] + xor_out[84][1][15];
assign sum_out[17][1][15] = xor_out[85][1][15] + xor_out[86][1][15] + xor_out[87][1][15] + xor_out[88][1][15] + xor_out[89][1][15];
assign sum_out[18][1][15] = xor_out[90][1][15] + xor_out[91][1][15] + xor_out[92][1][15] + xor_out[93][1][15] + xor_out[94][1][15];
assign sum_out[19][1][15] = xor_out[95][1][15] + xor_out[96][1][15] + xor_out[97][1][15] + xor_out[98][1][15] + xor_out[99][1][15];

assign sum_out[0][1][16] = xor_out[0][1][16] + xor_out[1][1][16] + xor_out[2][1][16] + xor_out[3][1][16] + xor_out[4][1][16];
assign sum_out[1][1][16] = xor_out[5][1][16] + xor_out[6][1][16] + xor_out[7][1][16] + xor_out[8][1][16] + xor_out[9][1][16];
assign sum_out[2][1][16] = xor_out[10][1][16] + xor_out[11][1][16] + xor_out[12][1][16] + xor_out[13][1][16] + xor_out[14][1][16];
assign sum_out[3][1][16] = xor_out[15][1][16] + xor_out[16][1][16] + xor_out[17][1][16] + xor_out[18][1][16] + xor_out[19][1][16];
assign sum_out[4][1][16] = xor_out[20][1][16] + xor_out[21][1][16] + xor_out[22][1][16] + xor_out[23][1][16] + xor_out[24][1][16];
assign sum_out[5][1][16] = xor_out[25][1][16] + xor_out[26][1][16] + xor_out[27][1][16] + xor_out[28][1][16] + xor_out[29][1][16];
assign sum_out[6][1][16] = xor_out[30][1][16] + xor_out[31][1][16] + xor_out[32][1][16] + xor_out[33][1][16] + xor_out[34][1][16];
assign sum_out[7][1][16] = xor_out[35][1][16] + xor_out[36][1][16] + xor_out[37][1][16] + xor_out[38][1][16] + xor_out[39][1][16];
assign sum_out[8][1][16] = xor_out[40][1][16] + xor_out[41][1][16] + xor_out[42][1][16] + xor_out[43][1][16] + xor_out[44][1][16];
assign sum_out[9][1][16] = xor_out[45][1][16] + xor_out[46][1][16] + xor_out[47][1][16] + xor_out[48][1][16] + xor_out[49][1][16];
assign sum_out[10][1][16] = xor_out[50][1][16] + xor_out[51][1][16] + xor_out[52][1][16] + xor_out[53][1][16] + xor_out[54][1][16];
assign sum_out[11][1][16] = xor_out[55][1][16] + xor_out[56][1][16] + xor_out[57][1][16] + xor_out[58][1][16] + xor_out[59][1][16];
assign sum_out[12][1][16] = xor_out[60][1][16] + xor_out[61][1][16] + xor_out[62][1][16] + xor_out[63][1][16] + xor_out[64][1][16];
assign sum_out[13][1][16] = xor_out[65][1][16] + xor_out[66][1][16] + xor_out[67][1][16] + xor_out[68][1][16] + xor_out[69][1][16];
assign sum_out[14][1][16] = xor_out[70][1][16] + xor_out[71][1][16] + xor_out[72][1][16] + xor_out[73][1][16] + xor_out[74][1][16];
assign sum_out[15][1][16] = xor_out[75][1][16] + xor_out[76][1][16] + xor_out[77][1][16] + xor_out[78][1][16] + xor_out[79][1][16];
assign sum_out[16][1][16] = xor_out[80][1][16] + xor_out[81][1][16] + xor_out[82][1][16] + xor_out[83][1][16] + xor_out[84][1][16];
assign sum_out[17][1][16] = xor_out[85][1][16] + xor_out[86][1][16] + xor_out[87][1][16] + xor_out[88][1][16] + xor_out[89][1][16];
assign sum_out[18][1][16] = xor_out[90][1][16] + xor_out[91][1][16] + xor_out[92][1][16] + xor_out[93][1][16] + xor_out[94][1][16];
assign sum_out[19][1][16] = xor_out[95][1][16] + xor_out[96][1][16] + xor_out[97][1][16] + xor_out[98][1][16] + xor_out[99][1][16];

assign sum_out[0][1][17] = xor_out[0][1][17] + xor_out[1][1][17] + xor_out[2][1][17] + xor_out[3][1][17] + xor_out[4][1][17];
assign sum_out[1][1][17] = xor_out[5][1][17] + xor_out[6][1][17] + xor_out[7][1][17] + xor_out[8][1][17] + xor_out[9][1][17];
assign sum_out[2][1][17] = xor_out[10][1][17] + xor_out[11][1][17] + xor_out[12][1][17] + xor_out[13][1][17] + xor_out[14][1][17];
assign sum_out[3][1][17] = xor_out[15][1][17] + xor_out[16][1][17] + xor_out[17][1][17] + xor_out[18][1][17] + xor_out[19][1][17];
assign sum_out[4][1][17] = xor_out[20][1][17] + xor_out[21][1][17] + xor_out[22][1][17] + xor_out[23][1][17] + xor_out[24][1][17];
assign sum_out[5][1][17] = xor_out[25][1][17] + xor_out[26][1][17] + xor_out[27][1][17] + xor_out[28][1][17] + xor_out[29][1][17];
assign sum_out[6][1][17] = xor_out[30][1][17] + xor_out[31][1][17] + xor_out[32][1][17] + xor_out[33][1][17] + xor_out[34][1][17];
assign sum_out[7][1][17] = xor_out[35][1][17] + xor_out[36][1][17] + xor_out[37][1][17] + xor_out[38][1][17] + xor_out[39][1][17];
assign sum_out[8][1][17] = xor_out[40][1][17] + xor_out[41][1][17] + xor_out[42][1][17] + xor_out[43][1][17] + xor_out[44][1][17];
assign sum_out[9][1][17] = xor_out[45][1][17] + xor_out[46][1][17] + xor_out[47][1][17] + xor_out[48][1][17] + xor_out[49][1][17];
assign sum_out[10][1][17] = xor_out[50][1][17] + xor_out[51][1][17] + xor_out[52][1][17] + xor_out[53][1][17] + xor_out[54][1][17];
assign sum_out[11][1][17] = xor_out[55][1][17] + xor_out[56][1][17] + xor_out[57][1][17] + xor_out[58][1][17] + xor_out[59][1][17];
assign sum_out[12][1][17] = xor_out[60][1][17] + xor_out[61][1][17] + xor_out[62][1][17] + xor_out[63][1][17] + xor_out[64][1][17];
assign sum_out[13][1][17] = xor_out[65][1][17] + xor_out[66][1][17] + xor_out[67][1][17] + xor_out[68][1][17] + xor_out[69][1][17];
assign sum_out[14][1][17] = xor_out[70][1][17] + xor_out[71][1][17] + xor_out[72][1][17] + xor_out[73][1][17] + xor_out[74][1][17];
assign sum_out[15][1][17] = xor_out[75][1][17] + xor_out[76][1][17] + xor_out[77][1][17] + xor_out[78][1][17] + xor_out[79][1][17];
assign sum_out[16][1][17] = xor_out[80][1][17] + xor_out[81][1][17] + xor_out[82][1][17] + xor_out[83][1][17] + xor_out[84][1][17];
assign sum_out[17][1][17] = xor_out[85][1][17] + xor_out[86][1][17] + xor_out[87][1][17] + xor_out[88][1][17] + xor_out[89][1][17];
assign sum_out[18][1][17] = xor_out[90][1][17] + xor_out[91][1][17] + xor_out[92][1][17] + xor_out[93][1][17] + xor_out[94][1][17];
assign sum_out[19][1][17] = xor_out[95][1][17] + xor_out[96][1][17] + xor_out[97][1][17] + xor_out[98][1][17] + xor_out[99][1][17];

assign sum_out[0][1][18] = xor_out[0][1][18] + xor_out[1][1][18] + xor_out[2][1][18] + xor_out[3][1][18] + xor_out[4][1][18];
assign sum_out[1][1][18] = xor_out[5][1][18] + xor_out[6][1][18] + xor_out[7][1][18] + xor_out[8][1][18] + xor_out[9][1][18];
assign sum_out[2][1][18] = xor_out[10][1][18] + xor_out[11][1][18] + xor_out[12][1][18] + xor_out[13][1][18] + xor_out[14][1][18];
assign sum_out[3][1][18] = xor_out[15][1][18] + xor_out[16][1][18] + xor_out[17][1][18] + xor_out[18][1][18] + xor_out[19][1][18];
assign sum_out[4][1][18] = xor_out[20][1][18] + xor_out[21][1][18] + xor_out[22][1][18] + xor_out[23][1][18] + xor_out[24][1][18];
assign sum_out[5][1][18] = xor_out[25][1][18] + xor_out[26][1][18] + xor_out[27][1][18] + xor_out[28][1][18] + xor_out[29][1][18];
assign sum_out[6][1][18] = xor_out[30][1][18] + xor_out[31][1][18] + xor_out[32][1][18] + xor_out[33][1][18] + xor_out[34][1][18];
assign sum_out[7][1][18] = xor_out[35][1][18] + xor_out[36][1][18] + xor_out[37][1][18] + xor_out[38][1][18] + xor_out[39][1][18];
assign sum_out[8][1][18] = xor_out[40][1][18] + xor_out[41][1][18] + xor_out[42][1][18] + xor_out[43][1][18] + xor_out[44][1][18];
assign sum_out[9][1][18] = xor_out[45][1][18] + xor_out[46][1][18] + xor_out[47][1][18] + xor_out[48][1][18] + xor_out[49][1][18];
assign sum_out[10][1][18] = xor_out[50][1][18] + xor_out[51][1][18] + xor_out[52][1][18] + xor_out[53][1][18] + xor_out[54][1][18];
assign sum_out[11][1][18] = xor_out[55][1][18] + xor_out[56][1][18] + xor_out[57][1][18] + xor_out[58][1][18] + xor_out[59][1][18];
assign sum_out[12][1][18] = xor_out[60][1][18] + xor_out[61][1][18] + xor_out[62][1][18] + xor_out[63][1][18] + xor_out[64][1][18];
assign sum_out[13][1][18] = xor_out[65][1][18] + xor_out[66][1][18] + xor_out[67][1][18] + xor_out[68][1][18] + xor_out[69][1][18];
assign sum_out[14][1][18] = xor_out[70][1][18] + xor_out[71][1][18] + xor_out[72][1][18] + xor_out[73][1][18] + xor_out[74][1][18];
assign sum_out[15][1][18] = xor_out[75][1][18] + xor_out[76][1][18] + xor_out[77][1][18] + xor_out[78][1][18] + xor_out[79][1][18];
assign sum_out[16][1][18] = xor_out[80][1][18] + xor_out[81][1][18] + xor_out[82][1][18] + xor_out[83][1][18] + xor_out[84][1][18];
assign sum_out[17][1][18] = xor_out[85][1][18] + xor_out[86][1][18] + xor_out[87][1][18] + xor_out[88][1][18] + xor_out[89][1][18];
assign sum_out[18][1][18] = xor_out[90][1][18] + xor_out[91][1][18] + xor_out[92][1][18] + xor_out[93][1][18] + xor_out[94][1][18];
assign sum_out[19][1][18] = xor_out[95][1][18] + xor_out[96][1][18] + xor_out[97][1][18] + xor_out[98][1][18] + xor_out[99][1][18];

assign sum_out[0][1][19] = xor_out[0][1][19] + xor_out[1][1][19] + xor_out[2][1][19] + xor_out[3][1][19] + xor_out[4][1][19];
assign sum_out[1][1][19] = xor_out[5][1][19] + xor_out[6][1][19] + xor_out[7][1][19] + xor_out[8][1][19] + xor_out[9][1][19];
assign sum_out[2][1][19] = xor_out[10][1][19] + xor_out[11][1][19] + xor_out[12][1][19] + xor_out[13][1][19] + xor_out[14][1][19];
assign sum_out[3][1][19] = xor_out[15][1][19] + xor_out[16][1][19] + xor_out[17][1][19] + xor_out[18][1][19] + xor_out[19][1][19];
assign sum_out[4][1][19] = xor_out[20][1][19] + xor_out[21][1][19] + xor_out[22][1][19] + xor_out[23][1][19] + xor_out[24][1][19];
assign sum_out[5][1][19] = xor_out[25][1][19] + xor_out[26][1][19] + xor_out[27][1][19] + xor_out[28][1][19] + xor_out[29][1][19];
assign sum_out[6][1][19] = xor_out[30][1][19] + xor_out[31][1][19] + xor_out[32][1][19] + xor_out[33][1][19] + xor_out[34][1][19];
assign sum_out[7][1][19] = xor_out[35][1][19] + xor_out[36][1][19] + xor_out[37][1][19] + xor_out[38][1][19] + xor_out[39][1][19];
assign sum_out[8][1][19] = xor_out[40][1][19] + xor_out[41][1][19] + xor_out[42][1][19] + xor_out[43][1][19] + xor_out[44][1][19];
assign sum_out[9][1][19] = xor_out[45][1][19] + xor_out[46][1][19] + xor_out[47][1][19] + xor_out[48][1][19] + xor_out[49][1][19];
assign sum_out[10][1][19] = xor_out[50][1][19] + xor_out[51][1][19] + xor_out[52][1][19] + xor_out[53][1][19] + xor_out[54][1][19];
assign sum_out[11][1][19] = xor_out[55][1][19] + xor_out[56][1][19] + xor_out[57][1][19] + xor_out[58][1][19] + xor_out[59][1][19];
assign sum_out[12][1][19] = xor_out[60][1][19] + xor_out[61][1][19] + xor_out[62][1][19] + xor_out[63][1][19] + xor_out[64][1][19];
assign sum_out[13][1][19] = xor_out[65][1][19] + xor_out[66][1][19] + xor_out[67][1][19] + xor_out[68][1][19] + xor_out[69][1][19];
assign sum_out[14][1][19] = xor_out[70][1][19] + xor_out[71][1][19] + xor_out[72][1][19] + xor_out[73][1][19] + xor_out[74][1][19];
assign sum_out[15][1][19] = xor_out[75][1][19] + xor_out[76][1][19] + xor_out[77][1][19] + xor_out[78][1][19] + xor_out[79][1][19];
assign sum_out[16][1][19] = xor_out[80][1][19] + xor_out[81][1][19] + xor_out[82][1][19] + xor_out[83][1][19] + xor_out[84][1][19];
assign sum_out[17][1][19] = xor_out[85][1][19] + xor_out[86][1][19] + xor_out[87][1][19] + xor_out[88][1][19] + xor_out[89][1][19];
assign sum_out[18][1][19] = xor_out[90][1][19] + xor_out[91][1][19] + xor_out[92][1][19] + xor_out[93][1][19] + xor_out[94][1][19];
assign sum_out[19][1][19] = xor_out[95][1][19] + xor_out[96][1][19] + xor_out[97][1][19] + xor_out[98][1][19] + xor_out[99][1][19];

assign sum_out[0][1][20] = xor_out[0][1][20] + xor_out[1][1][20] + xor_out[2][1][20] + xor_out[3][1][20] + xor_out[4][1][20];
assign sum_out[1][1][20] = xor_out[5][1][20] + xor_out[6][1][20] + xor_out[7][1][20] + xor_out[8][1][20] + xor_out[9][1][20];
assign sum_out[2][1][20] = xor_out[10][1][20] + xor_out[11][1][20] + xor_out[12][1][20] + xor_out[13][1][20] + xor_out[14][1][20];
assign sum_out[3][1][20] = xor_out[15][1][20] + xor_out[16][1][20] + xor_out[17][1][20] + xor_out[18][1][20] + xor_out[19][1][20];
assign sum_out[4][1][20] = xor_out[20][1][20] + xor_out[21][1][20] + xor_out[22][1][20] + xor_out[23][1][20] + xor_out[24][1][20];
assign sum_out[5][1][20] = xor_out[25][1][20] + xor_out[26][1][20] + xor_out[27][1][20] + xor_out[28][1][20] + xor_out[29][1][20];
assign sum_out[6][1][20] = xor_out[30][1][20] + xor_out[31][1][20] + xor_out[32][1][20] + xor_out[33][1][20] + xor_out[34][1][20];
assign sum_out[7][1][20] = xor_out[35][1][20] + xor_out[36][1][20] + xor_out[37][1][20] + xor_out[38][1][20] + xor_out[39][1][20];
assign sum_out[8][1][20] = xor_out[40][1][20] + xor_out[41][1][20] + xor_out[42][1][20] + xor_out[43][1][20] + xor_out[44][1][20];
assign sum_out[9][1][20] = xor_out[45][1][20] + xor_out[46][1][20] + xor_out[47][1][20] + xor_out[48][1][20] + xor_out[49][1][20];
assign sum_out[10][1][20] = xor_out[50][1][20] + xor_out[51][1][20] + xor_out[52][1][20] + xor_out[53][1][20] + xor_out[54][1][20];
assign sum_out[11][1][20] = xor_out[55][1][20] + xor_out[56][1][20] + xor_out[57][1][20] + xor_out[58][1][20] + xor_out[59][1][20];
assign sum_out[12][1][20] = xor_out[60][1][20] + xor_out[61][1][20] + xor_out[62][1][20] + xor_out[63][1][20] + xor_out[64][1][20];
assign sum_out[13][1][20] = xor_out[65][1][20] + xor_out[66][1][20] + xor_out[67][1][20] + xor_out[68][1][20] + xor_out[69][1][20];
assign sum_out[14][1][20] = xor_out[70][1][20] + xor_out[71][1][20] + xor_out[72][1][20] + xor_out[73][1][20] + xor_out[74][1][20];
assign sum_out[15][1][20] = xor_out[75][1][20] + xor_out[76][1][20] + xor_out[77][1][20] + xor_out[78][1][20] + xor_out[79][1][20];
assign sum_out[16][1][20] = xor_out[80][1][20] + xor_out[81][1][20] + xor_out[82][1][20] + xor_out[83][1][20] + xor_out[84][1][20];
assign sum_out[17][1][20] = xor_out[85][1][20] + xor_out[86][1][20] + xor_out[87][1][20] + xor_out[88][1][20] + xor_out[89][1][20];
assign sum_out[18][1][20] = xor_out[90][1][20] + xor_out[91][1][20] + xor_out[92][1][20] + xor_out[93][1][20] + xor_out[94][1][20];
assign sum_out[19][1][20] = xor_out[95][1][20] + xor_out[96][1][20] + xor_out[97][1][20] + xor_out[98][1][20] + xor_out[99][1][20];

assign sum_out[0][1][21] = xor_out[0][1][21] + xor_out[1][1][21] + xor_out[2][1][21] + xor_out[3][1][21] + xor_out[4][1][21];
assign sum_out[1][1][21] = xor_out[5][1][21] + xor_out[6][1][21] + xor_out[7][1][21] + xor_out[8][1][21] + xor_out[9][1][21];
assign sum_out[2][1][21] = xor_out[10][1][21] + xor_out[11][1][21] + xor_out[12][1][21] + xor_out[13][1][21] + xor_out[14][1][21];
assign sum_out[3][1][21] = xor_out[15][1][21] + xor_out[16][1][21] + xor_out[17][1][21] + xor_out[18][1][21] + xor_out[19][1][21];
assign sum_out[4][1][21] = xor_out[20][1][21] + xor_out[21][1][21] + xor_out[22][1][21] + xor_out[23][1][21] + xor_out[24][1][21];
assign sum_out[5][1][21] = xor_out[25][1][21] + xor_out[26][1][21] + xor_out[27][1][21] + xor_out[28][1][21] + xor_out[29][1][21];
assign sum_out[6][1][21] = xor_out[30][1][21] + xor_out[31][1][21] + xor_out[32][1][21] + xor_out[33][1][21] + xor_out[34][1][21];
assign sum_out[7][1][21] = xor_out[35][1][21] + xor_out[36][1][21] + xor_out[37][1][21] + xor_out[38][1][21] + xor_out[39][1][21];
assign sum_out[8][1][21] = xor_out[40][1][21] + xor_out[41][1][21] + xor_out[42][1][21] + xor_out[43][1][21] + xor_out[44][1][21];
assign sum_out[9][1][21] = xor_out[45][1][21] + xor_out[46][1][21] + xor_out[47][1][21] + xor_out[48][1][21] + xor_out[49][1][21];
assign sum_out[10][1][21] = xor_out[50][1][21] + xor_out[51][1][21] + xor_out[52][1][21] + xor_out[53][1][21] + xor_out[54][1][21];
assign sum_out[11][1][21] = xor_out[55][1][21] + xor_out[56][1][21] + xor_out[57][1][21] + xor_out[58][1][21] + xor_out[59][1][21];
assign sum_out[12][1][21] = xor_out[60][1][21] + xor_out[61][1][21] + xor_out[62][1][21] + xor_out[63][1][21] + xor_out[64][1][21];
assign sum_out[13][1][21] = xor_out[65][1][21] + xor_out[66][1][21] + xor_out[67][1][21] + xor_out[68][1][21] + xor_out[69][1][21];
assign sum_out[14][1][21] = xor_out[70][1][21] + xor_out[71][1][21] + xor_out[72][1][21] + xor_out[73][1][21] + xor_out[74][1][21];
assign sum_out[15][1][21] = xor_out[75][1][21] + xor_out[76][1][21] + xor_out[77][1][21] + xor_out[78][1][21] + xor_out[79][1][21];
assign sum_out[16][1][21] = xor_out[80][1][21] + xor_out[81][1][21] + xor_out[82][1][21] + xor_out[83][1][21] + xor_out[84][1][21];
assign sum_out[17][1][21] = xor_out[85][1][21] + xor_out[86][1][21] + xor_out[87][1][21] + xor_out[88][1][21] + xor_out[89][1][21];
assign sum_out[18][1][21] = xor_out[90][1][21] + xor_out[91][1][21] + xor_out[92][1][21] + xor_out[93][1][21] + xor_out[94][1][21];
assign sum_out[19][1][21] = xor_out[95][1][21] + xor_out[96][1][21] + xor_out[97][1][21] + xor_out[98][1][21] + xor_out[99][1][21];

assign sum_out[0][1][22] = xor_out[0][1][22] + xor_out[1][1][22] + xor_out[2][1][22] + xor_out[3][1][22] + xor_out[4][1][22];
assign sum_out[1][1][22] = xor_out[5][1][22] + xor_out[6][1][22] + xor_out[7][1][22] + xor_out[8][1][22] + xor_out[9][1][22];
assign sum_out[2][1][22] = xor_out[10][1][22] + xor_out[11][1][22] + xor_out[12][1][22] + xor_out[13][1][22] + xor_out[14][1][22];
assign sum_out[3][1][22] = xor_out[15][1][22] + xor_out[16][1][22] + xor_out[17][1][22] + xor_out[18][1][22] + xor_out[19][1][22];
assign sum_out[4][1][22] = xor_out[20][1][22] + xor_out[21][1][22] + xor_out[22][1][22] + xor_out[23][1][22] + xor_out[24][1][22];
assign sum_out[5][1][22] = xor_out[25][1][22] + xor_out[26][1][22] + xor_out[27][1][22] + xor_out[28][1][22] + xor_out[29][1][22];
assign sum_out[6][1][22] = xor_out[30][1][22] + xor_out[31][1][22] + xor_out[32][1][22] + xor_out[33][1][22] + xor_out[34][1][22];
assign sum_out[7][1][22] = xor_out[35][1][22] + xor_out[36][1][22] + xor_out[37][1][22] + xor_out[38][1][22] + xor_out[39][1][22];
assign sum_out[8][1][22] = xor_out[40][1][22] + xor_out[41][1][22] + xor_out[42][1][22] + xor_out[43][1][22] + xor_out[44][1][22];
assign sum_out[9][1][22] = xor_out[45][1][22] + xor_out[46][1][22] + xor_out[47][1][22] + xor_out[48][1][22] + xor_out[49][1][22];
assign sum_out[10][1][22] = xor_out[50][1][22] + xor_out[51][1][22] + xor_out[52][1][22] + xor_out[53][1][22] + xor_out[54][1][22];
assign sum_out[11][1][22] = xor_out[55][1][22] + xor_out[56][1][22] + xor_out[57][1][22] + xor_out[58][1][22] + xor_out[59][1][22];
assign sum_out[12][1][22] = xor_out[60][1][22] + xor_out[61][1][22] + xor_out[62][1][22] + xor_out[63][1][22] + xor_out[64][1][22];
assign sum_out[13][1][22] = xor_out[65][1][22] + xor_out[66][1][22] + xor_out[67][1][22] + xor_out[68][1][22] + xor_out[69][1][22];
assign sum_out[14][1][22] = xor_out[70][1][22] + xor_out[71][1][22] + xor_out[72][1][22] + xor_out[73][1][22] + xor_out[74][1][22];
assign sum_out[15][1][22] = xor_out[75][1][22] + xor_out[76][1][22] + xor_out[77][1][22] + xor_out[78][1][22] + xor_out[79][1][22];
assign sum_out[16][1][22] = xor_out[80][1][22] + xor_out[81][1][22] + xor_out[82][1][22] + xor_out[83][1][22] + xor_out[84][1][22];
assign sum_out[17][1][22] = xor_out[85][1][22] + xor_out[86][1][22] + xor_out[87][1][22] + xor_out[88][1][22] + xor_out[89][1][22];
assign sum_out[18][1][22] = xor_out[90][1][22] + xor_out[91][1][22] + xor_out[92][1][22] + xor_out[93][1][22] + xor_out[94][1][22];
assign sum_out[19][1][22] = xor_out[95][1][22] + xor_out[96][1][22] + xor_out[97][1][22] + xor_out[98][1][22] + xor_out[99][1][22];

assign sum_out[0][1][23] = xor_out[0][1][23] + xor_out[1][1][23] + xor_out[2][1][23] + xor_out[3][1][23] + xor_out[4][1][23];
assign sum_out[1][1][23] = xor_out[5][1][23] + xor_out[6][1][23] + xor_out[7][1][23] + xor_out[8][1][23] + xor_out[9][1][23];
assign sum_out[2][1][23] = xor_out[10][1][23] + xor_out[11][1][23] + xor_out[12][1][23] + xor_out[13][1][23] + xor_out[14][1][23];
assign sum_out[3][1][23] = xor_out[15][1][23] + xor_out[16][1][23] + xor_out[17][1][23] + xor_out[18][1][23] + xor_out[19][1][23];
assign sum_out[4][1][23] = xor_out[20][1][23] + xor_out[21][1][23] + xor_out[22][1][23] + xor_out[23][1][23] + xor_out[24][1][23];
assign sum_out[5][1][23] = xor_out[25][1][23] + xor_out[26][1][23] + xor_out[27][1][23] + xor_out[28][1][23] + xor_out[29][1][23];
assign sum_out[6][1][23] = xor_out[30][1][23] + xor_out[31][1][23] + xor_out[32][1][23] + xor_out[33][1][23] + xor_out[34][1][23];
assign sum_out[7][1][23] = xor_out[35][1][23] + xor_out[36][1][23] + xor_out[37][1][23] + xor_out[38][1][23] + xor_out[39][1][23];
assign sum_out[8][1][23] = xor_out[40][1][23] + xor_out[41][1][23] + xor_out[42][1][23] + xor_out[43][1][23] + xor_out[44][1][23];
assign sum_out[9][1][23] = xor_out[45][1][23] + xor_out[46][1][23] + xor_out[47][1][23] + xor_out[48][1][23] + xor_out[49][1][23];
assign sum_out[10][1][23] = xor_out[50][1][23] + xor_out[51][1][23] + xor_out[52][1][23] + xor_out[53][1][23] + xor_out[54][1][23];
assign sum_out[11][1][23] = xor_out[55][1][23] + xor_out[56][1][23] + xor_out[57][1][23] + xor_out[58][1][23] + xor_out[59][1][23];
assign sum_out[12][1][23] = xor_out[60][1][23] + xor_out[61][1][23] + xor_out[62][1][23] + xor_out[63][1][23] + xor_out[64][1][23];
assign sum_out[13][1][23] = xor_out[65][1][23] + xor_out[66][1][23] + xor_out[67][1][23] + xor_out[68][1][23] + xor_out[69][1][23];
assign sum_out[14][1][23] = xor_out[70][1][23] + xor_out[71][1][23] + xor_out[72][1][23] + xor_out[73][1][23] + xor_out[74][1][23];
assign sum_out[15][1][23] = xor_out[75][1][23] + xor_out[76][1][23] + xor_out[77][1][23] + xor_out[78][1][23] + xor_out[79][1][23];
assign sum_out[16][1][23] = xor_out[80][1][23] + xor_out[81][1][23] + xor_out[82][1][23] + xor_out[83][1][23] + xor_out[84][1][23];
assign sum_out[17][1][23] = xor_out[85][1][23] + xor_out[86][1][23] + xor_out[87][1][23] + xor_out[88][1][23] + xor_out[89][1][23];
assign sum_out[18][1][23] = xor_out[90][1][23] + xor_out[91][1][23] + xor_out[92][1][23] + xor_out[93][1][23] + xor_out[94][1][23];
assign sum_out[19][1][23] = xor_out[95][1][23] + xor_out[96][1][23] + xor_out[97][1][23] + xor_out[98][1][23] + xor_out[99][1][23];

assign sum_out[0][2][0] = xor_out[0][2][0] + xor_out[1][2][0] + xor_out[2][2][0] + xor_out[3][2][0] + xor_out[4][2][0];
assign sum_out[1][2][0] = xor_out[5][2][0] + xor_out[6][2][0] + xor_out[7][2][0] + xor_out[8][2][0] + xor_out[9][2][0];
assign sum_out[2][2][0] = xor_out[10][2][0] + xor_out[11][2][0] + xor_out[12][2][0] + xor_out[13][2][0] + xor_out[14][2][0];
assign sum_out[3][2][0] = xor_out[15][2][0] + xor_out[16][2][0] + xor_out[17][2][0] + xor_out[18][2][0] + xor_out[19][2][0];
assign sum_out[4][2][0] = xor_out[20][2][0] + xor_out[21][2][0] + xor_out[22][2][0] + xor_out[23][2][0] + xor_out[24][2][0];
assign sum_out[5][2][0] = xor_out[25][2][0] + xor_out[26][2][0] + xor_out[27][2][0] + xor_out[28][2][0] + xor_out[29][2][0];
assign sum_out[6][2][0] = xor_out[30][2][0] + xor_out[31][2][0] + xor_out[32][2][0] + xor_out[33][2][0] + xor_out[34][2][0];
assign sum_out[7][2][0] = xor_out[35][2][0] + xor_out[36][2][0] + xor_out[37][2][0] + xor_out[38][2][0] + xor_out[39][2][0];
assign sum_out[8][2][0] = xor_out[40][2][0] + xor_out[41][2][0] + xor_out[42][2][0] + xor_out[43][2][0] + xor_out[44][2][0];
assign sum_out[9][2][0] = xor_out[45][2][0] + xor_out[46][2][0] + xor_out[47][2][0] + xor_out[48][2][0] + xor_out[49][2][0];
assign sum_out[10][2][0] = xor_out[50][2][0] + xor_out[51][2][0] + xor_out[52][2][0] + xor_out[53][2][0] + xor_out[54][2][0];
assign sum_out[11][2][0] = xor_out[55][2][0] + xor_out[56][2][0] + xor_out[57][2][0] + xor_out[58][2][0] + xor_out[59][2][0];
assign sum_out[12][2][0] = xor_out[60][2][0] + xor_out[61][2][0] + xor_out[62][2][0] + xor_out[63][2][0] + xor_out[64][2][0];
assign sum_out[13][2][0] = xor_out[65][2][0] + xor_out[66][2][0] + xor_out[67][2][0] + xor_out[68][2][0] + xor_out[69][2][0];
assign sum_out[14][2][0] = xor_out[70][2][0] + xor_out[71][2][0] + xor_out[72][2][0] + xor_out[73][2][0] + xor_out[74][2][0];
assign sum_out[15][2][0] = xor_out[75][2][0] + xor_out[76][2][0] + xor_out[77][2][0] + xor_out[78][2][0] + xor_out[79][2][0];
assign sum_out[16][2][0] = xor_out[80][2][0] + xor_out[81][2][0] + xor_out[82][2][0] + xor_out[83][2][0] + xor_out[84][2][0];
assign sum_out[17][2][0] = xor_out[85][2][0] + xor_out[86][2][0] + xor_out[87][2][0] + xor_out[88][2][0] + xor_out[89][2][0];
assign sum_out[18][2][0] = xor_out[90][2][0] + xor_out[91][2][0] + xor_out[92][2][0] + xor_out[93][2][0] + xor_out[94][2][0];
assign sum_out[19][2][0] = xor_out[95][2][0] + xor_out[96][2][0] + xor_out[97][2][0] + xor_out[98][2][0] + xor_out[99][2][0];

assign sum_out[0][2][1] = xor_out[0][2][1] + xor_out[1][2][1] + xor_out[2][2][1] + xor_out[3][2][1] + xor_out[4][2][1];
assign sum_out[1][2][1] = xor_out[5][2][1] + xor_out[6][2][1] + xor_out[7][2][1] + xor_out[8][2][1] + xor_out[9][2][1];
assign sum_out[2][2][1] = xor_out[10][2][1] + xor_out[11][2][1] + xor_out[12][2][1] + xor_out[13][2][1] + xor_out[14][2][1];
assign sum_out[3][2][1] = xor_out[15][2][1] + xor_out[16][2][1] + xor_out[17][2][1] + xor_out[18][2][1] + xor_out[19][2][1];
assign sum_out[4][2][1] = xor_out[20][2][1] + xor_out[21][2][1] + xor_out[22][2][1] + xor_out[23][2][1] + xor_out[24][2][1];
assign sum_out[5][2][1] = xor_out[25][2][1] + xor_out[26][2][1] + xor_out[27][2][1] + xor_out[28][2][1] + xor_out[29][2][1];
assign sum_out[6][2][1] = xor_out[30][2][1] + xor_out[31][2][1] + xor_out[32][2][1] + xor_out[33][2][1] + xor_out[34][2][1];
assign sum_out[7][2][1] = xor_out[35][2][1] + xor_out[36][2][1] + xor_out[37][2][1] + xor_out[38][2][1] + xor_out[39][2][1];
assign sum_out[8][2][1] = xor_out[40][2][1] + xor_out[41][2][1] + xor_out[42][2][1] + xor_out[43][2][1] + xor_out[44][2][1];
assign sum_out[9][2][1] = xor_out[45][2][1] + xor_out[46][2][1] + xor_out[47][2][1] + xor_out[48][2][1] + xor_out[49][2][1];
assign sum_out[10][2][1] = xor_out[50][2][1] + xor_out[51][2][1] + xor_out[52][2][1] + xor_out[53][2][1] + xor_out[54][2][1];
assign sum_out[11][2][1] = xor_out[55][2][1] + xor_out[56][2][1] + xor_out[57][2][1] + xor_out[58][2][1] + xor_out[59][2][1];
assign sum_out[12][2][1] = xor_out[60][2][1] + xor_out[61][2][1] + xor_out[62][2][1] + xor_out[63][2][1] + xor_out[64][2][1];
assign sum_out[13][2][1] = xor_out[65][2][1] + xor_out[66][2][1] + xor_out[67][2][1] + xor_out[68][2][1] + xor_out[69][2][1];
assign sum_out[14][2][1] = xor_out[70][2][1] + xor_out[71][2][1] + xor_out[72][2][1] + xor_out[73][2][1] + xor_out[74][2][1];
assign sum_out[15][2][1] = xor_out[75][2][1] + xor_out[76][2][1] + xor_out[77][2][1] + xor_out[78][2][1] + xor_out[79][2][1];
assign sum_out[16][2][1] = xor_out[80][2][1] + xor_out[81][2][1] + xor_out[82][2][1] + xor_out[83][2][1] + xor_out[84][2][1];
assign sum_out[17][2][1] = xor_out[85][2][1] + xor_out[86][2][1] + xor_out[87][2][1] + xor_out[88][2][1] + xor_out[89][2][1];
assign sum_out[18][2][1] = xor_out[90][2][1] + xor_out[91][2][1] + xor_out[92][2][1] + xor_out[93][2][1] + xor_out[94][2][1];
assign sum_out[19][2][1] = xor_out[95][2][1] + xor_out[96][2][1] + xor_out[97][2][1] + xor_out[98][2][1] + xor_out[99][2][1];

assign sum_out[0][2][2] = xor_out[0][2][2] + xor_out[1][2][2] + xor_out[2][2][2] + xor_out[3][2][2] + xor_out[4][2][2];
assign sum_out[1][2][2] = xor_out[5][2][2] + xor_out[6][2][2] + xor_out[7][2][2] + xor_out[8][2][2] + xor_out[9][2][2];
assign sum_out[2][2][2] = xor_out[10][2][2] + xor_out[11][2][2] + xor_out[12][2][2] + xor_out[13][2][2] + xor_out[14][2][2];
assign sum_out[3][2][2] = xor_out[15][2][2] + xor_out[16][2][2] + xor_out[17][2][2] + xor_out[18][2][2] + xor_out[19][2][2];
assign sum_out[4][2][2] = xor_out[20][2][2] + xor_out[21][2][2] + xor_out[22][2][2] + xor_out[23][2][2] + xor_out[24][2][2];
assign sum_out[5][2][2] = xor_out[25][2][2] + xor_out[26][2][2] + xor_out[27][2][2] + xor_out[28][2][2] + xor_out[29][2][2];
assign sum_out[6][2][2] = xor_out[30][2][2] + xor_out[31][2][2] + xor_out[32][2][2] + xor_out[33][2][2] + xor_out[34][2][2];
assign sum_out[7][2][2] = xor_out[35][2][2] + xor_out[36][2][2] + xor_out[37][2][2] + xor_out[38][2][2] + xor_out[39][2][2];
assign sum_out[8][2][2] = xor_out[40][2][2] + xor_out[41][2][2] + xor_out[42][2][2] + xor_out[43][2][2] + xor_out[44][2][2];
assign sum_out[9][2][2] = xor_out[45][2][2] + xor_out[46][2][2] + xor_out[47][2][2] + xor_out[48][2][2] + xor_out[49][2][2];
assign sum_out[10][2][2] = xor_out[50][2][2] + xor_out[51][2][2] + xor_out[52][2][2] + xor_out[53][2][2] + xor_out[54][2][2];
assign sum_out[11][2][2] = xor_out[55][2][2] + xor_out[56][2][2] + xor_out[57][2][2] + xor_out[58][2][2] + xor_out[59][2][2];
assign sum_out[12][2][2] = xor_out[60][2][2] + xor_out[61][2][2] + xor_out[62][2][2] + xor_out[63][2][2] + xor_out[64][2][2];
assign sum_out[13][2][2] = xor_out[65][2][2] + xor_out[66][2][2] + xor_out[67][2][2] + xor_out[68][2][2] + xor_out[69][2][2];
assign sum_out[14][2][2] = xor_out[70][2][2] + xor_out[71][2][2] + xor_out[72][2][2] + xor_out[73][2][2] + xor_out[74][2][2];
assign sum_out[15][2][2] = xor_out[75][2][2] + xor_out[76][2][2] + xor_out[77][2][2] + xor_out[78][2][2] + xor_out[79][2][2];
assign sum_out[16][2][2] = xor_out[80][2][2] + xor_out[81][2][2] + xor_out[82][2][2] + xor_out[83][2][2] + xor_out[84][2][2];
assign sum_out[17][2][2] = xor_out[85][2][2] + xor_out[86][2][2] + xor_out[87][2][2] + xor_out[88][2][2] + xor_out[89][2][2];
assign sum_out[18][2][2] = xor_out[90][2][2] + xor_out[91][2][2] + xor_out[92][2][2] + xor_out[93][2][2] + xor_out[94][2][2];
assign sum_out[19][2][2] = xor_out[95][2][2] + xor_out[96][2][2] + xor_out[97][2][2] + xor_out[98][2][2] + xor_out[99][2][2];

assign sum_out[0][2][3] = xor_out[0][2][3] + xor_out[1][2][3] + xor_out[2][2][3] + xor_out[3][2][3] + xor_out[4][2][3];
assign sum_out[1][2][3] = xor_out[5][2][3] + xor_out[6][2][3] + xor_out[7][2][3] + xor_out[8][2][3] + xor_out[9][2][3];
assign sum_out[2][2][3] = xor_out[10][2][3] + xor_out[11][2][3] + xor_out[12][2][3] + xor_out[13][2][3] + xor_out[14][2][3];
assign sum_out[3][2][3] = xor_out[15][2][3] + xor_out[16][2][3] + xor_out[17][2][3] + xor_out[18][2][3] + xor_out[19][2][3];
assign sum_out[4][2][3] = xor_out[20][2][3] + xor_out[21][2][3] + xor_out[22][2][3] + xor_out[23][2][3] + xor_out[24][2][3];
assign sum_out[5][2][3] = xor_out[25][2][3] + xor_out[26][2][3] + xor_out[27][2][3] + xor_out[28][2][3] + xor_out[29][2][3];
assign sum_out[6][2][3] = xor_out[30][2][3] + xor_out[31][2][3] + xor_out[32][2][3] + xor_out[33][2][3] + xor_out[34][2][3];
assign sum_out[7][2][3] = xor_out[35][2][3] + xor_out[36][2][3] + xor_out[37][2][3] + xor_out[38][2][3] + xor_out[39][2][3];
assign sum_out[8][2][3] = xor_out[40][2][3] + xor_out[41][2][3] + xor_out[42][2][3] + xor_out[43][2][3] + xor_out[44][2][3];
assign sum_out[9][2][3] = xor_out[45][2][3] + xor_out[46][2][3] + xor_out[47][2][3] + xor_out[48][2][3] + xor_out[49][2][3];
assign sum_out[10][2][3] = xor_out[50][2][3] + xor_out[51][2][3] + xor_out[52][2][3] + xor_out[53][2][3] + xor_out[54][2][3];
assign sum_out[11][2][3] = xor_out[55][2][3] + xor_out[56][2][3] + xor_out[57][2][3] + xor_out[58][2][3] + xor_out[59][2][3];
assign sum_out[12][2][3] = xor_out[60][2][3] + xor_out[61][2][3] + xor_out[62][2][3] + xor_out[63][2][3] + xor_out[64][2][3];
assign sum_out[13][2][3] = xor_out[65][2][3] + xor_out[66][2][3] + xor_out[67][2][3] + xor_out[68][2][3] + xor_out[69][2][3];
assign sum_out[14][2][3] = xor_out[70][2][3] + xor_out[71][2][3] + xor_out[72][2][3] + xor_out[73][2][3] + xor_out[74][2][3];
assign sum_out[15][2][3] = xor_out[75][2][3] + xor_out[76][2][3] + xor_out[77][2][3] + xor_out[78][2][3] + xor_out[79][2][3];
assign sum_out[16][2][3] = xor_out[80][2][3] + xor_out[81][2][3] + xor_out[82][2][3] + xor_out[83][2][3] + xor_out[84][2][3];
assign sum_out[17][2][3] = xor_out[85][2][3] + xor_out[86][2][3] + xor_out[87][2][3] + xor_out[88][2][3] + xor_out[89][2][3];
assign sum_out[18][2][3] = xor_out[90][2][3] + xor_out[91][2][3] + xor_out[92][2][3] + xor_out[93][2][3] + xor_out[94][2][3];
assign sum_out[19][2][3] = xor_out[95][2][3] + xor_out[96][2][3] + xor_out[97][2][3] + xor_out[98][2][3] + xor_out[99][2][3];

assign sum_out[0][2][4] = xor_out[0][2][4] + xor_out[1][2][4] + xor_out[2][2][4] + xor_out[3][2][4] + xor_out[4][2][4];
assign sum_out[1][2][4] = xor_out[5][2][4] + xor_out[6][2][4] + xor_out[7][2][4] + xor_out[8][2][4] + xor_out[9][2][4];
assign sum_out[2][2][4] = xor_out[10][2][4] + xor_out[11][2][4] + xor_out[12][2][4] + xor_out[13][2][4] + xor_out[14][2][4];
assign sum_out[3][2][4] = xor_out[15][2][4] + xor_out[16][2][4] + xor_out[17][2][4] + xor_out[18][2][4] + xor_out[19][2][4];
assign sum_out[4][2][4] = xor_out[20][2][4] + xor_out[21][2][4] + xor_out[22][2][4] + xor_out[23][2][4] + xor_out[24][2][4];
assign sum_out[5][2][4] = xor_out[25][2][4] + xor_out[26][2][4] + xor_out[27][2][4] + xor_out[28][2][4] + xor_out[29][2][4];
assign sum_out[6][2][4] = xor_out[30][2][4] + xor_out[31][2][4] + xor_out[32][2][4] + xor_out[33][2][4] + xor_out[34][2][4];
assign sum_out[7][2][4] = xor_out[35][2][4] + xor_out[36][2][4] + xor_out[37][2][4] + xor_out[38][2][4] + xor_out[39][2][4];
assign sum_out[8][2][4] = xor_out[40][2][4] + xor_out[41][2][4] + xor_out[42][2][4] + xor_out[43][2][4] + xor_out[44][2][4];
assign sum_out[9][2][4] = xor_out[45][2][4] + xor_out[46][2][4] + xor_out[47][2][4] + xor_out[48][2][4] + xor_out[49][2][4];
assign sum_out[10][2][4] = xor_out[50][2][4] + xor_out[51][2][4] + xor_out[52][2][4] + xor_out[53][2][4] + xor_out[54][2][4];
assign sum_out[11][2][4] = xor_out[55][2][4] + xor_out[56][2][4] + xor_out[57][2][4] + xor_out[58][2][4] + xor_out[59][2][4];
assign sum_out[12][2][4] = xor_out[60][2][4] + xor_out[61][2][4] + xor_out[62][2][4] + xor_out[63][2][4] + xor_out[64][2][4];
assign sum_out[13][2][4] = xor_out[65][2][4] + xor_out[66][2][4] + xor_out[67][2][4] + xor_out[68][2][4] + xor_out[69][2][4];
assign sum_out[14][2][4] = xor_out[70][2][4] + xor_out[71][2][4] + xor_out[72][2][4] + xor_out[73][2][4] + xor_out[74][2][4];
assign sum_out[15][2][4] = xor_out[75][2][4] + xor_out[76][2][4] + xor_out[77][2][4] + xor_out[78][2][4] + xor_out[79][2][4];
assign sum_out[16][2][4] = xor_out[80][2][4] + xor_out[81][2][4] + xor_out[82][2][4] + xor_out[83][2][4] + xor_out[84][2][4];
assign sum_out[17][2][4] = xor_out[85][2][4] + xor_out[86][2][4] + xor_out[87][2][4] + xor_out[88][2][4] + xor_out[89][2][4];
assign sum_out[18][2][4] = xor_out[90][2][4] + xor_out[91][2][4] + xor_out[92][2][4] + xor_out[93][2][4] + xor_out[94][2][4];
assign sum_out[19][2][4] = xor_out[95][2][4] + xor_out[96][2][4] + xor_out[97][2][4] + xor_out[98][2][4] + xor_out[99][2][4];

assign sum_out[0][2][5] = xor_out[0][2][5] + xor_out[1][2][5] + xor_out[2][2][5] + xor_out[3][2][5] + xor_out[4][2][5];
assign sum_out[1][2][5] = xor_out[5][2][5] + xor_out[6][2][5] + xor_out[7][2][5] + xor_out[8][2][5] + xor_out[9][2][5];
assign sum_out[2][2][5] = xor_out[10][2][5] + xor_out[11][2][5] + xor_out[12][2][5] + xor_out[13][2][5] + xor_out[14][2][5];
assign sum_out[3][2][5] = xor_out[15][2][5] + xor_out[16][2][5] + xor_out[17][2][5] + xor_out[18][2][5] + xor_out[19][2][5];
assign sum_out[4][2][5] = xor_out[20][2][5] + xor_out[21][2][5] + xor_out[22][2][5] + xor_out[23][2][5] + xor_out[24][2][5];
assign sum_out[5][2][5] = xor_out[25][2][5] + xor_out[26][2][5] + xor_out[27][2][5] + xor_out[28][2][5] + xor_out[29][2][5];
assign sum_out[6][2][5] = xor_out[30][2][5] + xor_out[31][2][5] + xor_out[32][2][5] + xor_out[33][2][5] + xor_out[34][2][5];
assign sum_out[7][2][5] = xor_out[35][2][5] + xor_out[36][2][5] + xor_out[37][2][5] + xor_out[38][2][5] + xor_out[39][2][5];
assign sum_out[8][2][5] = xor_out[40][2][5] + xor_out[41][2][5] + xor_out[42][2][5] + xor_out[43][2][5] + xor_out[44][2][5];
assign sum_out[9][2][5] = xor_out[45][2][5] + xor_out[46][2][5] + xor_out[47][2][5] + xor_out[48][2][5] + xor_out[49][2][5];
assign sum_out[10][2][5] = xor_out[50][2][5] + xor_out[51][2][5] + xor_out[52][2][5] + xor_out[53][2][5] + xor_out[54][2][5];
assign sum_out[11][2][5] = xor_out[55][2][5] + xor_out[56][2][5] + xor_out[57][2][5] + xor_out[58][2][5] + xor_out[59][2][5];
assign sum_out[12][2][5] = xor_out[60][2][5] + xor_out[61][2][5] + xor_out[62][2][5] + xor_out[63][2][5] + xor_out[64][2][5];
assign sum_out[13][2][5] = xor_out[65][2][5] + xor_out[66][2][5] + xor_out[67][2][5] + xor_out[68][2][5] + xor_out[69][2][5];
assign sum_out[14][2][5] = xor_out[70][2][5] + xor_out[71][2][5] + xor_out[72][2][5] + xor_out[73][2][5] + xor_out[74][2][5];
assign sum_out[15][2][5] = xor_out[75][2][5] + xor_out[76][2][5] + xor_out[77][2][5] + xor_out[78][2][5] + xor_out[79][2][5];
assign sum_out[16][2][5] = xor_out[80][2][5] + xor_out[81][2][5] + xor_out[82][2][5] + xor_out[83][2][5] + xor_out[84][2][5];
assign sum_out[17][2][5] = xor_out[85][2][5] + xor_out[86][2][5] + xor_out[87][2][5] + xor_out[88][2][5] + xor_out[89][2][5];
assign sum_out[18][2][5] = xor_out[90][2][5] + xor_out[91][2][5] + xor_out[92][2][5] + xor_out[93][2][5] + xor_out[94][2][5];
assign sum_out[19][2][5] = xor_out[95][2][5] + xor_out[96][2][5] + xor_out[97][2][5] + xor_out[98][2][5] + xor_out[99][2][5];

assign sum_out[0][2][6] = xor_out[0][2][6] + xor_out[1][2][6] + xor_out[2][2][6] + xor_out[3][2][6] + xor_out[4][2][6];
assign sum_out[1][2][6] = xor_out[5][2][6] + xor_out[6][2][6] + xor_out[7][2][6] + xor_out[8][2][6] + xor_out[9][2][6];
assign sum_out[2][2][6] = xor_out[10][2][6] + xor_out[11][2][6] + xor_out[12][2][6] + xor_out[13][2][6] + xor_out[14][2][6];
assign sum_out[3][2][6] = xor_out[15][2][6] + xor_out[16][2][6] + xor_out[17][2][6] + xor_out[18][2][6] + xor_out[19][2][6];
assign sum_out[4][2][6] = xor_out[20][2][6] + xor_out[21][2][6] + xor_out[22][2][6] + xor_out[23][2][6] + xor_out[24][2][6];
assign sum_out[5][2][6] = xor_out[25][2][6] + xor_out[26][2][6] + xor_out[27][2][6] + xor_out[28][2][6] + xor_out[29][2][6];
assign sum_out[6][2][6] = xor_out[30][2][6] + xor_out[31][2][6] + xor_out[32][2][6] + xor_out[33][2][6] + xor_out[34][2][6];
assign sum_out[7][2][6] = xor_out[35][2][6] + xor_out[36][2][6] + xor_out[37][2][6] + xor_out[38][2][6] + xor_out[39][2][6];
assign sum_out[8][2][6] = xor_out[40][2][6] + xor_out[41][2][6] + xor_out[42][2][6] + xor_out[43][2][6] + xor_out[44][2][6];
assign sum_out[9][2][6] = xor_out[45][2][6] + xor_out[46][2][6] + xor_out[47][2][6] + xor_out[48][2][6] + xor_out[49][2][6];
assign sum_out[10][2][6] = xor_out[50][2][6] + xor_out[51][2][6] + xor_out[52][2][6] + xor_out[53][2][6] + xor_out[54][2][6];
assign sum_out[11][2][6] = xor_out[55][2][6] + xor_out[56][2][6] + xor_out[57][2][6] + xor_out[58][2][6] + xor_out[59][2][6];
assign sum_out[12][2][6] = xor_out[60][2][6] + xor_out[61][2][6] + xor_out[62][2][6] + xor_out[63][2][6] + xor_out[64][2][6];
assign sum_out[13][2][6] = xor_out[65][2][6] + xor_out[66][2][6] + xor_out[67][2][6] + xor_out[68][2][6] + xor_out[69][2][6];
assign sum_out[14][2][6] = xor_out[70][2][6] + xor_out[71][2][6] + xor_out[72][2][6] + xor_out[73][2][6] + xor_out[74][2][6];
assign sum_out[15][2][6] = xor_out[75][2][6] + xor_out[76][2][6] + xor_out[77][2][6] + xor_out[78][2][6] + xor_out[79][2][6];
assign sum_out[16][2][6] = xor_out[80][2][6] + xor_out[81][2][6] + xor_out[82][2][6] + xor_out[83][2][6] + xor_out[84][2][6];
assign sum_out[17][2][6] = xor_out[85][2][6] + xor_out[86][2][6] + xor_out[87][2][6] + xor_out[88][2][6] + xor_out[89][2][6];
assign sum_out[18][2][6] = xor_out[90][2][6] + xor_out[91][2][6] + xor_out[92][2][6] + xor_out[93][2][6] + xor_out[94][2][6];
assign sum_out[19][2][6] = xor_out[95][2][6] + xor_out[96][2][6] + xor_out[97][2][6] + xor_out[98][2][6] + xor_out[99][2][6];

assign sum_out[0][2][7] = xor_out[0][2][7] + xor_out[1][2][7] + xor_out[2][2][7] + xor_out[3][2][7] + xor_out[4][2][7];
assign sum_out[1][2][7] = xor_out[5][2][7] + xor_out[6][2][7] + xor_out[7][2][7] + xor_out[8][2][7] + xor_out[9][2][7];
assign sum_out[2][2][7] = xor_out[10][2][7] + xor_out[11][2][7] + xor_out[12][2][7] + xor_out[13][2][7] + xor_out[14][2][7];
assign sum_out[3][2][7] = xor_out[15][2][7] + xor_out[16][2][7] + xor_out[17][2][7] + xor_out[18][2][7] + xor_out[19][2][7];
assign sum_out[4][2][7] = xor_out[20][2][7] + xor_out[21][2][7] + xor_out[22][2][7] + xor_out[23][2][7] + xor_out[24][2][7];
assign sum_out[5][2][7] = xor_out[25][2][7] + xor_out[26][2][7] + xor_out[27][2][7] + xor_out[28][2][7] + xor_out[29][2][7];
assign sum_out[6][2][7] = xor_out[30][2][7] + xor_out[31][2][7] + xor_out[32][2][7] + xor_out[33][2][7] + xor_out[34][2][7];
assign sum_out[7][2][7] = xor_out[35][2][7] + xor_out[36][2][7] + xor_out[37][2][7] + xor_out[38][2][7] + xor_out[39][2][7];
assign sum_out[8][2][7] = xor_out[40][2][7] + xor_out[41][2][7] + xor_out[42][2][7] + xor_out[43][2][7] + xor_out[44][2][7];
assign sum_out[9][2][7] = xor_out[45][2][7] + xor_out[46][2][7] + xor_out[47][2][7] + xor_out[48][2][7] + xor_out[49][2][7];
assign sum_out[10][2][7] = xor_out[50][2][7] + xor_out[51][2][7] + xor_out[52][2][7] + xor_out[53][2][7] + xor_out[54][2][7];
assign sum_out[11][2][7] = xor_out[55][2][7] + xor_out[56][2][7] + xor_out[57][2][7] + xor_out[58][2][7] + xor_out[59][2][7];
assign sum_out[12][2][7] = xor_out[60][2][7] + xor_out[61][2][7] + xor_out[62][2][7] + xor_out[63][2][7] + xor_out[64][2][7];
assign sum_out[13][2][7] = xor_out[65][2][7] + xor_out[66][2][7] + xor_out[67][2][7] + xor_out[68][2][7] + xor_out[69][2][7];
assign sum_out[14][2][7] = xor_out[70][2][7] + xor_out[71][2][7] + xor_out[72][2][7] + xor_out[73][2][7] + xor_out[74][2][7];
assign sum_out[15][2][7] = xor_out[75][2][7] + xor_out[76][2][7] + xor_out[77][2][7] + xor_out[78][2][7] + xor_out[79][2][7];
assign sum_out[16][2][7] = xor_out[80][2][7] + xor_out[81][2][7] + xor_out[82][2][7] + xor_out[83][2][7] + xor_out[84][2][7];
assign sum_out[17][2][7] = xor_out[85][2][7] + xor_out[86][2][7] + xor_out[87][2][7] + xor_out[88][2][7] + xor_out[89][2][7];
assign sum_out[18][2][7] = xor_out[90][2][7] + xor_out[91][2][7] + xor_out[92][2][7] + xor_out[93][2][7] + xor_out[94][2][7];
assign sum_out[19][2][7] = xor_out[95][2][7] + xor_out[96][2][7] + xor_out[97][2][7] + xor_out[98][2][7] + xor_out[99][2][7];

assign sum_out[0][2][8] = xor_out[0][2][8] + xor_out[1][2][8] + xor_out[2][2][8] + xor_out[3][2][8] + xor_out[4][2][8];
assign sum_out[1][2][8] = xor_out[5][2][8] + xor_out[6][2][8] + xor_out[7][2][8] + xor_out[8][2][8] + xor_out[9][2][8];
assign sum_out[2][2][8] = xor_out[10][2][8] + xor_out[11][2][8] + xor_out[12][2][8] + xor_out[13][2][8] + xor_out[14][2][8];
assign sum_out[3][2][8] = xor_out[15][2][8] + xor_out[16][2][8] + xor_out[17][2][8] + xor_out[18][2][8] + xor_out[19][2][8];
assign sum_out[4][2][8] = xor_out[20][2][8] + xor_out[21][2][8] + xor_out[22][2][8] + xor_out[23][2][8] + xor_out[24][2][8];
assign sum_out[5][2][8] = xor_out[25][2][8] + xor_out[26][2][8] + xor_out[27][2][8] + xor_out[28][2][8] + xor_out[29][2][8];
assign sum_out[6][2][8] = xor_out[30][2][8] + xor_out[31][2][8] + xor_out[32][2][8] + xor_out[33][2][8] + xor_out[34][2][8];
assign sum_out[7][2][8] = xor_out[35][2][8] + xor_out[36][2][8] + xor_out[37][2][8] + xor_out[38][2][8] + xor_out[39][2][8];
assign sum_out[8][2][8] = xor_out[40][2][8] + xor_out[41][2][8] + xor_out[42][2][8] + xor_out[43][2][8] + xor_out[44][2][8];
assign sum_out[9][2][8] = xor_out[45][2][8] + xor_out[46][2][8] + xor_out[47][2][8] + xor_out[48][2][8] + xor_out[49][2][8];
assign sum_out[10][2][8] = xor_out[50][2][8] + xor_out[51][2][8] + xor_out[52][2][8] + xor_out[53][2][8] + xor_out[54][2][8];
assign sum_out[11][2][8] = xor_out[55][2][8] + xor_out[56][2][8] + xor_out[57][2][8] + xor_out[58][2][8] + xor_out[59][2][8];
assign sum_out[12][2][8] = xor_out[60][2][8] + xor_out[61][2][8] + xor_out[62][2][8] + xor_out[63][2][8] + xor_out[64][2][8];
assign sum_out[13][2][8] = xor_out[65][2][8] + xor_out[66][2][8] + xor_out[67][2][8] + xor_out[68][2][8] + xor_out[69][2][8];
assign sum_out[14][2][8] = xor_out[70][2][8] + xor_out[71][2][8] + xor_out[72][2][8] + xor_out[73][2][8] + xor_out[74][2][8];
assign sum_out[15][2][8] = xor_out[75][2][8] + xor_out[76][2][8] + xor_out[77][2][8] + xor_out[78][2][8] + xor_out[79][2][8];
assign sum_out[16][2][8] = xor_out[80][2][8] + xor_out[81][2][8] + xor_out[82][2][8] + xor_out[83][2][8] + xor_out[84][2][8];
assign sum_out[17][2][8] = xor_out[85][2][8] + xor_out[86][2][8] + xor_out[87][2][8] + xor_out[88][2][8] + xor_out[89][2][8];
assign sum_out[18][2][8] = xor_out[90][2][8] + xor_out[91][2][8] + xor_out[92][2][8] + xor_out[93][2][8] + xor_out[94][2][8];
assign sum_out[19][2][8] = xor_out[95][2][8] + xor_out[96][2][8] + xor_out[97][2][8] + xor_out[98][2][8] + xor_out[99][2][8];

assign sum_out[0][2][9] = xor_out[0][2][9] + xor_out[1][2][9] + xor_out[2][2][9] + xor_out[3][2][9] + xor_out[4][2][9];
assign sum_out[1][2][9] = xor_out[5][2][9] + xor_out[6][2][9] + xor_out[7][2][9] + xor_out[8][2][9] + xor_out[9][2][9];
assign sum_out[2][2][9] = xor_out[10][2][9] + xor_out[11][2][9] + xor_out[12][2][9] + xor_out[13][2][9] + xor_out[14][2][9];
assign sum_out[3][2][9] = xor_out[15][2][9] + xor_out[16][2][9] + xor_out[17][2][9] + xor_out[18][2][9] + xor_out[19][2][9];
assign sum_out[4][2][9] = xor_out[20][2][9] + xor_out[21][2][9] + xor_out[22][2][9] + xor_out[23][2][9] + xor_out[24][2][9];
assign sum_out[5][2][9] = xor_out[25][2][9] + xor_out[26][2][9] + xor_out[27][2][9] + xor_out[28][2][9] + xor_out[29][2][9];
assign sum_out[6][2][9] = xor_out[30][2][9] + xor_out[31][2][9] + xor_out[32][2][9] + xor_out[33][2][9] + xor_out[34][2][9];
assign sum_out[7][2][9] = xor_out[35][2][9] + xor_out[36][2][9] + xor_out[37][2][9] + xor_out[38][2][9] + xor_out[39][2][9];
assign sum_out[8][2][9] = xor_out[40][2][9] + xor_out[41][2][9] + xor_out[42][2][9] + xor_out[43][2][9] + xor_out[44][2][9];
assign sum_out[9][2][9] = xor_out[45][2][9] + xor_out[46][2][9] + xor_out[47][2][9] + xor_out[48][2][9] + xor_out[49][2][9];
assign sum_out[10][2][9] = xor_out[50][2][9] + xor_out[51][2][9] + xor_out[52][2][9] + xor_out[53][2][9] + xor_out[54][2][9];
assign sum_out[11][2][9] = xor_out[55][2][9] + xor_out[56][2][9] + xor_out[57][2][9] + xor_out[58][2][9] + xor_out[59][2][9];
assign sum_out[12][2][9] = xor_out[60][2][9] + xor_out[61][2][9] + xor_out[62][2][9] + xor_out[63][2][9] + xor_out[64][2][9];
assign sum_out[13][2][9] = xor_out[65][2][9] + xor_out[66][2][9] + xor_out[67][2][9] + xor_out[68][2][9] + xor_out[69][2][9];
assign sum_out[14][2][9] = xor_out[70][2][9] + xor_out[71][2][9] + xor_out[72][2][9] + xor_out[73][2][9] + xor_out[74][2][9];
assign sum_out[15][2][9] = xor_out[75][2][9] + xor_out[76][2][9] + xor_out[77][2][9] + xor_out[78][2][9] + xor_out[79][2][9];
assign sum_out[16][2][9] = xor_out[80][2][9] + xor_out[81][2][9] + xor_out[82][2][9] + xor_out[83][2][9] + xor_out[84][2][9];
assign sum_out[17][2][9] = xor_out[85][2][9] + xor_out[86][2][9] + xor_out[87][2][9] + xor_out[88][2][9] + xor_out[89][2][9];
assign sum_out[18][2][9] = xor_out[90][2][9] + xor_out[91][2][9] + xor_out[92][2][9] + xor_out[93][2][9] + xor_out[94][2][9];
assign sum_out[19][2][9] = xor_out[95][2][9] + xor_out[96][2][9] + xor_out[97][2][9] + xor_out[98][2][9] + xor_out[99][2][9];

assign sum_out[0][2][10] = xor_out[0][2][10] + xor_out[1][2][10] + xor_out[2][2][10] + xor_out[3][2][10] + xor_out[4][2][10];
assign sum_out[1][2][10] = xor_out[5][2][10] + xor_out[6][2][10] + xor_out[7][2][10] + xor_out[8][2][10] + xor_out[9][2][10];
assign sum_out[2][2][10] = xor_out[10][2][10] + xor_out[11][2][10] + xor_out[12][2][10] + xor_out[13][2][10] + xor_out[14][2][10];
assign sum_out[3][2][10] = xor_out[15][2][10] + xor_out[16][2][10] + xor_out[17][2][10] + xor_out[18][2][10] + xor_out[19][2][10];
assign sum_out[4][2][10] = xor_out[20][2][10] + xor_out[21][2][10] + xor_out[22][2][10] + xor_out[23][2][10] + xor_out[24][2][10];
assign sum_out[5][2][10] = xor_out[25][2][10] + xor_out[26][2][10] + xor_out[27][2][10] + xor_out[28][2][10] + xor_out[29][2][10];
assign sum_out[6][2][10] = xor_out[30][2][10] + xor_out[31][2][10] + xor_out[32][2][10] + xor_out[33][2][10] + xor_out[34][2][10];
assign sum_out[7][2][10] = xor_out[35][2][10] + xor_out[36][2][10] + xor_out[37][2][10] + xor_out[38][2][10] + xor_out[39][2][10];
assign sum_out[8][2][10] = xor_out[40][2][10] + xor_out[41][2][10] + xor_out[42][2][10] + xor_out[43][2][10] + xor_out[44][2][10];
assign sum_out[9][2][10] = xor_out[45][2][10] + xor_out[46][2][10] + xor_out[47][2][10] + xor_out[48][2][10] + xor_out[49][2][10];
assign sum_out[10][2][10] = xor_out[50][2][10] + xor_out[51][2][10] + xor_out[52][2][10] + xor_out[53][2][10] + xor_out[54][2][10];
assign sum_out[11][2][10] = xor_out[55][2][10] + xor_out[56][2][10] + xor_out[57][2][10] + xor_out[58][2][10] + xor_out[59][2][10];
assign sum_out[12][2][10] = xor_out[60][2][10] + xor_out[61][2][10] + xor_out[62][2][10] + xor_out[63][2][10] + xor_out[64][2][10];
assign sum_out[13][2][10] = xor_out[65][2][10] + xor_out[66][2][10] + xor_out[67][2][10] + xor_out[68][2][10] + xor_out[69][2][10];
assign sum_out[14][2][10] = xor_out[70][2][10] + xor_out[71][2][10] + xor_out[72][2][10] + xor_out[73][2][10] + xor_out[74][2][10];
assign sum_out[15][2][10] = xor_out[75][2][10] + xor_out[76][2][10] + xor_out[77][2][10] + xor_out[78][2][10] + xor_out[79][2][10];
assign sum_out[16][2][10] = xor_out[80][2][10] + xor_out[81][2][10] + xor_out[82][2][10] + xor_out[83][2][10] + xor_out[84][2][10];
assign sum_out[17][2][10] = xor_out[85][2][10] + xor_out[86][2][10] + xor_out[87][2][10] + xor_out[88][2][10] + xor_out[89][2][10];
assign sum_out[18][2][10] = xor_out[90][2][10] + xor_out[91][2][10] + xor_out[92][2][10] + xor_out[93][2][10] + xor_out[94][2][10];
assign sum_out[19][2][10] = xor_out[95][2][10] + xor_out[96][2][10] + xor_out[97][2][10] + xor_out[98][2][10] + xor_out[99][2][10];

assign sum_out[0][2][11] = xor_out[0][2][11] + xor_out[1][2][11] + xor_out[2][2][11] + xor_out[3][2][11] + xor_out[4][2][11];
assign sum_out[1][2][11] = xor_out[5][2][11] + xor_out[6][2][11] + xor_out[7][2][11] + xor_out[8][2][11] + xor_out[9][2][11];
assign sum_out[2][2][11] = xor_out[10][2][11] + xor_out[11][2][11] + xor_out[12][2][11] + xor_out[13][2][11] + xor_out[14][2][11];
assign sum_out[3][2][11] = xor_out[15][2][11] + xor_out[16][2][11] + xor_out[17][2][11] + xor_out[18][2][11] + xor_out[19][2][11];
assign sum_out[4][2][11] = xor_out[20][2][11] + xor_out[21][2][11] + xor_out[22][2][11] + xor_out[23][2][11] + xor_out[24][2][11];
assign sum_out[5][2][11] = xor_out[25][2][11] + xor_out[26][2][11] + xor_out[27][2][11] + xor_out[28][2][11] + xor_out[29][2][11];
assign sum_out[6][2][11] = xor_out[30][2][11] + xor_out[31][2][11] + xor_out[32][2][11] + xor_out[33][2][11] + xor_out[34][2][11];
assign sum_out[7][2][11] = xor_out[35][2][11] + xor_out[36][2][11] + xor_out[37][2][11] + xor_out[38][2][11] + xor_out[39][2][11];
assign sum_out[8][2][11] = xor_out[40][2][11] + xor_out[41][2][11] + xor_out[42][2][11] + xor_out[43][2][11] + xor_out[44][2][11];
assign sum_out[9][2][11] = xor_out[45][2][11] + xor_out[46][2][11] + xor_out[47][2][11] + xor_out[48][2][11] + xor_out[49][2][11];
assign sum_out[10][2][11] = xor_out[50][2][11] + xor_out[51][2][11] + xor_out[52][2][11] + xor_out[53][2][11] + xor_out[54][2][11];
assign sum_out[11][2][11] = xor_out[55][2][11] + xor_out[56][2][11] + xor_out[57][2][11] + xor_out[58][2][11] + xor_out[59][2][11];
assign sum_out[12][2][11] = xor_out[60][2][11] + xor_out[61][2][11] + xor_out[62][2][11] + xor_out[63][2][11] + xor_out[64][2][11];
assign sum_out[13][2][11] = xor_out[65][2][11] + xor_out[66][2][11] + xor_out[67][2][11] + xor_out[68][2][11] + xor_out[69][2][11];
assign sum_out[14][2][11] = xor_out[70][2][11] + xor_out[71][2][11] + xor_out[72][2][11] + xor_out[73][2][11] + xor_out[74][2][11];
assign sum_out[15][2][11] = xor_out[75][2][11] + xor_out[76][2][11] + xor_out[77][2][11] + xor_out[78][2][11] + xor_out[79][2][11];
assign sum_out[16][2][11] = xor_out[80][2][11] + xor_out[81][2][11] + xor_out[82][2][11] + xor_out[83][2][11] + xor_out[84][2][11];
assign sum_out[17][2][11] = xor_out[85][2][11] + xor_out[86][2][11] + xor_out[87][2][11] + xor_out[88][2][11] + xor_out[89][2][11];
assign sum_out[18][2][11] = xor_out[90][2][11] + xor_out[91][2][11] + xor_out[92][2][11] + xor_out[93][2][11] + xor_out[94][2][11];
assign sum_out[19][2][11] = xor_out[95][2][11] + xor_out[96][2][11] + xor_out[97][2][11] + xor_out[98][2][11] + xor_out[99][2][11];

assign sum_out[0][2][12] = xor_out[0][2][12] + xor_out[1][2][12] + xor_out[2][2][12] + xor_out[3][2][12] + xor_out[4][2][12];
assign sum_out[1][2][12] = xor_out[5][2][12] + xor_out[6][2][12] + xor_out[7][2][12] + xor_out[8][2][12] + xor_out[9][2][12];
assign sum_out[2][2][12] = xor_out[10][2][12] + xor_out[11][2][12] + xor_out[12][2][12] + xor_out[13][2][12] + xor_out[14][2][12];
assign sum_out[3][2][12] = xor_out[15][2][12] + xor_out[16][2][12] + xor_out[17][2][12] + xor_out[18][2][12] + xor_out[19][2][12];
assign sum_out[4][2][12] = xor_out[20][2][12] + xor_out[21][2][12] + xor_out[22][2][12] + xor_out[23][2][12] + xor_out[24][2][12];
assign sum_out[5][2][12] = xor_out[25][2][12] + xor_out[26][2][12] + xor_out[27][2][12] + xor_out[28][2][12] + xor_out[29][2][12];
assign sum_out[6][2][12] = xor_out[30][2][12] + xor_out[31][2][12] + xor_out[32][2][12] + xor_out[33][2][12] + xor_out[34][2][12];
assign sum_out[7][2][12] = xor_out[35][2][12] + xor_out[36][2][12] + xor_out[37][2][12] + xor_out[38][2][12] + xor_out[39][2][12];
assign sum_out[8][2][12] = xor_out[40][2][12] + xor_out[41][2][12] + xor_out[42][2][12] + xor_out[43][2][12] + xor_out[44][2][12];
assign sum_out[9][2][12] = xor_out[45][2][12] + xor_out[46][2][12] + xor_out[47][2][12] + xor_out[48][2][12] + xor_out[49][2][12];
assign sum_out[10][2][12] = xor_out[50][2][12] + xor_out[51][2][12] + xor_out[52][2][12] + xor_out[53][2][12] + xor_out[54][2][12];
assign sum_out[11][2][12] = xor_out[55][2][12] + xor_out[56][2][12] + xor_out[57][2][12] + xor_out[58][2][12] + xor_out[59][2][12];
assign sum_out[12][2][12] = xor_out[60][2][12] + xor_out[61][2][12] + xor_out[62][2][12] + xor_out[63][2][12] + xor_out[64][2][12];
assign sum_out[13][2][12] = xor_out[65][2][12] + xor_out[66][2][12] + xor_out[67][2][12] + xor_out[68][2][12] + xor_out[69][2][12];
assign sum_out[14][2][12] = xor_out[70][2][12] + xor_out[71][2][12] + xor_out[72][2][12] + xor_out[73][2][12] + xor_out[74][2][12];
assign sum_out[15][2][12] = xor_out[75][2][12] + xor_out[76][2][12] + xor_out[77][2][12] + xor_out[78][2][12] + xor_out[79][2][12];
assign sum_out[16][2][12] = xor_out[80][2][12] + xor_out[81][2][12] + xor_out[82][2][12] + xor_out[83][2][12] + xor_out[84][2][12];
assign sum_out[17][2][12] = xor_out[85][2][12] + xor_out[86][2][12] + xor_out[87][2][12] + xor_out[88][2][12] + xor_out[89][2][12];
assign sum_out[18][2][12] = xor_out[90][2][12] + xor_out[91][2][12] + xor_out[92][2][12] + xor_out[93][2][12] + xor_out[94][2][12];
assign sum_out[19][2][12] = xor_out[95][2][12] + xor_out[96][2][12] + xor_out[97][2][12] + xor_out[98][2][12] + xor_out[99][2][12];

assign sum_out[0][2][13] = xor_out[0][2][13] + xor_out[1][2][13] + xor_out[2][2][13] + xor_out[3][2][13] + xor_out[4][2][13];
assign sum_out[1][2][13] = xor_out[5][2][13] + xor_out[6][2][13] + xor_out[7][2][13] + xor_out[8][2][13] + xor_out[9][2][13];
assign sum_out[2][2][13] = xor_out[10][2][13] + xor_out[11][2][13] + xor_out[12][2][13] + xor_out[13][2][13] + xor_out[14][2][13];
assign sum_out[3][2][13] = xor_out[15][2][13] + xor_out[16][2][13] + xor_out[17][2][13] + xor_out[18][2][13] + xor_out[19][2][13];
assign sum_out[4][2][13] = xor_out[20][2][13] + xor_out[21][2][13] + xor_out[22][2][13] + xor_out[23][2][13] + xor_out[24][2][13];
assign sum_out[5][2][13] = xor_out[25][2][13] + xor_out[26][2][13] + xor_out[27][2][13] + xor_out[28][2][13] + xor_out[29][2][13];
assign sum_out[6][2][13] = xor_out[30][2][13] + xor_out[31][2][13] + xor_out[32][2][13] + xor_out[33][2][13] + xor_out[34][2][13];
assign sum_out[7][2][13] = xor_out[35][2][13] + xor_out[36][2][13] + xor_out[37][2][13] + xor_out[38][2][13] + xor_out[39][2][13];
assign sum_out[8][2][13] = xor_out[40][2][13] + xor_out[41][2][13] + xor_out[42][2][13] + xor_out[43][2][13] + xor_out[44][2][13];
assign sum_out[9][2][13] = xor_out[45][2][13] + xor_out[46][2][13] + xor_out[47][2][13] + xor_out[48][2][13] + xor_out[49][2][13];
assign sum_out[10][2][13] = xor_out[50][2][13] + xor_out[51][2][13] + xor_out[52][2][13] + xor_out[53][2][13] + xor_out[54][2][13];
assign sum_out[11][2][13] = xor_out[55][2][13] + xor_out[56][2][13] + xor_out[57][2][13] + xor_out[58][2][13] + xor_out[59][2][13];
assign sum_out[12][2][13] = xor_out[60][2][13] + xor_out[61][2][13] + xor_out[62][2][13] + xor_out[63][2][13] + xor_out[64][2][13];
assign sum_out[13][2][13] = xor_out[65][2][13] + xor_out[66][2][13] + xor_out[67][2][13] + xor_out[68][2][13] + xor_out[69][2][13];
assign sum_out[14][2][13] = xor_out[70][2][13] + xor_out[71][2][13] + xor_out[72][2][13] + xor_out[73][2][13] + xor_out[74][2][13];
assign sum_out[15][2][13] = xor_out[75][2][13] + xor_out[76][2][13] + xor_out[77][2][13] + xor_out[78][2][13] + xor_out[79][2][13];
assign sum_out[16][2][13] = xor_out[80][2][13] + xor_out[81][2][13] + xor_out[82][2][13] + xor_out[83][2][13] + xor_out[84][2][13];
assign sum_out[17][2][13] = xor_out[85][2][13] + xor_out[86][2][13] + xor_out[87][2][13] + xor_out[88][2][13] + xor_out[89][2][13];
assign sum_out[18][2][13] = xor_out[90][2][13] + xor_out[91][2][13] + xor_out[92][2][13] + xor_out[93][2][13] + xor_out[94][2][13];
assign sum_out[19][2][13] = xor_out[95][2][13] + xor_out[96][2][13] + xor_out[97][2][13] + xor_out[98][2][13] + xor_out[99][2][13];

assign sum_out[0][2][14] = xor_out[0][2][14] + xor_out[1][2][14] + xor_out[2][2][14] + xor_out[3][2][14] + xor_out[4][2][14];
assign sum_out[1][2][14] = xor_out[5][2][14] + xor_out[6][2][14] + xor_out[7][2][14] + xor_out[8][2][14] + xor_out[9][2][14];
assign sum_out[2][2][14] = xor_out[10][2][14] + xor_out[11][2][14] + xor_out[12][2][14] + xor_out[13][2][14] + xor_out[14][2][14];
assign sum_out[3][2][14] = xor_out[15][2][14] + xor_out[16][2][14] + xor_out[17][2][14] + xor_out[18][2][14] + xor_out[19][2][14];
assign sum_out[4][2][14] = xor_out[20][2][14] + xor_out[21][2][14] + xor_out[22][2][14] + xor_out[23][2][14] + xor_out[24][2][14];
assign sum_out[5][2][14] = xor_out[25][2][14] + xor_out[26][2][14] + xor_out[27][2][14] + xor_out[28][2][14] + xor_out[29][2][14];
assign sum_out[6][2][14] = xor_out[30][2][14] + xor_out[31][2][14] + xor_out[32][2][14] + xor_out[33][2][14] + xor_out[34][2][14];
assign sum_out[7][2][14] = xor_out[35][2][14] + xor_out[36][2][14] + xor_out[37][2][14] + xor_out[38][2][14] + xor_out[39][2][14];
assign sum_out[8][2][14] = xor_out[40][2][14] + xor_out[41][2][14] + xor_out[42][2][14] + xor_out[43][2][14] + xor_out[44][2][14];
assign sum_out[9][2][14] = xor_out[45][2][14] + xor_out[46][2][14] + xor_out[47][2][14] + xor_out[48][2][14] + xor_out[49][2][14];
assign sum_out[10][2][14] = xor_out[50][2][14] + xor_out[51][2][14] + xor_out[52][2][14] + xor_out[53][2][14] + xor_out[54][2][14];
assign sum_out[11][2][14] = xor_out[55][2][14] + xor_out[56][2][14] + xor_out[57][2][14] + xor_out[58][2][14] + xor_out[59][2][14];
assign sum_out[12][2][14] = xor_out[60][2][14] + xor_out[61][2][14] + xor_out[62][2][14] + xor_out[63][2][14] + xor_out[64][2][14];
assign sum_out[13][2][14] = xor_out[65][2][14] + xor_out[66][2][14] + xor_out[67][2][14] + xor_out[68][2][14] + xor_out[69][2][14];
assign sum_out[14][2][14] = xor_out[70][2][14] + xor_out[71][2][14] + xor_out[72][2][14] + xor_out[73][2][14] + xor_out[74][2][14];
assign sum_out[15][2][14] = xor_out[75][2][14] + xor_out[76][2][14] + xor_out[77][2][14] + xor_out[78][2][14] + xor_out[79][2][14];
assign sum_out[16][2][14] = xor_out[80][2][14] + xor_out[81][2][14] + xor_out[82][2][14] + xor_out[83][2][14] + xor_out[84][2][14];
assign sum_out[17][2][14] = xor_out[85][2][14] + xor_out[86][2][14] + xor_out[87][2][14] + xor_out[88][2][14] + xor_out[89][2][14];
assign sum_out[18][2][14] = xor_out[90][2][14] + xor_out[91][2][14] + xor_out[92][2][14] + xor_out[93][2][14] + xor_out[94][2][14];
assign sum_out[19][2][14] = xor_out[95][2][14] + xor_out[96][2][14] + xor_out[97][2][14] + xor_out[98][2][14] + xor_out[99][2][14];

assign sum_out[0][2][15] = xor_out[0][2][15] + xor_out[1][2][15] + xor_out[2][2][15] + xor_out[3][2][15] + xor_out[4][2][15];
assign sum_out[1][2][15] = xor_out[5][2][15] + xor_out[6][2][15] + xor_out[7][2][15] + xor_out[8][2][15] + xor_out[9][2][15];
assign sum_out[2][2][15] = xor_out[10][2][15] + xor_out[11][2][15] + xor_out[12][2][15] + xor_out[13][2][15] + xor_out[14][2][15];
assign sum_out[3][2][15] = xor_out[15][2][15] + xor_out[16][2][15] + xor_out[17][2][15] + xor_out[18][2][15] + xor_out[19][2][15];
assign sum_out[4][2][15] = xor_out[20][2][15] + xor_out[21][2][15] + xor_out[22][2][15] + xor_out[23][2][15] + xor_out[24][2][15];
assign sum_out[5][2][15] = xor_out[25][2][15] + xor_out[26][2][15] + xor_out[27][2][15] + xor_out[28][2][15] + xor_out[29][2][15];
assign sum_out[6][2][15] = xor_out[30][2][15] + xor_out[31][2][15] + xor_out[32][2][15] + xor_out[33][2][15] + xor_out[34][2][15];
assign sum_out[7][2][15] = xor_out[35][2][15] + xor_out[36][2][15] + xor_out[37][2][15] + xor_out[38][2][15] + xor_out[39][2][15];
assign sum_out[8][2][15] = xor_out[40][2][15] + xor_out[41][2][15] + xor_out[42][2][15] + xor_out[43][2][15] + xor_out[44][2][15];
assign sum_out[9][2][15] = xor_out[45][2][15] + xor_out[46][2][15] + xor_out[47][2][15] + xor_out[48][2][15] + xor_out[49][2][15];
assign sum_out[10][2][15] = xor_out[50][2][15] + xor_out[51][2][15] + xor_out[52][2][15] + xor_out[53][2][15] + xor_out[54][2][15];
assign sum_out[11][2][15] = xor_out[55][2][15] + xor_out[56][2][15] + xor_out[57][2][15] + xor_out[58][2][15] + xor_out[59][2][15];
assign sum_out[12][2][15] = xor_out[60][2][15] + xor_out[61][2][15] + xor_out[62][2][15] + xor_out[63][2][15] + xor_out[64][2][15];
assign sum_out[13][2][15] = xor_out[65][2][15] + xor_out[66][2][15] + xor_out[67][2][15] + xor_out[68][2][15] + xor_out[69][2][15];
assign sum_out[14][2][15] = xor_out[70][2][15] + xor_out[71][2][15] + xor_out[72][2][15] + xor_out[73][2][15] + xor_out[74][2][15];
assign sum_out[15][2][15] = xor_out[75][2][15] + xor_out[76][2][15] + xor_out[77][2][15] + xor_out[78][2][15] + xor_out[79][2][15];
assign sum_out[16][2][15] = xor_out[80][2][15] + xor_out[81][2][15] + xor_out[82][2][15] + xor_out[83][2][15] + xor_out[84][2][15];
assign sum_out[17][2][15] = xor_out[85][2][15] + xor_out[86][2][15] + xor_out[87][2][15] + xor_out[88][2][15] + xor_out[89][2][15];
assign sum_out[18][2][15] = xor_out[90][2][15] + xor_out[91][2][15] + xor_out[92][2][15] + xor_out[93][2][15] + xor_out[94][2][15];
assign sum_out[19][2][15] = xor_out[95][2][15] + xor_out[96][2][15] + xor_out[97][2][15] + xor_out[98][2][15] + xor_out[99][2][15];

assign sum_out[0][2][16] = xor_out[0][2][16] + xor_out[1][2][16] + xor_out[2][2][16] + xor_out[3][2][16] + xor_out[4][2][16];
assign sum_out[1][2][16] = xor_out[5][2][16] + xor_out[6][2][16] + xor_out[7][2][16] + xor_out[8][2][16] + xor_out[9][2][16];
assign sum_out[2][2][16] = xor_out[10][2][16] + xor_out[11][2][16] + xor_out[12][2][16] + xor_out[13][2][16] + xor_out[14][2][16];
assign sum_out[3][2][16] = xor_out[15][2][16] + xor_out[16][2][16] + xor_out[17][2][16] + xor_out[18][2][16] + xor_out[19][2][16];
assign sum_out[4][2][16] = xor_out[20][2][16] + xor_out[21][2][16] + xor_out[22][2][16] + xor_out[23][2][16] + xor_out[24][2][16];
assign sum_out[5][2][16] = xor_out[25][2][16] + xor_out[26][2][16] + xor_out[27][2][16] + xor_out[28][2][16] + xor_out[29][2][16];
assign sum_out[6][2][16] = xor_out[30][2][16] + xor_out[31][2][16] + xor_out[32][2][16] + xor_out[33][2][16] + xor_out[34][2][16];
assign sum_out[7][2][16] = xor_out[35][2][16] + xor_out[36][2][16] + xor_out[37][2][16] + xor_out[38][2][16] + xor_out[39][2][16];
assign sum_out[8][2][16] = xor_out[40][2][16] + xor_out[41][2][16] + xor_out[42][2][16] + xor_out[43][2][16] + xor_out[44][2][16];
assign sum_out[9][2][16] = xor_out[45][2][16] + xor_out[46][2][16] + xor_out[47][2][16] + xor_out[48][2][16] + xor_out[49][2][16];
assign sum_out[10][2][16] = xor_out[50][2][16] + xor_out[51][2][16] + xor_out[52][2][16] + xor_out[53][2][16] + xor_out[54][2][16];
assign sum_out[11][2][16] = xor_out[55][2][16] + xor_out[56][2][16] + xor_out[57][2][16] + xor_out[58][2][16] + xor_out[59][2][16];
assign sum_out[12][2][16] = xor_out[60][2][16] + xor_out[61][2][16] + xor_out[62][2][16] + xor_out[63][2][16] + xor_out[64][2][16];
assign sum_out[13][2][16] = xor_out[65][2][16] + xor_out[66][2][16] + xor_out[67][2][16] + xor_out[68][2][16] + xor_out[69][2][16];
assign sum_out[14][2][16] = xor_out[70][2][16] + xor_out[71][2][16] + xor_out[72][2][16] + xor_out[73][2][16] + xor_out[74][2][16];
assign sum_out[15][2][16] = xor_out[75][2][16] + xor_out[76][2][16] + xor_out[77][2][16] + xor_out[78][2][16] + xor_out[79][2][16];
assign sum_out[16][2][16] = xor_out[80][2][16] + xor_out[81][2][16] + xor_out[82][2][16] + xor_out[83][2][16] + xor_out[84][2][16];
assign sum_out[17][2][16] = xor_out[85][2][16] + xor_out[86][2][16] + xor_out[87][2][16] + xor_out[88][2][16] + xor_out[89][2][16];
assign sum_out[18][2][16] = xor_out[90][2][16] + xor_out[91][2][16] + xor_out[92][2][16] + xor_out[93][2][16] + xor_out[94][2][16];
assign sum_out[19][2][16] = xor_out[95][2][16] + xor_out[96][2][16] + xor_out[97][2][16] + xor_out[98][2][16] + xor_out[99][2][16];

assign sum_out[0][2][17] = xor_out[0][2][17] + xor_out[1][2][17] + xor_out[2][2][17] + xor_out[3][2][17] + xor_out[4][2][17];
assign sum_out[1][2][17] = xor_out[5][2][17] + xor_out[6][2][17] + xor_out[7][2][17] + xor_out[8][2][17] + xor_out[9][2][17];
assign sum_out[2][2][17] = xor_out[10][2][17] + xor_out[11][2][17] + xor_out[12][2][17] + xor_out[13][2][17] + xor_out[14][2][17];
assign sum_out[3][2][17] = xor_out[15][2][17] + xor_out[16][2][17] + xor_out[17][2][17] + xor_out[18][2][17] + xor_out[19][2][17];
assign sum_out[4][2][17] = xor_out[20][2][17] + xor_out[21][2][17] + xor_out[22][2][17] + xor_out[23][2][17] + xor_out[24][2][17];
assign sum_out[5][2][17] = xor_out[25][2][17] + xor_out[26][2][17] + xor_out[27][2][17] + xor_out[28][2][17] + xor_out[29][2][17];
assign sum_out[6][2][17] = xor_out[30][2][17] + xor_out[31][2][17] + xor_out[32][2][17] + xor_out[33][2][17] + xor_out[34][2][17];
assign sum_out[7][2][17] = xor_out[35][2][17] + xor_out[36][2][17] + xor_out[37][2][17] + xor_out[38][2][17] + xor_out[39][2][17];
assign sum_out[8][2][17] = xor_out[40][2][17] + xor_out[41][2][17] + xor_out[42][2][17] + xor_out[43][2][17] + xor_out[44][2][17];
assign sum_out[9][2][17] = xor_out[45][2][17] + xor_out[46][2][17] + xor_out[47][2][17] + xor_out[48][2][17] + xor_out[49][2][17];
assign sum_out[10][2][17] = xor_out[50][2][17] + xor_out[51][2][17] + xor_out[52][2][17] + xor_out[53][2][17] + xor_out[54][2][17];
assign sum_out[11][2][17] = xor_out[55][2][17] + xor_out[56][2][17] + xor_out[57][2][17] + xor_out[58][2][17] + xor_out[59][2][17];
assign sum_out[12][2][17] = xor_out[60][2][17] + xor_out[61][2][17] + xor_out[62][2][17] + xor_out[63][2][17] + xor_out[64][2][17];
assign sum_out[13][2][17] = xor_out[65][2][17] + xor_out[66][2][17] + xor_out[67][2][17] + xor_out[68][2][17] + xor_out[69][2][17];
assign sum_out[14][2][17] = xor_out[70][2][17] + xor_out[71][2][17] + xor_out[72][2][17] + xor_out[73][2][17] + xor_out[74][2][17];
assign sum_out[15][2][17] = xor_out[75][2][17] + xor_out[76][2][17] + xor_out[77][2][17] + xor_out[78][2][17] + xor_out[79][2][17];
assign sum_out[16][2][17] = xor_out[80][2][17] + xor_out[81][2][17] + xor_out[82][2][17] + xor_out[83][2][17] + xor_out[84][2][17];
assign sum_out[17][2][17] = xor_out[85][2][17] + xor_out[86][2][17] + xor_out[87][2][17] + xor_out[88][2][17] + xor_out[89][2][17];
assign sum_out[18][2][17] = xor_out[90][2][17] + xor_out[91][2][17] + xor_out[92][2][17] + xor_out[93][2][17] + xor_out[94][2][17];
assign sum_out[19][2][17] = xor_out[95][2][17] + xor_out[96][2][17] + xor_out[97][2][17] + xor_out[98][2][17] + xor_out[99][2][17];

assign sum_out[0][2][18] = xor_out[0][2][18] + xor_out[1][2][18] + xor_out[2][2][18] + xor_out[3][2][18] + xor_out[4][2][18];
assign sum_out[1][2][18] = xor_out[5][2][18] + xor_out[6][2][18] + xor_out[7][2][18] + xor_out[8][2][18] + xor_out[9][2][18];
assign sum_out[2][2][18] = xor_out[10][2][18] + xor_out[11][2][18] + xor_out[12][2][18] + xor_out[13][2][18] + xor_out[14][2][18];
assign sum_out[3][2][18] = xor_out[15][2][18] + xor_out[16][2][18] + xor_out[17][2][18] + xor_out[18][2][18] + xor_out[19][2][18];
assign sum_out[4][2][18] = xor_out[20][2][18] + xor_out[21][2][18] + xor_out[22][2][18] + xor_out[23][2][18] + xor_out[24][2][18];
assign sum_out[5][2][18] = xor_out[25][2][18] + xor_out[26][2][18] + xor_out[27][2][18] + xor_out[28][2][18] + xor_out[29][2][18];
assign sum_out[6][2][18] = xor_out[30][2][18] + xor_out[31][2][18] + xor_out[32][2][18] + xor_out[33][2][18] + xor_out[34][2][18];
assign sum_out[7][2][18] = xor_out[35][2][18] + xor_out[36][2][18] + xor_out[37][2][18] + xor_out[38][2][18] + xor_out[39][2][18];
assign sum_out[8][2][18] = xor_out[40][2][18] + xor_out[41][2][18] + xor_out[42][2][18] + xor_out[43][2][18] + xor_out[44][2][18];
assign sum_out[9][2][18] = xor_out[45][2][18] + xor_out[46][2][18] + xor_out[47][2][18] + xor_out[48][2][18] + xor_out[49][2][18];
assign sum_out[10][2][18] = xor_out[50][2][18] + xor_out[51][2][18] + xor_out[52][2][18] + xor_out[53][2][18] + xor_out[54][2][18];
assign sum_out[11][2][18] = xor_out[55][2][18] + xor_out[56][2][18] + xor_out[57][2][18] + xor_out[58][2][18] + xor_out[59][2][18];
assign sum_out[12][2][18] = xor_out[60][2][18] + xor_out[61][2][18] + xor_out[62][2][18] + xor_out[63][2][18] + xor_out[64][2][18];
assign sum_out[13][2][18] = xor_out[65][2][18] + xor_out[66][2][18] + xor_out[67][2][18] + xor_out[68][2][18] + xor_out[69][2][18];
assign sum_out[14][2][18] = xor_out[70][2][18] + xor_out[71][2][18] + xor_out[72][2][18] + xor_out[73][2][18] + xor_out[74][2][18];
assign sum_out[15][2][18] = xor_out[75][2][18] + xor_out[76][2][18] + xor_out[77][2][18] + xor_out[78][2][18] + xor_out[79][2][18];
assign sum_out[16][2][18] = xor_out[80][2][18] + xor_out[81][2][18] + xor_out[82][2][18] + xor_out[83][2][18] + xor_out[84][2][18];
assign sum_out[17][2][18] = xor_out[85][2][18] + xor_out[86][2][18] + xor_out[87][2][18] + xor_out[88][2][18] + xor_out[89][2][18];
assign sum_out[18][2][18] = xor_out[90][2][18] + xor_out[91][2][18] + xor_out[92][2][18] + xor_out[93][2][18] + xor_out[94][2][18];
assign sum_out[19][2][18] = xor_out[95][2][18] + xor_out[96][2][18] + xor_out[97][2][18] + xor_out[98][2][18] + xor_out[99][2][18];

assign sum_out[0][2][19] = xor_out[0][2][19] + xor_out[1][2][19] + xor_out[2][2][19] + xor_out[3][2][19] + xor_out[4][2][19];
assign sum_out[1][2][19] = xor_out[5][2][19] + xor_out[6][2][19] + xor_out[7][2][19] + xor_out[8][2][19] + xor_out[9][2][19];
assign sum_out[2][2][19] = xor_out[10][2][19] + xor_out[11][2][19] + xor_out[12][2][19] + xor_out[13][2][19] + xor_out[14][2][19];
assign sum_out[3][2][19] = xor_out[15][2][19] + xor_out[16][2][19] + xor_out[17][2][19] + xor_out[18][2][19] + xor_out[19][2][19];
assign sum_out[4][2][19] = xor_out[20][2][19] + xor_out[21][2][19] + xor_out[22][2][19] + xor_out[23][2][19] + xor_out[24][2][19];
assign sum_out[5][2][19] = xor_out[25][2][19] + xor_out[26][2][19] + xor_out[27][2][19] + xor_out[28][2][19] + xor_out[29][2][19];
assign sum_out[6][2][19] = xor_out[30][2][19] + xor_out[31][2][19] + xor_out[32][2][19] + xor_out[33][2][19] + xor_out[34][2][19];
assign sum_out[7][2][19] = xor_out[35][2][19] + xor_out[36][2][19] + xor_out[37][2][19] + xor_out[38][2][19] + xor_out[39][2][19];
assign sum_out[8][2][19] = xor_out[40][2][19] + xor_out[41][2][19] + xor_out[42][2][19] + xor_out[43][2][19] + xor_out[44][2][19];
assign sum_out[9][2][19] = xor_out[45][2][19] + xor_out[46][2][19] + xor_out[47][2][19] + xor_out[48][2][19] + xor_out[49][2][19];
assign sum_out[10][2][19] = xor_out[50][2][19] + xor_out[51][2][19] + xor_out[52][2][19] + xor_out[53][2][19] + xor_out[54][2][19];
assign sum_out[11][2][19] = xor_out[55][2][19] + xor_out[56][2][19] + xor_out[57][2][19] + xor_out[58][2][19] + xor_out[59][2][19];
assign sum_out[12][2][19] = xor_out[60][2][19] + xor_out[61][2][19] + xor_out[62][2][19] + xor_out[63][2][19] + xor_out[64][2][19];
assign sum_out[13][2][19] = xor_out[65][2][19] + xor_out[66][2][19] + xor_out[67][2][19] + xor_out[68][2][19] + xor_out[69][2][19];
assign sum_out[14][2][19] = xor_out[70][2][19] + xor_out[71][2][19] + xor_out[72][2][19] + xor_out[73][2][19] + xor_out[74][2][19];
assign sum_out[15][2][19] = xor_out[75][2][19] + xor_out[76][2][19] + xor_out[77][2][19] + xor_out[78][2][19] + xor_out[79][2][19];
assign sum_out[16][2][19] = xor_out[80][2][19] + xor_out[81][2][19] + xor_out[82][2][19] + xor_out[83][2][19] + xor_out[84][2][19];
assign sum_out[17][2][19] = xor_out[85][2][19] + xor_out[86][2][19] + xor_out[87][2][19] + xor_out[88][2][19] + xor_out[89][2][19];
assign sum_out[18][2][19] = xor_out[90][2][19] + xor_out[91][2][19] + xor_out[92][2][19] + xor_out[93][2][19] + xor_out[94][2][19];
assign sum_out[19][2][19] = xor_out[95][2][19] + xor_out[96][2][19] + xor_out[97][2][19] + xor_out[98][2][19] + xor_out[99][2][19];

assign sum_out[0][2][20] = xor_out[0][2][20] + xor_out[1][2][20] + xor_out[2][2][20] + xor_out[3][2][20] + xor_out[4][2][20];
assign sum_out[1][2][20] = xor_out[5][2][20] + xor_out[6][2][20] + xor_out[7][2][20] + xor_out[8][2][20] + xor_out[9][2][20];
assign sum_out[2][2][20] = xor_out[10][2][20] + xor_out[11][2][20] + xor_out[12][2][20] + xor_out[13][2][20] + xor_out[14][2][20];
assign sum_out[3][2][20] = xor_out[15][2][20] + xor_out[16][2][20] + xor_out[17][2][20] + xor_out[18][2][20] + xor_out[19][2][20];
assign sum_out[4][2][20] = xor_out[20][2][20] + xor_out[21][2][20] + xor_out[22][2][20] + xor_out[23][2][20] + xor_out[24][2][20];
assign sum_out[5][2][20] = xor_out[25][2][20] + xor_out[26][2][20] + xor_out[27][2][20] + xor_out[28][2][20] + xor_out[29][2][20];
assign sum_out[6][2][20] = xor_out[30][2][20] + xor_out[31][2][20] + xor_out[32][2][20] + xor_out[33][2][20] + xor_out[34][2][20];
assign sum_out[7][2][20] = xor_out[35][2][20] + xor_out[36][2][20] + xor_out[37][2][20] + xor_out[38][2][20] + xor_out[39][2][20];
assign sum_out[8][2][20] = xor_out[40][2][20] + xor_out[41][2][20] + xor_out[42][2][20] + xor_out[43][2][20] + xor_out[44][2][20];
assign sum_out[9][2][20] = xor_out[45][2][20] + xor_out[46][2][20] + xor_out[47][2][20] + xor_out[48][2][20] + xor_out[49][2][20];
assign sum_out[10][2][20] = xor_out[50][2][20] + xor_out[51][2][20] + xor_out[52][2][20] + xor_out[53][2][20] + xor_out[54][2][20];
assign sum_out[11][2][20] = xor_out[55][2][20] + xor_out[56][2][20] + xor_out[57][2][20] + xor_out[58][2][20] + xor_out[59][2][20];
assign sum_out[12][2][20] = xor_out[60][2][20] + xor_out[61][2][20] + xor_out[62][2][20] + xor_out[63][2][20] + xor_out[64][2][20];
assign sum_out[13][2][20] = xor_out[65][2][20] + xor_out[66][2][20] + xor_out[67][2][20] + xor_out[68][2][20] + xor_out[69][2][20];
assign sum_out[14][2][20] = xor_out[70][2][20] + xor_out[71][2][20] + xor_out[72][2][20] + xor_out[73][2][20] + xor_out[74][2][20];
assign sum_out[15][2][20] = xor_out[75][2][20] + xor_out[76][2][20] + xor_out[77][2][20] + xor_out[78][2][20] + xor_out[79][2][20];
assign sum_out[16][2][20] = xor_out[80][2][20] + xor_out[81][2][20] + xor_out[82][2][20] + xor_out[83][2][20] + xor_out[84][2][20];
assign sum_out[17][2][20] = xor_out[85][2][20] + xor_out[86][2][20] + xor_out[87][2][20] + xor_out[88][2][20] + xor_out[89][2][20];
assign sum_out[18][2][20] = xor_out[90][2][20] + xor_out[91][2][20] + xor_out[92][2][20] + xor_out[93][2][20] + xor_out[94][2][20];
assign sum_out[19][2][20] = xor_out[95][2][20] + xor_out[96][2][20] + xor_out[97][2][20] + xor_out[98][2][20] + xor_out[99][2][20];

assign sum_out[0][2][21] = xor_out[0][2][21] + xor_out[1][2][21] + xor_out[2][2][21] + xor_out[3][2][21] + xor_out[4][2][21];
assign sum_out[1][2][21] = xor_out[5][2][21] + xor_out[6][2][21] + xor_out[7][2][21] + xor_out[8][2][21] + xor_out[9][2][21];
assign sum_out[2][2][21] = xor_out[10][2][21] + xor_out[11][2][21] + xor_out[12][2][21] + xor_out[13][2][21] + xor_out[14][2][21];
assign sum_out[3][2][21] = xor_out[15][2][21] + xor_out[16][2][21] + xor_out[17][2][21] + xor_out[18][2][21] + xor_out[19][2][21];
assign sum_out[4][2][21] = xor_out[20][2][21] + xor_out[21][2][21] + xor_out[22][2][21] + xor_out[23][2][21] + xor_out[24][2][21];
assign sum_out[5][2][21] = xor_out[25][2][21] + xor_out[26][2][21] + xor_out[27][2][21] + xor_out[28][2][21] + xor_out[29][2][21];
assign sum_out[6][2][21] = xor_out[30][2][21] + xor_out[31][2][21] + xor_out[32][2][21] + xor_out[33][2][21] + xor_out[34][2][21];
assign sum_out[7][2][21] = xor_out[35][2][21] + xor_out[36][2][21] + xor_out[37][2][21] + xor_out[38][2][21] + xor_out[39][2][21];
assign sum_out[8][2][21] = xor_out[40][2][21] + xor_out[41][2][21] + xor_out[42][2][21] + xor_out[43][2][21] + xor_out[44][2][21];
assign sum_out[9][2][21] = xor_out[45][2][21] + xor_out[46][2][21] + xor_out[47][2][21] + xor_out[48][2][21] + xor_out[49][2][21];
assign sum_out[10][2][21] = xor_out[50][2][21] + xor_out[51][2][21] + xor_out[52][2][21] + xor_out[53][2][21] + xor_out[54][2][21];
assign sum_out[11][2][21] = xor_out[55][2][21] + xor_out[56][2][21] + xor_out[57][2][21] + xor_out[58][2][21] + xor_out[59][2][21];
assign sum_out[12][2][21] = xor_out[60][2][21] + xor_out[61][2][21] + xor_out[62][2][21] + xor_out[63][2][21] + xor_out[64][2][21];
assign sum_out[13][2][21] = xor_out[65][2][21] + xor_out[66][2][21] + xor_out[67][2][21] + xor_out[68][2][21] + xor_out[69][2][21];
assign sum_out[14][2][21] = xor_out[70][2][21] + xor_out[71][2][21] + xor_out[72][2][21] + xor_out[73][2][21] + xor_out[74][2][21];
assign sum_out[15][2][21] = xor_out[75][2][21] + xor_out[76][2][21] + xor_out[77][2][21] + xor_out[78][2][21] + xor_out[79][2][21];
assign sum_out[16][2][21] = xor_out[80][2][21] + xor_out[81][2][21] + xor_out[82][2][21] + xor_out[83][2][21] + xor_out[84][2][21];
assign sum_out[17][2][21] = xor_out[85][2][21] + xor_out[86][2][21] + xor_out[87][2][21] + xor_out[88][2][21] + xor_out[89][2][21];
assign sum_out[18][2][21] = xor_out[90][2][21] + xor_out[91][2][21] + xor_out[92][2][21] + xor_out[93][2][21] + xor_out[94][2][21];
assign sum_out[19][2][21] = xor_out[95][2][21] + xor_out[96][2][21] + xor_out[97][2][21] + xor_out[98][2][21] + xor_out[99][2][21];

assign sum_out[0][2][22] = xor_out[0][2][22] + xor_out[1][2][22] + xor_out[2][2][22] + xor_out[3][2][22] + xor_out[4][2][22];
assign sum_out[1][2][22] = xor_out[5][2][22] + xor_out[6][2][22] + xor_out[7][2][22] + xor_out[8][2][22] + xor_out[9][2][22];
assign sum_out[2][2][22] = xor_out[10][2][22] + xor_out[11][2][22] + xor_out[12][2][22] + xor_out[13][2][22] + xor_out[14][2][22];
assign sum_out[3][2][22] = xor_out[15][2][22] + xor_out[16][2][22] + xor_out[17][2][22] + xor_out[18][2][22] + xor_out[19][2][22];
assign sum_out[4][2][22] = xor_out[20][2][22] + xor_out[21][2][22] + xor_out[22][2][22] + xor_out[23][2][22] + xor_out[24][2][22];
assign sum_out[5][2][22] = xor_out[25][2][22] + xor_out[26][2][22] + xor_out[27][2][22] + xor_out[28][2][22] + xor_out[29][2][22];
assign sum_out[6][2][22] = xor_out[30][2][22] + xor_out[31][2][22] + xor_out[32][2][22] + xor_out[33][2][22] + xor_out[34][2][22];
assign sum_out[7][2][22] = xor_out[35][2][22] + xor_out[36][2][22] + xor_out[37][2][22] + xor_out[38][2][22] + xor_out[39][2][22];
assign sum_out[8][2][22] = xor_out[40][2][22] + xor_out[41][2][22] + xor_out[42][2][22] + xor_out[43][2][22] + xor_out[44][2][22];
assign sum_out[9][2][22] = xor_out[45][2][22] + xor_out[46][2][22] + xor_out[47][2][22] + xor_out[48][2][22] + xor_out[49][2][22];
assign sum_out[10][2][22] = xor_out[50][2][22] + xor_out[51][2][22] + xor_out[52][2][22] + xor_out[53][2][22] + xor_out[54][2][22];
assign sum_out[11][2][22] = xor_out[55][2][22] + xor_out[56][2][22] + xor_out[57][2][22] + xor_out[58][2][22] + xor_out[59][2][22];
assign sum_out[12][2][22] = xor_out[60][2][22] + xor_out[61][2][22] + xor_out[62][2][22] + xor_out[63][2][22] + xor_out[64][2][22];
assign sum_out[13][2][22] = xor_out[65][2][22] + xor_out[66][2][22] + xor_out[67][2][22] + xor_out[68][2][22] + xor_out[69][2][22];
assign sum_out[14][2][22] = xor_out[70][2][22] + xor_out[71][2][22] + xor_out[72][2][22] + xor_out[73][2][22] + xor_out[74][2][22];
assign sum_out[15][2][22] = xor_out[75][2][22] + xor_out[76][2][22] + xor_out[77][2][22] + xor_out[78][2][22] + xor_out[79][2][22];
assign sum_out[16][2][22] = xor_out[80][2][22] + xor_out[81][2][22] + xor_out[82][2][22] + xor_out[83][2][22] + xor_out[84][2][22];
assign sum_out[17][2][22] = xor_out[85][2][22] + xor_out[86][2][22] + xor_out[87][2][22] + xor_out[88][2][22] + xor_out[89][2][22];
assign sum_out[18][2][22] = xor_out[90][2][22] + xor_out[91][2][22] + xor_out[92][2][22] + xor_out[93][2][22] + xor_out[94][2][22];
assign sum_out[19][2][22] = xor_out[95][2][22] + xor_out[96][2][22] + xor_out[97][2][22] + xor_out[98][2][22] + xor_out[99][2][22];

assign sum_out[0][2][23] = xor_out[0][2][23] + xor_out[1][2][23] + xor_out[2][2][23] + xor_out[3][2][23] + xor_out[4][2][23];
assign sum_out[1][2][23] = xor_out[5][2][23] + xor_out[6][2][23] + xor_out[7][2][23] + xor_out[8][2][23] + xor_out[9][2][23];
assign sum_out[2][2][23] = xor_out[10][2][23] + xor_out[11][2][23] + xor_out[12][2][23] + xor_out[13][2][23] + xor_out[14][2][23];
assign sum_out[3][2][23] = xor_out[15][2][23] + xor_out[16][2][23] + xor_out[17][2][23] + xor_out[18][2][23] + xor_out[19][2][23];
assign sum_out[4][2][23] = xor_out[20][2][23] + xor_out[21][2][23] + xor_out[22][2][23] + xor_out[23][2][23] + xor_out[24][2][23];
assign sum_out[5][2][23] = xor_out[25][2][23] + xor_out[26][2][23] + xor_out[27][2][23] + xor_out[28][2][23] + xor_out[29][2][23];
assign sum_out[6][2][23] = xor_out[30][2][23] + xor_out[31][2][23] + xor_out[32][2][23] + xor_out[33][2][23] + xor_out[34][2][23];
assign sum_out[7][2][23] = xor_out[35][2][23] + xor_out[36][2][23] + xor_out[37][2][23] + xor_out[38][2][23] + xor_out[39][2][23];
assign sum_out[8][2][23] = xor_out[40][2][23] + xor_out[41][2][23] + xor_out[42][2][23] + xor_out[43][2][23] + xor_out[44][2][23];
assign sum_out[9][2][23] = xor_out[45][2][23] + xor_out[46][2][23] + xor_out[47][2][23] + xor_out[48][2][23] + xor_out[49][2][23];
assign sum_out[10][2][23] = xor_out[50][2][23] + xor_out[51][2][23] + xor_out[52][2][23] + xor_out[53][2][23] + xor_out[54][2][23];
assign sum_out[11][2][23] = xor_out[55][2][23] + xor_out[56][2][23] + xor_out[57][2][23] + xor_out[58][2][23] + xor_out[59][2][23];
assign sum_out[12][2][23] = xor_out[60][2][23] + xor_out[61][2][23] + xor_out[62][2][23] + xor_out[63][2][23] + xor_out[64][2][23];
assign sum_out[13][2][23] = xor_out[65][2][23] + xor_out[66][2][23] + xor_out[67][2][23] + xor_out[68][2][23] + xor_out[69][2][23];
assign sum_out[14][2][23] = xor_out[70][2][23] + xor_out[71][2][23] + xor_out[72][2][23] + xor_out[73][2][23] + xor_out[74][2][23];
assign sum_out[15][2][23] = xor_out[75][2][23] + xor_out[76][2][23] + xor_out[77][2][23] + xor_out[78][2][23] + xor_out[79][2][23];
assign sum_out[16][2][23] = xor_out[80][2][23] + xor_out[81][2][23] + xor_out[82][2][23] + xor_out[83][2][23] + xor_out[84][2][23];
assign sum_out[17][2][23] = xor_out[85][2][23] + xor_out[86][2][23] + xor_out[87][2][23] + xor_out[88][2][23] + xor_out[89][2][23];
assign sum_out[18][2][23] = xor_out[90][2][23] + xor_out[91][2][23] + xor_out[92][2][23] + xor_out[93][2][23] + xor_out[94][2][23];
assign sum_out[19][2][23] = xor_out[95][2][23] + xor_out[96][2][23] + xor_out[97][2][23] + xor_out[98][2][23] + xor_out[99][2][23];

assign sum_out[0][3][0] = xor_out[0][3][0] + xor_out[1][3][0] + xor_out[2][3][0] + xor_out[3][3][0] + xor_out[4][3][0];
assign sum_out[1][3][0] = xor_out[5][3][0] + xor_out[6][3][0] + xor_out[7][3][0] + xor_out[8][3][0] + xor_out[9][3][0];
assign sum_out[2][3][0] = xor_out[10][3][0] + xor_out[11][3][0] + xor_out[12][3][0] + xor_out[13][3][0] + xor_out[14][3][0];
assign sum_out[3][3][0] = xor_out[15][3][0] + xor_out[16][3][0] + xor_out[17][3][0] + xor_out[18][3][0] + xor_out[19][3][0];
assign sum_out[4][3][0] = xor_out[20][3][0] + xor_out[21][3][0] + xor_out[22][3][0] + xor_out[23][3][0] + xor_out[24][3][0];
assign sum_out[5][3][0] = xor_out[25][3][0] + xor_out[26][3][0] + xor_out[27][3][0] + xor_out[28][3][0] + xor_out[29][3][0];
assign sum_out[6][3][0] = xor_out[30][3][0] + xor_out[31][3][0] + xor_out[32][3][0] + xor_out[33][3][0] + xor_out[34][3][0];
assign sum_out[7][3][0] = xor_out[35][3][0] + xor_out[36][3][0] + xor_out[37][3][0] + xor_out[38][3][0] + xor_out[39][3][0];
assign sum_out[8][3][0] = xor_out[40][3][0] + xor_out[41][3][0] + xor_out[42][3][0] + xor_out[43][3][0] + xor_out[44][3][0];
assign sum_out[9][3][0] = xor_out[45][3][0] + xor_out[46][3][0] + xor_out[47][3][0] + xor_out[48][3][0] + xor_out[49][3][0];
assign sum_out[10][3][0] = xor_out[50][3][0] + xor_out[51][3][0] + xor_out[52][3][0] + xor_out[53][3][0] + xor_out[54][3][0];
assign sum_out[11][3][0] = xor_out[55][3][0] + xor_out[56][3][0] + xor_out[57][3][0] + xor_out[58][3][0] + xor_out[59][3][0];
assign sum_out[12][3][0] = xor_out[60][3][0] + xor_out[61][3][0] + xor_out[62][3][0] + xor_out[63][3][0] + xor_out[64][3][0];
assign sum_out[13][3][0] = xor_out[65][3][0] + xor_out[66][3][0] + xor_out[67][3][0] + xor_out[68][3][0] + xor_out[69][3][0];
assign sum_out[14][3][0] = xor_out[70][3][0] + xor_out[71][3][0] + xor_out[72][3][0] + xor_out[73][3][0] + xor_out[74][3][0];
assign sum_out[15][3][0] = xor_out[75][3][0] + xor_out[76][3][0] + xor_out[77][3][0] + xor_out[78][3][0] + xor_out[79][3][0];
assign sum_out[16][3][0] = xor_out[80][3][0] + xor_out[81][3][0] + xor_out[82][3][0] + xor_out[83][3][0] + xor_out[84][3][0];
assign sum_out[17][3][0] = xor_out[85][3][0] + xor_out[86][3][0] + xor_out[87][3][0] + xor_out[88][3][0] + xor_out[89][3][0];
assign sum_out[18][3][0] = xor_out[90][3][0] + xor_out[91][3][0] + xor_out[92][3][0] + xor_out[93][3][0] + xor_out[94][3][0];
assign sum_out[19][3][0] = xor_out[95][3][0] + xor_out[96][3][0] + xor_out[97][3][0] + xor_out[98][3][0] + xor_out[99][3][0];

assign sum_out[0][3][1] = xor_out[0][3][1] + xor_out[1][3][1] + xor_out[2][3][1] + xor_out[3][3][1] + xor_out[4][3][1];
assign sum_out[1][3][1] = xor_out[5][3][1] + xor_out[6][3][1] + xor_out[7][3][1] + xor_out[8][3][1] + xor_out[9][3][1];
assign sum_out[2][3][1] = xor_out[10][3][1] + xor_out[11][3][1] + xor_out[12][3][1] + xor_out[13][3][1] + xor_out[14][3][1];
assign sum_out[3][3][1] = xor_out[15][3][1] + xor_out[16][3][1] + xor_out[17][3][1] + xor_out[18][3][1] + xor_out[19][3][1];
assign sum_out[4][3][1] = xor_out[20][3][1] + xor_out[21][3][1] + xor_out[22][3][1] + xor_out[23][3][1] + xor_out[24][3][1];
assign sum_out[5][3][1] = xor_out[25][3][1] + xor_out[26][3][1] + xor_out[27][3][1] + xor_out[28][3][1] + xor_out[29][3][1];
assign sum_out[6][3][1] = xor_out[30][3][1] + xor_out[31][3][1] + xor_out[32][3][1] + xor_out[33][3][1] + xor_out[34][3][1];
assign sum_out[7][3][1] = xor_out[35][3][1] + xor_out[36][3][1] + xor_out[37][3][1] + xor_out[38][3][1] + xor_out[39][3][1];
assign sum_out[8][3][1] = xor_out[40][3][1] + xor_out[41][3][1] + xor_out[42][3][1] + xor_out[43][3][1] + xor_out[44][3][1];
assign sum_out[9][3][1] = xor_out[45][3][1] + xor_out[46][3][1] + xor_out[47][3][1] + xor_out[48][3][1] + xor_out[49][3][1];
assign sum_out[10][3][1] = xor_out[50][3][1] + xor_out[51][3][1] + xor_out[52][3][1] + xor_out[53][3][1] + xor_out[54][3][1];
assign sum_out[11][3][1] = xor_out[55][3][1] + xor_out[56][3][1] + xor_out[57][3][1] + xor_out[58][3][1] + xor_out[59][3][1];
assign sum_out[12][3][1] = xor_out[60][3][1] + xor_out[61][3][1] + xor_out[62][3][1] + xor_out[63][3][1] + xor_out[64][3][1];
assign sum_out[13][3][1] = xor_out[65][3][1] + xor_out[66][3][1] + xor_out[67][3][1] + xor_out[68][3][1] + xor_out[69][3][1];
assign sum_out[14][3][1] = xor_out[70][3][1] + xor_out[71][3][1] + xor_out[72][3][1] + xor_out[73][3][1] + xor_out[74][3][1];
assign sum_out[15][3][1] = xor_out[75][3][1] + xor_out[76][3][1] + xor_out[77][3][1] + xor_out[78][3][1] + xor_out[79][3][1];
assign sum_out[16][3][1] = xor_out[80][3][1] + xor_out[81][3][1] + xor_out[82][3][1] + xor_out[83][3][1] + xor_out[84][3][1];
assign sum_out[17][3][1] = xor_out[85][3][1] + xor_out[86][3][1] + xor_out[87][3][1] + xor_out[88][3][1] + xor_out[89][3][1];
assign sum_out[18][3][1] = xor_out[90][3][1] + xor_out[91][3][1] + xor_out[92][3][1] + xor_out[93][3][1] + xor_out[94][3][1];
assign sum_out[19][3][1] = xor_out[95][3][1] + xor_out[96][3][1] + xor_out[97][3][1] + xor_out[98][3][1] + xor_out[99][3][1];

assign sum_out[0][3][2] = xor_out[0][3][2] + xor_out[1][3][2] + xor_out[2][3][2] + xor_out[3][3][2] + xor_out[4][3][2];
assign sum_out[1][3][2] = xor_out[5][3][2] + xor_out[6][3][2] + xor_out[7][3][2] + xor_out[8][3][2] + xor_out[9][3][2];
assign sum_out[2][3][2] = xor_out[10][3][2] + xor_out[11][3][2] + xor_out[12][3][2] + xor_out[13][3][2] + xor_out[14][3][2];
assign sum_out[3][3][2] = xor_out[15][3][2] + xor_out[16][3][2] + xor_out[17][3][2] + xor_out[18][3][2] + xor_out[19][3][2];
assign sum_out[4][3][2] = xor_out[20][3][2] + xor_out[21][3][2] + xor_out[22][3][2] + xor_out[23][3][2] + xor_out[24][3][2];
assign sum_out[5][3][2] = xor_out[25][3][2] + xor_out[26][3][2] + xor_out[27][3][2] + xor_out[28][3][2] + xor_out[29][3][2];
assign sum_out[6][3][2] = xor_out[30][3][2] + xor_out[31][3][2] + xor_out[32][3][2] + xor_out[33][3][2] + xor_out[34][3][2];
assign sum_out[7][3][2] = xor_out[35][3][2] + xor_out[36][3][2] + xor_out[37][3][2] + xor_out[38][3][2] + xor_out[39][3][2];
assign sum_out[8][3][2] = xor_out[40][3][2] + xor_out[41][3][2] + xor_out[42][3][2] + xor_out[43][3][2] + xor_out[44][3][2];
assign sum_out[9][3][2] = xor_out[45][3][2] + xor_out[46][3][2] + xor_out[47][3][2] + xor_out[48][3][2] + xor_out[49][3][2];
assign sum_out[10][3][2] = xor_out[50][3][2] + xor_out[51][3][2] + xor_out[52][3][2] + xor_out[53][3][2] + xor_out[54][3][2];
assign sum_out[11][3][2] = xor_out[55][3][2] + xor_out[56][3][2] + xor_out[57][3][2] + xor_out[58][3][2] + xor_out[59][3][2];
assign sum_out[12][3][2] = xor_out[60][3][2] + xor_out[61][3][2] + xor_out[62][3][2] + xor_out[63][3][2] + xor_out[64][3][2];
assign sum_out[13][3][2] = xor_out[65][3][2] + xor_out[66][3][2] + xor_out[67][3][2] + xor_out[68][3][2] + xor_out[69][3][2];
assign sum_out[14][3][2] = xor_out[70][3][2] + xor_out[71][3][2] + xor_out[72][3][2] + xor_out[73][3][2] + xor_out[74][3][2];
assign sum_out[15][3][2] = xor_out[75][3][2] + xor_out[76][3][2] + xor_out[77][3][2] + xor_out[78][3][2] + xor_out[79][3][2];
assign sum_out[16][3][2] = xor_out[80][3][2] + xor_out[81][3][2] + xor_out[82][3][2] + xor_out[83][3][2] + xor_out[84][3][2];
assign sum_out[17][3][2] = xor_out[85][3][2] + xor_out[86][3][2] + xor_out[87][3][2] + xor_out[88][3][2] + xor_out[89][3][2];
assign sum_out[18][3][2] = xor_out[90][3][2] + xor_out[91][3][2] + xor_out[92][3][2] + xor_out[93][3][2] + xor_out[94][3][2];
assign sum_out[19][3][2] = xor_out[95][3][2] + xor_out[96][3][2] + xor_out[97][3][2] + xor_out[98][3][2] + xor_out[99][3][2];

assign sum_out[0][3][3] = xor_out[0][3][3] + xor_out[1][3][3] + xor_out[2][3][3] + xor_out[3][3][3] + xor_out[4][3][3];
assign sum_out[1][3][3] = xor_out[5][3][3] + xor_out[6][3][3] + xor_out[7][3][3] + xor_out[8][3][3] + xor_out[9][3][3];
assign sum_out[2][3][3] = xor_out[10][3][3] + xor_out[11][3][3] + xor_out[12][3][3] + xor_out[13][3][3] + xor_out[14][3][3];
assign sum_out[3][3][3] = xor_out[15][3][3] + xor_out[16][3][3] + xor_out[17][3][3] + xor_out[18][3][3] + xor_out[19][3][3];
assign sum_out[4][3][3] = xor_out[20][3][3] + xor_out[21][3][3] + xor_out[22][3][3] + xor_out[23][3][3] + xor_out[24][3][3];
assign sum_out[5][3][3] = xor_out[25][3][3] + xor_out[26][3][3] + xor_out[27][3][3] + xor_out[28][3][3] + xor_out[29][3][3];
assign sum_out[6][3][3] = xor_out[30][3][3] + xor_out[31][3][3] + xor_out[32][3][3] + xor_out[33][3][3] + xor_out[34][3][3];
assign sum_out[7][3][3] = xor_out[35][3][3] + xor_out[36][3][3] + xor_out[37][3][3] + xor_out[38][3][3] + xor_out[39][3][3];
assign sum_out[8][3][3] = xor_out[40][3][3] + xor_out[41][3][3] + xor_out[42][3][3] + xor_out[43][3][3] + xor_out[44][3][3];
assign sum_out[9][3][3] = xor_out[45][3][3] + xor_out[46][3][3] + xor_out[47][3][3] + xor_out[48][3][3] + xor_out[49][3][3];
assign sum_out[10][3][3] = xor_out[50][3][3] + xor_out[51][3][3] + xor_out[52][3][3] + xor_out[53][3][3] + xor_out[54][3][3];
assign sum_out[11][3][3] = xor_out[55][3][3] + xor_out[56][3][3] + xor_out[57][3][3] + xor_out[58][3][3] + xor_out[59][3][3];
assign sum_out[12][3][3] = xor_out[60][3][3] + xor_out[61][3][3] + xor_out[62][3][3] + xor_out[63][3][3] + xor_out[64][3][3];
assign sum_out[13][3][3] = xor_out[65][3][3] + xor_out[66][3][3] + xor_out[67][3][3] + xor_out[68][3][3] + xor_out[69][3][3];
assign sum_out[14][3][3] = xor_out[70][3][3] + xor_out[71][3][3] + xor_out[72][3][3] + xor_out[73][3][3] + xor_out[74][3][3];
assign sum_out[15][3][3] = xor_out[75][3][3] + xor_out[76][3][3] + xor_out[77][3][3] + xor_out[78][3][3] + xor_out[79][3][3];
assign sum_out[16][3][3] = xor_out[80][3][3] + xor_out[81][3][3] + xor_out[82][3][3] + xor_out[83][3][3] + xor_out[84][3][3];
assign sum_out[17][3][3] = xor_out[85][3][3] + xor_out[86][3][3] + xor_out[87][3][3] + xor_out[88][3][3] + xor_out[89][3][3];
assign sum_out[18][3][3] = xor_out[90][3][3] + xor_out[91][3][3] + xor_out[92][3][3] + xor_out[93][3][3] + xor_out[94][3][3];
assign sum_out[19][3][3] = xor_out[95][3][3] + xor_out[96][3][3] + xor_out[97][3][3] + xor_out[98][3][3] + xor_out[99][3][3];

assign sum_out[0][3][4] = xor_out[0][3][4] + xor_out[1][3][4] + xor_out[2][3][4] + xor_out[3][3][4] + xor_out[4][3][4];
assign sum_out[1][3][4] = xor_out[5][3][4] + xor_out[6][3][4] + xor_out[7][3][4] + xor_out[8][3][4] + xor_out[9][3][4];
assign sum_out[2][3][4] = xor_out[10][3][4] + xor_out[11][3][4] + xor_out[12][3][4] + xor_out[13][3][4] + xor_out[14][3][4];
assign sum_out[3][3][4] = xor_out[15][3][4] + xor_out[16][3][4] + xor_out[17][3][4] + xor_out[18][3][4] + xor_out[19][3][4];
assign sum_out[4][3][4] = xor_out[20][3][4] + xor_out[21][3][4] + xor_out[22][3][4] + xor_out[23][3][4] + xor_out[24][3][4];
assign sum_out[5][3][4] = xor_out[25][3][4] + xor_out[26][3][4] + xor_out[27][3][4] + xor_out[28][3][4] + xor_out[29][3][4];
assign sum_out[6][3][4] = xor_out[30][3][4] + xor_out[31][3][4] + xor_out[32][3][4] + xor_out[33][3][4] + xor_out[34][3][4];
assign sum_out[7][3][4] = xor_out[35][3][4] + xor_out[36][3][4] + xor_out[37][3][4] + xor_out[38][3][4] + xor_out[39][3][4];
assign sum_out[8][3][4] = xor_out[40][3][4] + xor_out[41][3][4] + xor_out[42][3][4] + xor_out[43][3][4] + xor_out[44][3][4];
assign sum_out[9][3][4] = xor_out[45][3][4] + xor_out[46][3][4] + xor_out[47][3][4] + xor_out[48][3][4] + xor_out[49][3][4];
assign sum_out[10][3][4] = xor_out[50][3][4] + xor_out[51][3][4] + xor_out[52][3][4] + xor_out[53][3][4] + xor_out[54][3][4];
assign sum_out[11][3][4] = xor_out[55][3][4] + xor_out[56][3][4] + xor_out[57][3][4] + xor_out[58][3][4] + xor_out[59][3][4];
assign sum_out[12][3][4] = xor_out[60][3][4] + xor_out[61][3][4] + xor_out[62][3][4] + xor_out[63][3][4] + xor_out[64][3][4];
assign sum_out[13][3][4] = xor_out[65][3][4] + xor_out[66][3][4] + xor_out[67][3][4] + xor_out[68][3][4] + xor_out[69][3][4];
assign sum_out[14][3][4] = xor_out[70][3][4] + xor_out[71][3][4] + xor_out[72][3][4] + xor_out[73][3][4] + xor_out[74][3][4];
assign sum_out[15][3][4] = xor_out[75][3][4] + xor_out[76][3][4] + xor_out[77][3][4] + xor_out[78][3][4] + xor_out[79][3][4];
assign sum_out[16][3][4] = xor_out[80][3][4] + xor_out[81][3][4] + xor_out[82][3][4] + xor_out[83][3][4] + xor_out[84][3][4];
assign sum_out[17][3][4] = xor_out[85][3][4] + xor_out[86][3][4] + xor_out[87][3][4] + xor_out[88][3][4] + xor_out[89][3][4];
assign sum_out[18][3][4] = xor_out[90][3][4] + xor_out[91][3][4] + xor_out[92][3][4] + xor_out[93][3][4] + xor_out[94][3][4];
assign sum_out[19][3][4] = xor_out[95][3][4] + xor_out[96][3][4] + xor_out[97][3][4] + xor_out[98][3][4] + xor_out[99][3][4];

assign sum_out[0][3][5] = xor_out[0][3][5] + xor_out[1][3][5] + xor_out[2][3][5] + xor_out[3][3][5] + xor_out[4][3][5];
assign sum_out[1][3][5] = xor_out[5][3][5] + xor_out[6][3][5] + xor_out[7][3][5] + xor_out[8][3][5] + xor_out[9][3][5];
assign sum_out[2][3][5] = xor_out[10][3][5] + xor_out[11][3][5] + xor_out[12][3][5] + xor_out[13][3][5] + xor_out[14][3][5];
assign sum_out[3][3][5] = xor_out[15][3][5] + xor_out[16][3][5] + xor_out[17][3][5] + xor_out[18][3][5] + xor_out[19][3][5];
assign sum_out[4][3][5] = xor_out[20][3][5] + xor_out[21][3][5] + xor_out[22][3][5] + xor_out[23][3][5] + xor_out[24][3][5];
assign sum_out[5][3][5] = xor_out[25][3][5] + xor_out[26][3][5] + xor_out[27][3][5] + xor_out[28][3][5] + xor_out[29][3][5];
assign sum_out[6][3][5] = xor_out[30][3][5] + xor_out[31][3][5] + xor_out[32][3][5] + xor_out[33][3][5] + xor_out[34][3][5];
assign sum_out[7][3][5] = xor_out[35][3][5] + xor_out[36][3][5] + xor_out[37][3][5] + xor_out[38][3][5] + xor_out[39][3][5];
assign sum_out[8][3][5] = xor_out[40][3][5] + xor_out[41][3][5] + xor_out[42][3][5] + xor_out[43][3][5] + xor_out[44][3][5];
assign sum_out[9][3][5] = xor_out[45][3][5] + xor_out[46][3][5] + xor_out[47][3][5] + xor_out[48][3][5] + xor_out[49][3][5];
assign sum_out[10][3][5] = xor_out[50][3][5] + xor_out[51][3][5] + xor_out[52][3][5] + xor_out[53][3][5] + xor_out[54][3][5];
assign sum_out[11][3][5] = xor_out[55][3][5] + xor_out[56][3][5] + xor_out[57][3][5] + xor_out[58][3][5] + xor_out[59][3][5];
assign sum_out[12][3][5] = xor_out[60][3][5] + xor_out[61][3][5] + xor_out[62][3][5] + xor_out[63][3][5] + xor_out[64][3][5];
assign sum_out[13][3][5] = xor_out[65][3][5] + xor_out[66][3][5] + xor_out[67][3][5] + xor_out[68][3][5] + xor_out[69][3][5];
assign sum_out[14][3][5] = xor_out[70][3][5] + xor_out[71][3][5] + xor_out[72][3][5] + xor_out[73][3][5] + xor_out[74][3][5];
assign sum_out[15][3][5] = xor_out[75][3][5] + xor_out[76][3][5] + xor_out[77][3][5] + xor_out[78][3][5] + xor_out[79][3][5];
assign sum_out[16][3][5] = xor_out[80][3][5] + xor_out[81][3][5] + xor_out[82][3][5] + xor_out[83][3][5] + xor_out[84][3][5];
assign sum_out[17][3][5] = xor_out[85][3][5] + xor_out[86][3][5] + xor_out[87][3][5] + xor_out[88][3][5] + xor_out[89][3][5];
assign sum_out[18][3][5] = xor_out[90][3][5] + xor_out[91][3][5] + xor_out[92][3][5] + xor_out[93][3][5] + xor_out[94][3][5];
assign sum_out[19][3][5] = xor_out[95][3][5] + xor_out[96][3][5] + xor_out[97][3][5] + xor_out[98][3][5] + xor_out[99][3][5];

assign sum_out[0][3][6] = xor_out[0][3][6] + xor_out[1][3][6] + xor_out[2][3][6] + xor_out[3][3][6] + xor_out[4][3][6];
assign sum_out[1][3][6] = xor_out[5][3][6] + xor_out[6][3][6] + xor_out[7][3][6] + xor_out[8][3][6] + xor_out[9][3][6];
assign sum_out[2][3][6] = xor_out[10][3][6] + xor_out[11][3][6] + xor_out[12][3][6] + xor_out[13][3][6] + xor_out[14][3][6];
assign sum_out[3][3][6] = xor_out[15][3][6] + xor_out[16][3][6] + xor_out[17][3][6] + xor_out[18][3][6] + xor_out[19][3][6];
assign sum_out[4][3][6] = xor_out[20][3][6] + xor_out[21][3][6] + xor_out[22][3][6] + xor_out[23][3][6] + xor_out[24][3][6];
assign sum_out[5][3][6] = xor_out[25][3][6] + xor_out[26][3][6] + xor_out[27][3][6] + xor_out[28][3][6] + xor_out[29][3][6];
assign sum_out[6][3][6] = xor_out[30][3][6] + xor_out[31][3][6] + xor_out[32][3][6] + xor_out[33][3][6] + xor_out[34][3][6];
assign sum_out[7][3][6] = xor_out[35][3][6] + xor_out[36][3][6] + xor_out[37][3][6] + xor_out[38][3][6] + xor_out[39][3][6];
assign sum_out[8][3][6] = xor_out[40][3][6] + xor_out[41][3][6] + xor_out[42][3][6] + xor_out[43][3][6] + xor_out[44][3][6];
assign sum_out[9][3][6] = xor_out[45][3][6] + xor_out[46][3][6] + xor_out[47][3][6] + xor_out[48][3][6] + xor_out[49][3][6];
assign sum_out[10][3][6] = xor_out[50][3][6] + xor_out[51][3][6] + xor_out[52][3][6] + xor_out[53][3][6] + xor_out[54][3][6];
assign sum_out[11][3][6] = xor_out[55][3][6] + xor_out[56][3][6] + xor_out[57][3][6] + xor_out[58][3][6] + xor_out[59][3][6];
assign sum_out[12][3][6] = xor_out[60][3][6] + xor_out[61][3][6] + xor_out[62][3][6] + xor_out[63][3][6] + xor_out[64][3][6];
assign sum_out[13][3][6] = xor_out[65][3][6] + xor_out[66][3][6] + xor_out[67][3][6] + xor_out[68][3][6] + xor_out[69][3][6];
assign sum_out[14][3][6] = xor_out[70][3][6] + xor_out[71][3][6] + xor_out[72][3][6] + xor_out[73][3][6] + xor_out[74][3][6];
assign sum_out[15][3][6] = xor_out[75][3][6] + xor_out[76][3][6] + xor_out[77][3][6] + xor_out[78][3][6] + xor_out[79][3][6];
assign sum_out[16][3][6] = xor_out[80][3][6] + xor_out[81][3][6] + xor_out[82][3][6] + xor_out[83][3][6] + xor_out[84][3][6];
assign sum_out[17][3][6] = xor_out[85][3][6] + xor_out[86][3][6] + xor_out[87][3][6] + xor_out[88][3][6] + xor_out[89][3][6];
assign sum_out[18][3][6] = xor_out[90][3][6] + xor_out[91][3][6] + xor_out[92][3][6] + xor_out[93][3][6] + xor_out[94][3][6];
assign sum_out[19][3][6] = xor_out[95][3][6] + xor_out[96][3][6] + xor_out[97][3][6] + xor_out[98][3][6] + xor_out[99][3][6];

assign sum_out[0][3][7] = xor_out[0][3][7] + xor_out[1][3][7] + xor_out[2][3][7] + xor_out[3][3][7] + xor_out[4][3][7];
assign sum_out[1][3][7] = xor_out[5][3][7] + xor_out[6][3][7] + xor_out[7][3][7] + xor_out[8][3][7] + xor_out[9][3][7];
assign sum_out[2][3][7] = xor_out[10][3][7] + xor_out[11][3][7] + xor_out[12][3][7] + xor_out[13][3][7] + xor_out[14][3][7];
assign sum_out[3][3][7] = xor_out[15][3][7] + xor_out[16][3][7] + xor_out[17][3][7] + xor_out[18][3][7] + xor_out[19][3][7];
assign sum_out[4][3][7] = xor_out[20][3][7] + xor_out[21][3][7] + xor_out[22][3][7] + xor_out[23][3][7] + xor_out[24][3][7];
assign sum_out[5][3][7] = xor_out[25][3][7] + xor_out[26][3][7] + xor_out[27][3][7] + xor_out[28][3][7] + xor_out[29][3][7];
assign sum_out[6][3][7] = xor_out[30][3][7] + xor_out[31][3][7] + xor_out[32][3][7] + xor_out[33][3][7] + xor_out[34][3][7];
assign sum_out[7][3][7] = xor_out[35][3][7] + xor_out[36][3][7] + xor_out[37][3][7] + xor_out[38][3][7] + xor_out[39][3][7];
assign sum_out[8][3][7] = xor_out[40][3][7] + xor_out[41][3][7] + xor_out[42][3][7] + xor_out[43][3][7] + xor_out[44][3][7];
assign sum_out[9][3][7] = xor_out[45][3][7] + xor_out[46][3][7] + xor_out[47][3][7] + xor_out[48][3][7] + xor_out[49][3][7];
assign sum_out[10][3][7] = xor_out[50][3][7] + xor_out[51][3][7] + xor_out[52][3][7] + xor_out[53][3][7] + xor_out[54][3][7];
assign sum_out[11][3][7] = xor_out[55][3][7] + xor_out[56][3][7] + xor_out[57][3][7] + xor_out[58][3][7] + xor_out[59][3][7];
assign sum_out[12][3][7] = xor_out[60][3][7] + xor_out[61][3][7] + xor_out[62][3][7] + xor_out[63][3][7] + xor_out[64][3][7];
assign sum_out[13][3][7] = xor_out[65][3][7] + xor_out[66][3][7] + xor_out[67][3][7] + xor_out[68][3][7] + xor_out[69][3][7];
assign sum_out[14][3][7] = xor_out[70][3][7] + xor_out[71][3][7] + xor_out[72][3][7] + xor_out[73][3][7] + xor_out[74][3][7];
assign sum_out[15][3][7] = xor_out[75][3][7] + xor_out[76][3][7] + xor_out[77][3][7] + xor_out[78][3][7] + xor_out[79][3][7];
assign sum_out[16][3][7] = xor_out[80][3][7] + xor_out[81][3][7] + xor_out[82][3][7] + xor_out[83][3][7] + xor_out[84][3][7];
assign sum_out[17][3][7] = xor_out[85][3][7] + xor_out[86][3][7] + xor_out[87][3][7] + xor_out[88][3][7] + xor_out[89][3][7];
assign sum_out[18][3][7] = xor_out[90][3][7] + xor_out[91][3][7] + xor_out[92][3][7] + xor_out[93][3][7] + xor_out[94][3][7];
assign sum_out[19][3][7] = xor_out[95][3][7] + xor_out[96][3][7] + xor_out[97][3][7] + xor_out[98][3][7] + xor_out[99][3][7];

assign sum_out[0][3][8] = xor_out[0][3][8] + xor_out[1][3][8] + xor_out[2][3][8] + xor_out[3][3][8] + xor_out[4][3][8];
assign sum_out[1][3][8] = xor_out[5][3][8] + xor_out[6][3][8] + xor_out[7][3][8] + xor_out[8][3][8] + xor_out[9][3][8];
assign sum_out[2][3][8] = xor_out[10][3][8] + xor_out[11][3][8] + xor_out[12][3][8] + xor_out[13][3][8] + xor_out[14][3][8];
assign sum_out[3][3][8] = xor_out[15][3][8] + xor_out[16][3][8] + xor_out[17][3][8] + xor_out[18][3][8] + xor_out[19][3][8];
assign sum_out[4][3][8] = xor_out[20][3][8] + xor_out[21][3][8] + xor_out[22][3][8] + xor_out[23][3][8] + xor_out[24][3][8];
assign sum_out[5][3][8] = xor_out[25][3][8] + xor_out[26][3][8] + xor_out[27][3][8] + xor_out[28][3][8] + xor_out[29][3][8];
assign sum_out[6][3][8] = xor_out[30][3][8] + xor_out[31][3][8] + xor_out[32][3][8] + xor_out[33][3][8] + xor_out[34][3][8];
assign sum_out[7][3][8] = xor_out[35][3][8] + xor_out[36][3][8] + xor_out[37][3][8] + xor_out[38][3][8] + xor_out[39][3][8];
assign sum_out[8][3][8] = xor_out[40][3][8] + xor_out[41][3][8] + xor_out[42][3][8] + xor_out[43][3][8] + xor_out[44][3][8];
assign sum_out[9][3][8] = xor_out[45][3][8] + xor_out[46][3][8] + xor_out[47][3][8] + xor_out[48][3][8] + xor_out[49][3][8];
assign sum_out[10][3][8] = xor_out[50][3][8] + xor_out[51][3][8] + xor_out[52][3][8] + xor_out[53][3][8] + xor_out[54][3][8];
assign sum_out[11][3][8] = xor_out[55][3][8] + xor_out[56][3][8] + xor_out[57][3][8] + xor_out[58][3][8] + xor_out[59][3][8];
assign sum_out[12][3][8] = xor_out[60][3][8] + xor_out[61][3][8] + xor_out[62][3][8] + xor_out[63][3][8] + xor_out[64][3][8];
assign sum_out[13][3][8] = xor_out[65][3][8] + xor_out[66][3][8] + xor_out[67][3][8] + xor_out[68][3][8] + xor_out[69][3][8];
assign sum_out[14][3][8] = xor_out[70][3][8] + xor_out[71][3][8] + xor_out[72][3][8] + xor_out[73][3][8] + xor_out[74][3][8];
assign sum_out[15][3][8] = xor_out[75][3][8] + xor_out[76][3][8] + xor_out[77][3][8] + xor_out[78][3][8] + xor_out[79][3][8];
assign sum_out[16][3][8] = xor_out[80][3][8] + xor_out[81][3][8] + xor_out[82][3][8] + xor_out[83][3][8] + xor_out[84][3][8];
assign sum_out[17][3][8] = xor_out[85][3][8] + xor_out[86][3][8] + xor_out[87][3][8] + xor_out[88][3][8] + xor_out[89][3][8];
assign sum_out[18][3][8] = xor_out[90][3][8] + xor_out[91][3][8] + xor_out[92][3][8] + xor_out[93][3][8] + xor_out[94][3][8];
assign sum_out[19][3][8] = xor_out[95][3][8] + xor_out[96][3][8] + xor_out[97][3][8] + xor_out[98][3][8] + xor_out[99][3][8];

assign sum_out[0][3][9] = xor_out[0][3][9] + xor_out[1][3][9] + xor_out[2][3][9] + xor_out[3][3][9] + xor_out[4][3][9];
assign sum_out[1][3][9] = xor_out[5][3][9] + xor_out[6][3][9] + xor_out[7][3][9] + xor_out[8][3][9] + xor_out[9][3][9];
assign sum_out[2][3][9] = xor_out[10][3][9] + xor_out[11][3][9] + xor_out[12][3][9] + xor_out[13][3][9] + xor_out[14][3][9];
assign sum_out[3][3][9] = xor_out[15][3][9] + xor_out[16][3][9] + xor_out[17][3][9] + xor_out[18][3][9] + xor_out[19][3][9];
assign sum_out[4][3][9] = xor_out[20][3][9] + xor_out[21][3][9] + xor_out[22][3][9] + xor_out[23][3][9] + xor_out[24][3][9];
assign sum_out[5][3][9] = xor_out[25][3][9] + xor_out[26][3][9] + xor_out[27][3][9] + xor_out[28][3][9] + xor_out[29][3][9];
assign sum_out[6][3][9] = xor_out[30][3][9] + xor_out[31][3][9] + xor_out[32][3][9] + xor_out[33][3][9] + xor_out[34][3][9];
assign sum_out[7][3][9] = xor_out[35][3][9] + xor_out[36][3][9] + xor_out[37][3][9] + xor_out[38][3][9] + xor_out[39][3][9];
assign sum_out[8][3][9] = xor_out[40][3][9] + xor_out[41][3][9] + xor_out[42][3][9] + xor_out[43][3][9] + xor_out[44][3][9];
assign sum_out[9][3][9] = xor_out[45][3][9] + xor_out[46][3][9] + xor_out[47][3][9] + xor_out[48][3][9] + xor_out[49][3][9];
assign sum_out[10][3][9] = xor_out[50][3][9] + xor_out[51][3][9] + xor_out[52][3][9] + xor_out[53][3][9] + xor_out[54][3][9];
assign sum_out[11][3][9] = xor_out[55][3][9] + xor_out[56][3][9] + xor_out[57][3][9] + xor_out[58][3][9] + xor_out[59][3][9];
assign sum_out[12][3][9] = xor_out[60][3][9] + xor_out[61][3][9] + xor_out[62][3][9] + xor_out[63][3][9] + xor_out[64][3][9];
assign sum_out[13][3][9] = xor_out[65][3][9] + xor_out[66][3][9] + xor_out[67][3][9] + xor_out[68][3][9] + xor_out[69][3][9];
assign sum_out[14][3][9] = xor_out[70][3][9] + xor_out[71][3][9] + xor_out[72][3][9] + xor_out[73][3][9] + xor_out[74][3][9];
assign sum_out[15][3][9] = xor_out[75][3][9] + xor_out[76][3][9] + xor_out[77][3][9] + xor_out[78][3][9] + xor_out[79][3][9];
assign sum_out[16][3][9] = xor_out[80][3][9] + xor_out[81][3][9] + xor_out[82][3][9] + xor_out[83][3][9] + xor_out[84][3][9];
assign sum_out[17][3][9] = xor_out[85][3][9] + xor_out[86][3][9] + xor_out[87][3][9] + xor_out[88][3][9] + xor_out[89][3][9];
assign sum_out[18][3][9] = xor_out[90][3][9] + xor_out[91][3][9] + xor_out[92][3][9] + xor_out[93][3][9] + xor_out[94][3][9];
assign sum_out[19][3][9] = xor_out[95][3][9] + xor_out[96][3][9] + xor_out[97][3][9] + xor_out[98][3][9] + xor_out[99][3][9];

assign sum_out[0][3][10] = xor_out[0][3][10] + xor_out[1][3][10] + xor_out[2][3][10] + xor_out[3][3][10] + xor_out[4][3][10];
assign sum_out[1][3][10] = xor_out[5][3][10] + xor_out[6][3][10] + xor_out[7][3][10] + xor_out[8][3][10] + xor_out[9][3][10];
assign sum_out[2][3][10] = xor_out[10][3][10] + xor_out[11][3][10] + xor_out[12][3][10] + xor_out[13][3][10] + xor_out[14][3][10];
assign sum_out[3][3][10] = xor_out[15][3][10] + xor_out[16][3][10] + xor_out[17][3][10] + xor_out[18][3][10] + xor_out[19][3][10];
assign sum_out[4][3][10] = xor_out[20][3][10] + xor_out[21][3][10] + xor_out[22][3][10] + xor_out[23][3][10] + xor_out[24][3][10];
assign sum_out[5][3][10] = xor_out[25][3][10] + xor_out[26][3][10] + xor_out[27][3][10] + xor_out[28][3][10] + xor_out[29][3][10];
assign sum_out[6][3][10] = xor_out[30][3][10] + xor_out[31][3][10] + xor_out[32][3][10] + xor_out[33][3][10] + xor_out[34][3][10];
assign sum_out[7][3][10] = xor_out[35][3][10] + xor_out[36][3][10] + xor_out[37][3][10] + xor_out[38][3][10] + xor_out[39][3][10];
assign sum_out[8][3][10] = xor_out[40][3][10] + xor_out[41][3][10] + xor_out[42][3][10] + xor_out[43][3][10] + xor_out[44][3][10];
assign sum_out[9][3][10] = xor_out[45][3][10] + xor_out[46][3][10] + xor_out[47][3][10] + xor_out[48][3][10] + xor_out[49][3][10];
assign sum_out[10][3][10] = xor_out[50][3][10] + xor_out[51][3][10] + xor_out[52][3][10] + xor_out[53][3][10] + xor_out[54][3][10];
assign sum_out[11][3][10] = xor_out[55][3][10] + xor_out[56][3][10] + xor_out[57][3][10] + xor_out[58][3][10] + xor_out[59][3][10];
assign sum_out[12][3][10] = xor_out[60][3][10] + xor_out[61][3][10] + xor_out[62][3][10] + xor_out[63][3][10] + xor_out[64][3][10];
assign sum_out[13][3][10] = xor_out[65][3][10] + xor_out[66][3][10] + xor_out[67][3][10] + xor_out[68][3][10] + xor_out[69][3][10];
assign sum_out[14][3][10] = xor_out[70][3][10] + xor_out[71][3][10] + xor_out[72][3][10] + xor_out[73][3][10] + xor_out[74][3][10];
assign sum_out[15][3][10] = xor_out[75][3][10] + xor_out[76][3][10] + xor_out[77][3][10] + xor_out[78][3][10] + xor_out[79][3][10];
assign sum_out[16][3][10] = xor_out[80][3][10] + xor_out[81][3][10] + xor_out[82][3][10] + xor_out[83][3][10] + xor_out[84][3][10];
assign sum_out[17][3][10] = xor_out[85][3][10] + xor_out[86][3][10] + xor_out[87][3][10] + xor_out[88][3][10] + xor_out[89][3][10];
assign sum_out[18][3][10] = xor_out[90][3][10] + xor_out[91][3][10] + xor_out[92][3][10] + xor_out[93][3][10] + xor_out[94][3][10];
assign sum_out[19][3][10] = xor_out[95][3][10] + xor_out[96][3][10] + xor_out[97][3][10] + xor_out[98][3][10] + xor_out[99][3][10];

assign sum_out[0][3][11] = xor_out[0][3][11] + xor_out[1][3][11] + xor_out[2][3][11] + xor_out[3][3][11] + xor_out[4][3][11];
assign sum_out[1][3][11] = xor_out[5][3][11] + xor_out[6][3][11] + xor_out[7][3][11] + xor_out[8][3][11] + xor_out[9][3][11];
assign sum_out[2][3][11] = xor_out[10][3][11] + xor_out[11][3][11] + xor_out[12][3][11] + xor_out[13][3][11] + xor_out[14][3][11];
assign sum_out[3][3][11] = xor_out[15][3][11] + xor_out[16][3][11] + xor_out[17][3][11] + xor_out[18][3][11] + xor_out[19][3][11];
assign sum_out[4][3][11] = xor_out[20][3][11] + xor_out[21][3][11] + xor_out[22][3][11] + xor_out[23][3][11] + xor_out[24][3][11];
assign sum_out[5][3][11] = xor_out[25][3][11] + xor_out[26][3][11] + xor_out[27][3][11] + xor_out[28][3][11] + xor_out[29][3][11];
assign sum_out[6][3][11] = xor_out[30][3][11] + xor_out[31][3][11] + xor_out[32][3][11] + xor_out[33][3][11] + xor_out[34][3][11];
assign sum_out[7][3][11] = xor_out[35][3][11] + xor_out[36][3][11] + xor_out[37][3][11] + xor_out[38][3][11] + xor_out[39][3][11];
assign sum_out[8][3][11] = xor_out[40][3][11] + xor_out[41][3][11] + xor_out[42][3][11] + xor_out[43][3][11] + xor_out[44][3][11];
assign sum_out[9][3][11] = xor_out[45][3][11] + xor_out[46][3][11] + xor_out[47][3][11] + xor_out[48][3][11] + xor_out[49][3][11];
assign sum_out[10][3][11] = xor_out[50][3][11] + xor_out[51][3][11] + xor_out[52][3][11] + xor_out[53][3][11] + xor_out[54][3][11];
assign sum_out[11][3][11] = xor_out[55][3][11] + xor_out[56][3][11] + xor_out[57][3][11] + xor_out[58][3][11] + xor_out[59][3][11];
assign sum_out[12][3][11] = xor_out[60][3][11] + xor_out[61][3][11] + xor_out[62][3][11] + xor_out[63][3][11] + xor_out[64][3][11];
assign sum_out[13][3][11] = xor_out[65][3][11] + xor_out[66][3][11] + xor_out[67][3][11] + xor_out[68][3][11] + xor_out[69][3][11];
assign sum_out[14][3][11] = xor_out[70][3][11] + xor_out[71][3][11] + xor_out[72][3][11] + xor_out[73][3][11] + xor_out[74][3][11];
assign sum_out[15][3][11] = xor_out[75][3][11] + xor_out[76][3][11] + xor_out[77][3][11] + xor_out[78][3][11] + xor_out[79][3][11];
assign sum_out[16][3][11] = xor_out[80][3][11] + xor_out[81][3][11] + xor_out[82][3][11] + xor_out[83][3][11] + xor_out[84][3][11];
assign sum_out[17][3][11] = xor_out[85][3][11] + xor_out[86][3][11] + xor_out[87][3][11] + xor_out[88][3][11] + xor_out[89][3][11];
assign sum_out[18][3][11] = xor_out[90][3][11] + xor_out[91][3][11] + xor_out[92][3][11] + xor_out[93][3][11] + xor_out[94][3][11];
assign sum_out[19][3][11] = xor_out[95][3][11] + xor_out[96][3][11] + xor_out[97][3][11] + xor_out[98][3][11] + xor_out[99][3][11];

assign sum_out[0][3][12] = xor_out[0][3][12] + xor_out[1][3][12] + xor_out[2][3][12] + xor_out[3][3][12] + xor_out[4][3][12];
assign sum_out[1][3][12] = xor_out[5][3][12] + xor_out[6][3][12] + xor_out[7][3][12] + xor_out[8][3][12] + xor_out[9][3][12];
assign sum_out[2][3][12] = xor_out[10][3][12] + xor_out[11][3][12] + xor_out[12][3][12] + xor_out[13][3][12] + xor_out[14][3][12];
assign sum_out[3][3][12] = xor_out[15][3][12] + xor_out[16][3][12] + xor_out[17][3][12] + xor_out[18][3][12] + xor_out[19][3][12];
assign sum_out[4][3][12] = xor_out[20][3][12] + xor_out[21][3][12] + xor_out[22][3][12] + xor_out[23][3][12] + xor_out[24][3][12];
assign sum_out[5][3][12] = xor_out[25][3][12] + xor_out[26][3][12] + xor_out[27][3][12] + xor_out[28][3][12] + xor_out[29][3][12];
assign sum_out[6][3][12] = xor_out[30][3][12] + xor_out[31][3][12] + xor_out[32][3][12] + xor_out[33][3][12] + xor_out[34][3][12];
assign sum_out[7][3][12] = xor_out[35][3][12] + xor_out[36][3][12] + xor_out[37][3][12] + xor_out[38][3][12] + xor_out[39][3][12];
assign sum_out[8][3][12] = xor_out[40][3][12] + xor_out[41][3][12] + xor_out[42][3][12] + xor_out[43][3][12] + xor_out[44][3][12];
assign sum_out[9][3][12] = xor_out[45][3][12] + xor_out[46][3][12] + xor_out[47][3][12] + xor_out[48][3][12] + xor_out[49][3][12];
assign sum_out[10][3][12] = xor_out[50][3][12] + xor_out[51][3][12] + xor_out[52][3][12] + xor_out[53][3][12] + xor_out[54][3][12];
assign sum_out[11][3][12] = xor_out[55][3][12] + xor_out[56][3][12] + xor_out[57][3][12] + xor_out[58][3][12] + xor_out[59][3][12];
assign sum_out[12][3][12] = xor_out[60][3][12] + xor_out[61][3][12] + xor_out[62][3][12] + xor_out[63][3][12] + xor_out[64][3][12];
assign sum_out[13][3][12] = xor_out[65][3][12] + xor_out[66][3][12] + xor_out[67][3][12] + xor_out[68][3][12] + xor_out[69][3][12];
assign sum_out[14][3][12] = xor_out[70][3][12] + xor_out[71][3][12] + xor_out[72][3][12] + xor_out[73][3][12] + xor_out[74][3][12];
assign sum_out[15][3][12] = xor_out[75][3][12] + xor_out[76][3][12] + xor_out[77][3][12] + xor_out[78][3][12] + xor_out[79][3][12];
assign sum_out[16][3][12] = xor_out[80][3][12] + xor_out[81][3][12] + xor_out[82][3][12] + xor_out[83][3][12] + xor_out[84][3][12];
assign sum_out[17][3][12] = xor_out[85][3][12] + xor_out[86][3][12] + xor_out[87][3][12] + xor_out[88][3][12] + xor_out[89][3][12];
assign sum_out[18][3][12] = xor_out[90][3][12] + xor_out[91][3][12] + xor_out[92][3][12] + xor_out[93][3][12] + xor_out[94][3][12];
assign sum_out[19][3][12] = xor_out[95][3][12] + xor_out[96][3][12] + xor_out[97][3][12] + xor_out[98][3][12] + xor_out[99][3][12];

assign sum_out[0][3][13] = xor_out[0][3][13] + xor_out[1][3][13] + xor_out[2][3][13] + xor_out[3][3][13] + xor_out[4][3][13];
assign sum_out[1][3][13] = xor_out[5][3][13] + xor_out[6][3][13] + xor_out[7][3][13] + xor_out[8][3][13] + xor_out[9][3][13];
assign sum_out[2][3][13] = xor_out[10][3][13] + xor_out[11][3][13] + xor_out[12][3][13] + xor_out[13][3][13] + xor_out[14][3][13];
assign sum_out[3][3][13] = xor_out[15][3][13] + xor_out[16][3][13] + xor_out[17][3][13] + xor_out[18][3][13] + xor_out[19][3][13];
assign sum_out[4][3][13] = xor_out[20][3][13] + xor_out[21][3][13] + xor_out[22][3][13] + xor_out[23][3][13] + xor_out[24][3][13];
assign sum_out[5][3][13] = xor_out[25][3][13] + xor_out[26][3][13] + xor_out[27][3][13] + xor_out[28][3][13] + xor_out[29][3][13];
assign sum_out[6][3][13] = xor_out[30][3][13] + xor_out[31][3][13] + xor_out[32][3][13] + xor_out[33][3][13] + xor_out[34][3][13];
assign sum_out[7][3][13] = xor_out[35][3][13] + xor_out[36][3][13] + xor_out[37][3][13] + xor_out[38][3][13] + xor_out[39][3][13];
assign sum_out[8][3][13] = xor_out[40][3][13] + xor_out[41][3][13] + xor_out[42][3][13] + xor_out[43][3][13] + xor_out[44][3][13];
assign sum_out[9][3][13] = xor_out[45][3][13] + xor_out[46][3][13] + xor_out[47][3][13] + xor_out[48][3][13] + xor_out[49][3][13];
assign sum_out[10][3][13] = xor_out[50][3][13] + xor_out[51][3][13] + xor_out[52][3][13] + xor_out[53][3][13] + xor_out[54][3][13];
assign sum_out[11][3][13] = xor_out[55][3][13] + xor_out[56][3][13] + xor_out[57][3][13] + xor_out[58][3][13] + xor_out[59][3][13];
assign sum_out[12][3][13] = xor_out[60][3][13] + xor_out[61][3][13] + xor_out[62][3][13] + xor_out[63][3][13] + xor_out[64][3][13];
assign sum_out[13][3][13] = xor_out[65][3][13] + xor_out[66][3][13] + xor_out[67][3][13] + xor_out[68][3][13] + xor_out[69][3][13];
assign sum_out[14][3][13] = xor_out[70][3][13] + xor_out[71][3][13] + xor_out[72][3][13] + xor_out[73][3][13] + xor_out[74][3][13];
assign sum_out[15][3][13] = xor_out[75][3][13] + xor_out[76][3][13] + xor_out[77][3][13] + xor_out[78][3][13] + xor_out[79][3][13];
assign sum_out[16][3][13] = xor_out[80][3][13] + xor_out[81][3][13] + xor_out[82][3][13] + xor_out[83][3][13] + xor_out[84][3][13];
assign sum_out[17][3][13] = xor_out[85][3][13] + xor_out[86][3][13] + xor_out[87][3][13] + xor_out[88][3][13] + xor_out[89][3][13];
assign sum_out[18][3][13] = xor_out[90][3][13] + xor_out[91][3][13] + xor_out[92][3][13] + xor_out[93][3][13] + xor_out[94][3][13];
assign sum_out[19][3][13] = xor_out[95][3][13] + xor_out[96][3][13] + xor_out[97][3][13] + xor_out[98][3][13] + xor_out[99][3][13];

assign sum_out[0][3][14] = xor_out[0][3][14] + xor_out[1][3][14] + xor_out[2][3][14] + xor_out[3][3][14] + xor_out[4][3][14];
assign sum_out[1][3][14] = xor_out[5][3][14] + xor_out[6][3][14] + xor_out[7][3][14] + xor_out[8][3][14] + xor_out[9][3][14];
assign sum_out[2][3][14] = xor_out[10][3][14] + xor_out[11][3][14] + xor_out[12][3][14] + xor_out[13][3][14] + xor_out[14][3][14];
assign sum_out[3][3][14] = xor_out[15][3][14] + xor_out[16][3][14] + xor_out[17][3][14] + xor_out[18][3][14] + xor_out[19][3][14];
assign sum_out[4][3][14] = xor_out[20][3][14] + xor_out[21][3][14] + xor_out[22][3][14] + xor_out[23][3][14] + xor_out[24][3][14];
assign sum_out[5][3][14] = xor_out[25][3][14] + xor_out[26][3][14] + xor_out[27][3][14] + xor_out[28][3][14] + xor_out[29][3][14];
assign sum_out[6][3][14] = xor_out[30][3][14] + xor_out[31][3][14] + xor_out[32][3][14] + xor_out[33][3][14] + xor_out[34][3][14];
assign sum_out[7][3][14] = xor_out[35][3][14] + xor_out[36][3][14] + xor_out[37][3][14] + xor_out[38][3][14] + xor_out[39][3][14];
assign sum_out[8][3][14] = xor_out[40][3][14] + xor_out[41][3][14] + xor_out[42][3][14] + xor_out[43][3][14] + xor_out[44][3][14];
assign sum_out[9][3][14] = xor_out[45][3][14] + xor_out[46][3][14] + xor_out[47][3][14] + xor_out[48][3][14] + xor_out[49][3][14];
assign sum_out[10][3][14] = xor_out[50][3][14] + xor_out[51][3][14] + xor_out[52][3][14] + xor_out[53][3][14] + xor_out[54][3][14];
assign sum_out[11][3][14] = xor_out[55][3][14] + xor_out[56][3][14] + xor_out[57][3][14] + xor_out[58][3][14] + xor_out[59][3][14];
assign sum_out[12][3][14] = xor_out[60][3][14] + xor_out[61][3][14] + xor_out[62][3][14] + xor_out[63][3][14] + xor_out[64][3][14];
assign sum_out[13][3][14] = xor_out[65][3][14] + xor_out[66][3][14] + xor_out[67][3][14] + xor_out[68][3][14] + xor_out[69][3][14];
assign sum_out[14][3][14] = xor_out[70][3][14] + xor_out[71][3][14] + xor_out[72][3][14] + xor_out[73][3][14] + xor_out[74][3][14];
assign sum_out[15][3][14] = xor_out[75][3][14] + xor_out[76][3][14] + xor_out[77][3][14] + xor_out[78][3][14] + xor_out[79][3][14];
assign sum_out[16][3][14] = xor_out[80][3][14] + xor_out[81][3][14] + xor_out[82][3][14] + xor_out[83][3][14] + xor_out[84][3][14];
assign sum_out[17][3][14] = xor_out[85][3][14] + xor_out[86][3][14] + xor_out[87][3][14] + xor_out[88][3][14] + xor_out[89][3][14];
assign sum_out[18][3][14] = xor_out[90][3][14] + xor_out[91][3][14] + xor_out[92][3][14] + xor_out[93][3][14] + xor_out[94][3][14];
assign sum_out[19][3][14] = xor_out[95][3][14] + xor_out[96][3][14] + xor_out[97][3][14] + xor_out[98][3][14] + xor_out[99][3][14];

assign sum_out[0][3][15] = xor_out[0][3][15] + xor_out[1][3][15] + xor_out[2][3][15] + xor_out[3][3][15] + xor_out[4][3][15];
assign sum_out[1][3][15] = xor_out[5][3][15] + xor_out[6][3][15] + xor_out[7][3][15] + xor_out[8][3][15] + xor_out[9][3][15];
assign sum_out[2][3][15] = xor_out[10][3][15] + xor_out[11][3][15] + xor_out[12][3][15] + xor_out[13][3][15] + xor_out[14][3][15];
assign sum_out[3][3][15] = xor_out[15][3][15] + xor_out[16][3][15] + xor_out[17][3][15] + xor_out[18][3][15] + xor_out[19][3][15];
assign sum_out[4][3][15] = xor_out[20][3][15] + xor_out[21][3][15] + xor_out[22][3][15] + xor_out[23][3][15] + xor_out[24][3][15];
assign sum_out[5][3][15] = xor_out[25][3][15] + xor_out[26][3][15] + xor_out[27][3][15] + xor_out[28][3][15] + xor_out[29][3][15];
assign sum_out[6][3][15] = xor_out[30][3][15] + xor_out[31][3][15] + xor_out[32][3][15] + xor_out[33][3][15] + xor_out[34][3][15];
assign sum_out[7][3][15] = xor_out[35][3][15] + xor_out[36][3][15] + xor_out[37][3][15] + xor_out[38][3][15] + xor_out[39][3][15];
assign sum_out[8][3][15] = xor_out[40][3][15] + xor_out[41][3][15] + xor_out[42][3][15] + xor_out[43][3][15] + xor_out[44][3][15];
assign sum_out[9][3][15] = xor_out[45][3][15] + xor_out[46][3][15] + xor_out[47][3][15] + xor_out[48][3][15] + xor_out[49][3][15];
assign sum_out[10][3][15] = xor_out[50][3][15] + xor_out[51][3][15] + xor_out[52][3][15] + xor_out[53][3][15] + xor_out[54][3][15];
assign sum_out[11][3][15] = xor_out[55][3][15] + xor_out[56][3][15] + xor_out[57][3][15] + xor_out[58][3][15] + xor_out[59][3][15];
assign sum_out[12][3][15] = xor_out[60][3][15] + xor_out[61][3][15] + xor_out[62][3][15] + xor_out[63][3][15] + xor_out[64][3][15];
assign sum_out[13][3][15] = xor_out[65][3][15] + xor_out[66][3][15] + xor_out[67][3][15] + xor_out[68][3][15] + xor_out[69][3][15];
assign sum_out[14][3][15] = xor_out[70][3][15] + xor_out[71][3][15] + xor_out[72][3][15] + xor_out[73][3][15] + xor_out[74][3][15];
assign sum_out[15][3][15] = xor_out[75][3][15] + xor_out[76][3][15] + xor_out[77][3][15] + xor_out[78][3][15] + xor_out[79][3][15];
assign sum_out[16][3][15] = xor_out[80][3][15] + xor_out[81][3][15] + xor_out[82][3][15] + xor_out[83][3][15] + xor_out[84][3][15];
assign sum_out[17][3][15] = xor_out[85][3][15] + xor_out[86][3][15] + xor_out[87][3][15] + xor_out[88][3][15] + xor_out[89][3][15];
assign sum_out[18][3][15] = xor_out[90][3][15] + xor_out[91][3][15] + xor_out[92][3][15] + xor_out[93][3][15] + xor_out[94][3][15];
assign sum_out[19][3][15] = xor_out[95][3][15] + xor_out[96][3][15] + xor_out[97][3][15] + xor_out[98][3][15] + xor_out[99][3][15];

assign sum_out[0][3][16] = xor_out[0][3][16] + xor_out[1][3][16] + xor_out[2][3][16] + xor_out[3][3][16] + xor_out[4][3][16];
assign sum_out[1][3][16] = xor_out[5][3][16] + xor_out[6][3][16] + xor_out[7][3][16] + xor_out[8][3][16] + xor_out[9][3][16];
assign sum_out[2][3][16] = xor_out[10][3][16] + xor_out[11][3][16] + xor_out[12][3][16] + xor_out[13][3][16] + xor_out[14][3][16];
assign sum_out[3][3][16] = xor_out[15][3][16] + xor_out[16][3][16] + xor_out[17][3][16] + xor_out[18][3][16] + xor_out[19][3][16];
assign sum_out[4][3][16] = xor_out[20][3][16] + xor_out[21][3][16] + xor_out[22][3][16] + xor_out[23][3][16] + xor_out[24][3][16];
assign sum_out[5][3][16] = xor_out[25][3][16] + xor_out[26][3][16] + xor_out[27][3][16] + xor_out[28][3][16] + xor_out[29][3][16];
assign sum_out[6][3][16] = xor_out[30][3][16] + xor_out[31][3][16] + xor_out[32][3][16] + xor_out[33][3][16] + xor_out[34][3][16];
assign sum_out[7][3][16] = xor_out[35][3][16] + xor_out[36][3][16] + xor_out[37][3][16] + xor_out[38][3][16] + xor_out[39][3][16];
assign sum_out[8][3][16] = xor_out[40][3][16] + xor_out[41][3][16] + xor_out[42][3][16] + xor_out[43][3][16] + xor_out[44][3][16];
assign sum_out[9][3][16] = xor_out[45][3][16] + xor_out[46][3][16] + xor_out[47][3][16] + xor_out[48][3][16] + xor_out[49][3][16];
assign sum_out[10][3][16] = xor_out[50][3][16] + xor_out[51][3][16] + xor_out[52][3][16] + xor_out[53][3][16] + xor_out[54][3][16];
assign sum_out[11][3][16] = xor_out[55][3][16] + xor_out[56][3][16] + xor_out[57][3][16] + xor_out[58][3][16] + xor_out[59][3][16];
assign sum_out[12][3][16] = xor_out[60][3][16] + xor_out[61][3][16] + xor_out[62][3][16] + xor_out[63][3][16] + xor_out[64][3][16];
assign sum_out[13][3][16] = xor_out[65][3][16] + xor_out[66][3][16] + xor_out[67][3][16] + xor_out[68][3][16] + xor_out[69][3][16];
assign sum_out[14][3][16] = xor_out[70][3][16] + xor_out[71][3][16] + xor_out[72][3][16] + xor_out[73][3][16] + xor_out[74][3][16];
assign sum_out[15][3][16] = xor_out[75][3][16] + xor_out[76][3][16] + xor_out[77][3][16] + xor_out[78][3][16] + xor_out[79][3][16];
assign sum_out[16][3][16] = xor_out[80][3][16] + xor_out[81][3][16] + xor_out[82][3][16] + xor_out[83][3][16] + xor_out[84][3][16];
assign sum_out[17][3][16] = xor_out[85][3][16] + xor_out[86][3][16] + xor_out[87][3][16] + xor_out[88][3][16] + xor_out[89][3][16];
assign sum_out[18][3][16] = xor_out[90][3][16] + xor_out[91][3][16] + xor_out[92][3][16] + xor_out[93][3][16] + xor_out[94][3][16];
assign sum_out[19][3][16] = xor_out[95][3][16] + xor_out[96][3][16] + xor_out[97][3][16] + xor_out[98][3][16] + xor_out[99][3][16];

assign sum_out[0][3][17] = xor_out[0][3][17] + xor_out[1][3][17] + xor_out[2][3][17] + xor_out[3][3][17] + xor_out[4][3][17];
assign sum_out[1][3][17] = xor_out[5][3][17] + xor_out[6][3][17] + xor_out[7][3][17] + xor_out[8][3][17] + xor_out[9][3][17];
assign sum_out[2][3][17] = xor_out[10][3][17] + xor_out[11][3][17] + xor_out[12][3][17] + xor_out[13][3][17] + xor_out[14][3][17];
assign sum_out[3][3][17] = xor_out[15][3][17] + xor_out[16][3][17] + xor_out[17][3][17] + xor_out[18][3][17] + xor_out[19][3][17];
assign sum_out[4][3][17] = xor_out[20][3][17] + xor_out[21][3][17] + xor_out[22][3][17] + xor_out[23][3][17] + xor_out[24][3][17];
assign sum_out[5][3][17] = xor_out[25][3][17] + xor_out[26][3][17] + xor_out[27][3][17] + xor_out[28][3][17] + xor_out[29][3][17];
assign sum_out[6][3][17] = xor_out[30][3][17] + xor_out[31][3][17] + xor_out[32][3][17] + xor_out[33][3][17] + xor_out[34][3][17];
assign sum_out[7][3][17] = xor_out[35][3][17] + xor_out[36][3][17] + xor_out[37][3][17] + xor_out[38][3][17] + xor_out[39][3][17];
assign sum_out[8][3][17] = xor_out[40][3][17] + xor_out[41][3][17] + xor_out[42][3][17] + xor_out[43][3][17] + xor_out[44][3][17];
assign sum_out[9][3][17] = xor_out[45][3][17] + xor_out[46][3][17] + xor_out[47][3][17] + xor_out[48][3][17] + xor_out[49][3][17];
assign sum_out[10][3][17] = xor_out[50][3][17] + xor_out[51][3][17] + xor_out[52][3][17] + xor_out[53][3][17] + xor_out[54][3][17];
assign sum_out[11][3][17] = xor_out[55][3][17] + xor_out[56][3][17] + xor_out[57][3][17] + xor_out[58][3][17] + xor_out[59][3][17];
assign sum_out[12][3][17] = xor_out[60][3][17] + xor_out[61][3][17] + xor_out[62][3][17] + xor_out[63][3][17] + xor_out[64][3][17];
assign sum_out[13][3][17] = xor_out[65][3][17] + xor_out[66][3][17] + xor_out[67][3][17] + xor_out[68][3][17] + xor_out[69][3][17];
assign sum_out[14][3][17] = xor_out[70][3][17] + xor_out[71][3][17] + xor_out[72][3][17] + xor_out[73][3][17] + xor_out[74][3][17];
assign sum_out[15][3][17] = xor_out[75][3][17] + xor_out[76][3][17] + xor_out[77][3][17] + xor_out[78][3][17] + xor_out[79][3][17];
assign sum_out[16][3][17] = xor_out[80][3][17] + xor_out[81][3][17] + xor_out[82][3][17] + xor_out[83][3][17] + xor_out[84][3][17];
assign sum_out[17][3][17] = xor_out[85][3][17] + xor_out[86][3][17] + xor_out[87][3][17] + xor_out[88][3][17] + xor_out[89][3][17];
assign sum_out[18][3][17] = xor_out[90][3][17] + xor_out[91][3][17] + xor_out[92][3][17] + xor_out[93][3][17] + xor_out[94][3][17];
assign sum_out[19][3][17] = xor_out[95][3][17] + xor_out[96][3][17] + xor_out[97][3][17] + xor_out[98][3][17] + xor_out[99][3][17];

assign sum_out[0][3][18] = xor_out[0][3][18] + xor_out[1][3][18] + xor_out[2][3][18] + xor_out[3][3][18] + xor_out[4][3][18];
assign sum_out[1][3][18] = xor_out[5][3][18] + xor_out[6][3][18] + xor_out[7][3][18] + xor_out[8][3][18] + xor_out[9][3][18];
assign sum_out[2][3][18] = xor_out[10][3][18] + xor_out[11][3][18] + xor_out[12][3][18] + xor_out[13][3][18] + xor_out[14][3][18];
assign sum_out[3][3][18] = xor_out[15][3][18] + xor_out[16][3][18] + xor_out[17][3][18] + xor_out[18][3][18] + xor_out[19][3][18];
assign sum_out[4][3][18] = xor_out[20][3][18] + xor_out[21][3][18] + xor_out[22][3][18] + xor_out[23][3][18] + xor_out[24][3][18];
assign sum_out[5][3][18] = xor_out[25][3][18] + xor_out[26][3][18] + xor_out[27][3][18] + xor_out[28][3][18] + xor_out[29][3][18];
assign sum_out[6][3][18] = xor_out[30][3][18] + xor_out[31][3][18] + xor_out[32][3][18] + xor_out[33][3][18] + xor_out[34][3][18];
assign sum_out[7][3][18] = xor_out[35][3][18] + xor_out[36][3][18] + xor_out[37][3][18] + xor_out[38][3][18] + xor_out[39][3][18];
assign sum_out[8][3][18] = xor_out[40][3][18] + xor_out[41][3][18] + xor_out[42][3][18] + xor_out[43][3][18] + xor_out[44][3][18];
assign sum_out[9][3][18] = xor_out[45][3][18] + xor_out[46][3][18] + xor_out[47][3][18] + xor_out[48][3][18] + xor_out[49][3][18];
assign sum_out[10][3][18] = xor_out[50][3][18] + xor_out[51][3][18] + xor_out[52][3][18] + xor_out[53][3][18] + xor_out[54][3][18];
assign sum_out[11][3][18] = xor_out[55][3][18] + xor_out[56][3][18] + xor_out[57][3][18] + xor_out[58][3][18] + xor_out[59][3][18];
assign sum_out[12][3][18] = xor_out[60][3][18] + xor_out[61][3][18] + xor_out[62][3][18] + xor_out[63][3][18] + xor_out[64][3][18];
assign sum_out[13][3][18] = xor_out[65][3][18] + xor_out[66][3][18] + xor_out[67][3][18] + xor_out[68][3][18] + xor_out[69][3][18];
assign sum_out[14][3][18] = xor_out[70][3][18] + xor_out[71][3][18] + xor_out[72][3][18] + xor_out[73][3][18] + xor_out[74][3][18];
assign sum_out[15][3][18] = xor_out[75][3][18] + xor_out[76][3][18] + xor_out[77][3][18] + xor_out[78][3][18] + xor_out[79][3][18];
assign sum_out[16][3][18] = xor_out[80][3][18] + xor_out[81][3][18] + xor_out[82][3][18] + xor_out[83][3][18] + xor_out[84][3][18];
assign sum_out[17][3][18] = xor_out[85][3][18] + xor_out[86][3][18] + xor_out[87][3][18] + xor_out[88][3][18] + xor_out[89][3][18];
assign sum_out[18][3][18] = xor_out[90][3][18] + xor_out[91][3][18] + xor_out[92][3][18] + xor_out[93][3][18] + xor_out[94][3][18];
assign sum_out[19][3][18] = xor_out[95][3][18] + xor_out[96][3][18] + xor_out[97][3][18] + xor_out[98][3][18] + xor_out[99][3][18];

assign sum_out[0][3][19] = xor_out[0][3][19] + xor_out[1][3][19] + xor_out[2][3][19] + xor_out[3][3][19] + xor_out[4][3][19];
assign sum_out[1][3][19] = xor_out[5][3][19] + xor_out[6][3][19] + xor_out[7][3][19] + xor_out[8][3][19] + xor_out[9][3][19];
assign sum_out[2][3][19] = xor_out[10][3][19] + xor_out[11][3][19] + xor_out[12][3][19] + xor_out[13][3][19] + xor_out[14][3][19];
assign sum_out[3][3][19] = xor_out[15][3][19] + xor_out[16][3][19] + xor_out[17][3][19] + xor_out[18][3][19] + xor_out[19][3][19];
assign sum_out[4][3][19] = xor_out[20][3][19] + xor_out[21][3][19] + xor_out[22][3][19] + xor_out[23][3][19] + xor_out[24][3][19];
assign sum_out[5][3][19] = xor_out[25][3][19] + xor_out[26][3][19] + xor_out[27][3][19] + xor_out[28][3][19] + xor_out[29][3][19];
assign sum_out[6][3][19] = xor_out[30][3][19] + xor_out[31][3][19] + xor_out[32][3][19] + xor_out[33][3][19] + xor_out[34][3][19];
assign sum_out[7][3][19] = xor_out[35][3][19] + xor_out[36][3][19] + xor_out[37][3][19] + xor_out[38][3][19] + xor_out[39][3][19];
assign sum_out[8][3][19] = xor_out[40][3][19] + xor_out[41][3][19] + xor_out[42][3][19] + xor_out[43][3][19] + xor_out[44][3][19];
assign sum_out[9][3][19] = xor_out[45][3][19] + xor_out[46][3][19] + xor_out[47][3][19] + xor_out[48][3][19] + xor_out[49][3][19];
assign sum_out[10][3][19] = xor_out[50][3][19] + xor_out[51][3][19] + xor_out[52][3][19] + xor_out[53][3][19] + xor_out[54][3][19];
assign sum_out[11][3][19] = xor_out[55][3][19] + xor_out[56][3][19] + xor_out[57][3][19] + xor_out[58][3][19] + xor_out[59][3][19];
assign sum_out[12][3][19] = xor_out[60][3][19] + xor_out[61][3][19] + xor_out[62][3][19] + xor_out[63][3][19] + xor_out[64][3][19];
assign sum_out[13][3][19] = xor_out[65][3][19] + xor_out[66][3][19] + xor_out[67][3][19] + xor_out[68][3][19] + xor_out[69][3][19];
assign sum_out[14][3][19] = xor_out[70][3][19] + xor_out[71][3][19] + xor_out[72][3][19] + xor_out[73][3][19] + xor_out[74][3][19];
assign sum_out[15][3][19] = xor_out[75][3][19] + xor_out[76][3][19] + xor_out[77][3][19] + xor_out[78][3][19] + xor_out[79][3][19];
assign sum_out[16][3][19] = xor_out[80][3][19] + xor_out[81][3][19] + xor_out[82][3][19] + xor_out[83][3][19] + xor_out[84][3][19];
assign sum_out[17][3][19] = xor_out[85][3][19] + xor_out[86][3][19] + xor_out[87][3][19] + xor_out[88][3][19] + xor_out[89][3][19];
assign sum_out[18][3][19] = xor_out[90][3][19] + xor_out[91][3][19] + xor_out[92][3][19] + xor_out[93][3][19] + xor_out[94][3][19];
assign sum_out[19][3][19] = xor_out[95][3][19] + xor_out[96][3][19] + xor_out[97][3][19] + xor_out[98][3][19] + xor_out[99][3][19];

assign sum_out[0][3][20] = xor_out[0][3][20] + xor_out[1][3][20] + xor_out[2][3][20] + xor_out[3][3][20] + xor_out[4][3][20];
assign sum_out[1][3][20] = xor_out[5][3][20] + xor_out[6][3][20] + xor_out[7][3][20] + xor_out[8][3][20] + xor_out[9][3][20];
assign sum_out[2][3][20] = xor_out[10][3][20] + xor_out[11][3][20] + xor_out[12][3][20] + xor_out[13][3][20] + xor_out[14][3][20];
assign sum_out[3][3][20] = xor_out[15][3][20] + xor_out[16][3][20] + xor_out[17][3][20] + xor_out[18][3][20] + xor_out[19][3][20];
assign sum_out[4][3][20] = xor_out[20][3][20] + xor_out[21][3][20] + xor_out[22][3][20] + xor_out[23][3][20] + xor_out[24][3][20];
assign sum_out[5][3][20] = xor_out[25][3][20] + xor_out[26][3][20] + xor_out[27][3][20] + xor_out[28][3][20] + xor_out[29][3][20];
assign sum_out[6][3][20] = xor_out[30][3][20] + xor_out[31][3][20] + xor_out[32][3][20] + xor_out[33][3][20] + xor_out[34][3][20];
assign sum_out[7][3][20] = xor_out[35][3][20] + xor_out[36][3][20] + xor_out[37][3][20] + xor_out[38][3][20] + xor_out[39][3][20];
assign sum_out[8][3][20] = xor_out[40][3][20] + xor_out[41][3][20] + xor_out[42][3][20] + xor_out[43][3][20] + xor_out[44][3][20];
assign sum_out[9][3][20] = xor_out[45][3][20] + xor_out[46][3][20] + xor_out[47][3][20] + xor_out[48][3][20] + xor_out[49][3][20];
assign sum_out[10][3][20] = xor_out[50][3][20] + xor_out[51][3][20] + xor_out[52][3][20] + xor_out[53][3][20] + xor_out[54][3][20];
assign sum_out[11][3][20] = xor_out[55][3][20] + xor_out[56][3][20] + xor_out[57][3][20] + xor_out[58][3][20] + xor_out[59][3][20];
assign sum_out[12][3][20] = xor_out[60][3][20] + xor_out[61][3][20] + xor_out[62][3][20] + xor_out[63][3][20] + xor_out[64][3][20];
assign sum_out[13][3][20] = xor_out[65][3][20] + xor_out[66][3][20] + xor_out[67][3][20] + xor_out[68][3][20] + xor_out[69][3][20];
assign sum_out[14][3][20] = xor_out[70][3][20] + xor_out[71][3][20] + xor_out[72][3][20] + xor_out[73][3][20] + xor_out[74][3][20];
assign sum_out[15][3][20] = xor_out[75][3][20] + xor_out[76][3][20] + xor_out[77][3][20] + xor_out[78][3][20] + xor_out[79][3][20];
assign sum_out[16][3][20] = xor_out[80][3][20] + xor_out[81][3][20] + xor_out[82][3][20] + xor_out[83][3][20] + xor_out[84][3][20];
assign sum_out[17][3][20] = xor_out[85][3][20] + xor_out[86][3][20] + xor_out[87][3][20] + xor_out[88][3][20] + xor_out[89][3][20];
assign sum_out[18][3][20] = xor_out[90][3][20] + xor_out[91][3][20] + xor_out[92][3][20] + xor_out[93][3][20] + xor_out[94][3][20];
assign sum_out[19][3][20] = xor_out[95][3][20] + xor_out[96][3][20] + xor_out[97][3][20] + xor_out[98][3][20] + xor_out[99][3][20];

assign sum_out[0][3][21] = xor_out[0][3][21] + xor_out[1][3][21] + xor_out[2][3][21] + xor_out[3][3][21] + xor_out[4][3][21];
assign sum_out[1][3][21] = xor_out[5][3][21] + xor_out[6][3][21] + xor_out[7][3][21] + xor_out[8][3][21] + xor_out[9][3][21];
assign sum_out[2][3][21] = xor_out[10][3][21] + xor_out[11][3][21] + xor_out[12][3][21] + xor_out[13][3][21] + xor_out[14][3][21];
assign sum_out[3][3][21] = xor_out[15][3][21] + xor_out[16][3][21] + xor_out[17][3][21] + xor_out[18][3][21] + xor_out[19][3][21];
assign sum_out[4][3][21] = xor_out[20][3][21] + xor_out[21][3][21] + xor_out[22][3][21] + xor_out[23][3][21] + xor_out[24][3][21];
assign sum_out[5][3][21] = xor_out[25][3][21] + xor_out[26][3][21] + xor_out[27][3][21] + xor_out[28][3][21] + xor_out[29][3][21];
assign sum_out[6][3][21] = xor_out[30][3][21] + xor_out[31][3][21] + xor_out[32][3][21] + xor_out[33][3][21] + xor_out[34][3][21];
assign sum_out[7][3][21] = xor_out[35][3][21] + xor_out[36][3][21] + xor_out[37][3][21] + xor_out[38][3][21] + xor_out[39][3][21];
assign sum_out[8][3][21] = xor_out[40][3][21] + xor_out[41][3][21] + xor_out[42][3][21] + xor_out[43][3][21] + xor_out[44][3][21];
assign sum_out[9][3][21] = xor_out[45][3][21] + xor_out[46][3][21] + xor_out[47][3][21] + xor_out[48][3][21] + xor_out[49][3][21];
assign sum_out[10][3][21] = xor_out[50][3][21] + xor_out[51][3][21] + xor_out[52][3][21] + xor_out[53][3][21] + xor_out[54][3][21];
assign sum_out[11][3][21] = xor_out[55][3][21] + xor_out[56][3][21] + xor_out[57][3][21] + xor_out[58][3][21] + xor_out[59][3][21];
assign sum_out[12][3][21] = xor_out[60][3][21] + xor_out[61][3][21] + xor_out[62][3][21] + xor_out[63][3][21] + xor_out[64][3][21];
assign sum_out[13][3][21] = xor_out[65][3][21] + xor_out[66][3][21] + xor_out[67][3][21] + xor_out[68][3][21] + xor_out[69][3][21];
assign sum_out[14][3][21] = xor_out[70][3][21] + xor_out[71][3][21] + xor_out[72][3][21] + xor_out[73][3][21] + xor_out[74][3][21];
assign sum_out[15][3][21] = xor_out[75][3][21] + xor_out[76][3][21] + xor_out[77][3][21] + xor_out[78][3][21] + xor_out[79][3][21];
assign sum_out[16][3][21] = xor_out[80][3][21] + xor_out[81][3][21] + xor_out[82][3][21] + xor_out[83][3][21] + xor_out[84][3][21];
assign sum_out[17][3][21] = xor_out[85][3][21] + xor_out[86][3][21] + xor_out[87][3][21] + xor_out[88][3][21] + xor_out[89][3][21];
assign sum_out[18][3][21] = xor_out[90][3][21] + xor_out[91][3][21] + xor_out[92][3][21] + xor_out[93][3][21] + xor_out[94][3][21];
assign sum_out[19][3][21] = xor_out[95][3][21] + xor_out[96][3][21] + xor_out[97][3][21] + xor_out[98][3][21] + xor_out[99][3][21];

assign sum_out[0][3][22] = xor_out[0][3][22] + xor_out[1][3][22] + xor_out[2][3][22] + xor_out[3][3][22] + xor_out[4][3][22];
assign sum_out[1][3][22] = xor_out[5][3][22] + xor_out[6][3][22] + xor_out[7][3][22] + xor_out[8][3][22] + xor_out[9][3][22];
assign sum_out[2][3][22] = xor_out[10][3][22] + xor_out[11][3][22] + xor_out[12][3][22] + xor_out[13][3][22] + xor_out[14][3][22];
assign sum_out[3][3][22] = xor_out[15][3][22] + xor_out[16][3][22] + xor_out[17][3][22] + xor_out[18][3][22] + xor_out[19][3][22];
assign sum_out[4][3][22] = xor_out[20][3][22] + xor_out[21][3][22] + xor_out[22][3][22] + xor_out[23][3][22] + xor_out[24][3][22];
assign sum_out[5][3][22] = xor_out[25][3][22] + xor_out[26][3][22] + xor_out[27][3][22] + xor_out[28][3][22] + xor_out[29][3][22];
assign sum_out[6][3][22] = xor_out[30][3][22] + xor_out[31][3][22] + xor_out[32][3][22] + xor_out[33][3][22] + xor_out[34][3][22];
assign sum_out[7][3][22] = xor_out[35][3][22] + xor_out[36][3][22] + xor_out[37][3][22] + xor_out[38][3][22] + xor_out[39][3][22];
assign sum_out[8][3][22] = xor_out[40][3][22] + xor_out[41][3][22] + xor_out[42][3][22] + xor_out[43][3][22] + xor_out[44][3][22];
assign sum_out[9][3][22] = xor_out[45][3][22] + xor_out[46][3][22] + xor_out[47][3][22] + xor_out[48][3][22] + xor_out[49][3][22];
assign sum_out[10][3][22] = xor_out[50][3][22] + xor_out[51][3][22] + xor_out[52][3][22] + xor_out[53][3][22] + xor_out[54][3][22];
assign sum_out[11][3][22] = xor_out[55][3][22] + xor_out[56][3][22] + xor_out[57][3][22] + xor_out[58][3][22] + xor_out[59][3][22];
assign sum_out[12][3][22] = xor_out[60][3][22] + xor_out[61][3][22] + xor_out[62][3][22] + xor_out[63][3][22] + xor_out[64][3][22];
assign sum_out[13][3][22] = xor_out[65][3][22] + xor_out[66][3][22] + xor_out[67][3][22] + xor_out[68][3][22] + xor_out[69][3][22];
assign sum_out[14][3][22] = xor_out[70][3][22] + xor_out[71][3][22] + xor_out[72][3][22] + xor_out[73][3][22] + xor_out[74][3][22];
assign sum_out[15][3][22] = xor_out[75][3][22] + xor_out[76][3][22] + xor_out[77][3][22] + xor_out[78][3][22] + xor_out[79][3][22];
assign sum_out[16][3][22] = xor_out[80][3][22] + xor_out[81][3][22] + xor_out[82][3][22] + xor_out[83][3][22] + xor_out[84][3][22];
assign sum_out[17][3][22] = xor_out[85][3][22] + xor_out[86][3][22] + xor_out[87][3][22] + xor_out[88][3][22] + xor_out[89][3][22];
assign sum_out[18][3][22] = xor_out[90][3][22] + xor_out[91][3][22] + xor_out[92][3][22] + xor_out[93][3][22] + xor_out[94][3][22];
assign sum_out[19][3][22] = xor_out[95][3][22] + xor_out[96][3][22] + xor_out[97][3][22] + xor_out[98][3][22] + xor_out[99][3][22];

assign sum_out[0][3][23] = xor_out[0][3][23] + xor_out[1][3][23] + xor_out[2][3][23] + xor_out[3][3][23] + xor_out[4][3][23];
assign sum_out[1][3][23] = xor_out[5][3][23] + xor_out[6][3][23] + xor_out[7][3][23] + xor_out[8][3][23] + xor_out[9][3][23];
assign sum_out[2][3][23] = xor_out[10][3][23] + xor_out[11][3][23] + xor_out[12][3][23] + xor_out[13][3][23] + xor_out[14][3][23];
assign sum_out[3][3][23] = xor_out[15][3][23] + xor_out[16][3][23] + xor_out[17][3][23] + xor_out[18][3][23] + xor_out[19][3][23];
assign sum_out[4][3][23] = xor_out[20][3][23] + xor_out[21][3][23] + xor_out[22][3][23] + xor_out[23][3][23] + xor_out[24][3][23];
assign sum_out[5][3][23] = xor_out[25][3][23] + xor_out[26][3][23] + xor_out[27][3][23] + xor_out[28][3][23] + xor_out[29][3][23];
assign sum_out[6][3][23] = xor_out[30][3][23] + xor_out[31][3][23] + xor_out[32][3][23] + xor_out[33][3][23] + xor_out[34][3][23];
assign sum_out[7][3][23] = xor_out[35][3][23] + xor_out[36][3][23] + xor_out[37][3][23] + xor_out[38][3][23] + xor_out[39][3][23];
assign sum_out[8][3][23] = xor_out[40][3][23] + xor_out[41][3][23] + xor_out[42][3][23] + xor_out[43][3][23] + xor_out[44][3][23];
assign sum_out[9][3][23] = xor_out[45][3][23] + xor_out[46][3][23] + xor_out[47][3][23] + xor_out[48][3][23] + xor_out[49][3][23];
assign sum_out[10][3][23] = xor_out[50][3][23] + xor_out[51][3][23] + xor_out[52][3][23] + xor_out[53][3][23] + xor_out[54][3][23];
assign sum_out[11][3][23] = xor_out[55][3][23] + xor_out[56][3][23] + xor_out[57][3][23] + xor_out[58][3][23] + xor_out[59][3][23];
assign sum_out[12][3][23] = xor_out[60][3][23] + xor_out[61][3][23] + xor_out[62][3][23] + xor_out[63][3][23] + xor_out[64][3][23];
assign sum_out[13][3][23] = xor_out[65][3][23] + xor_out[66][3][23] + xor_out[67][3][23] + xor_out[68][3][23] + xor_out[69][3][23];
assign sum_out[14][3][23] = xor_out[70][3][23] + xor_out[71][3][23] + xor_out[72][3][23] + xor_out[73][3][23] + xor_out[74][3][23];
assign sum_out[15][3][23] = xor_out[75][3][23] + xor_out[76][3][23] + xor_out[77][3][23] + xor_out[78][3][23] + xor_out[79][3][23];
assign sum_out[16][3][23] = xor_out[80][3][23] + xor_out[81][3][23] + xor_out[82][3][23] + xor_out[83][3][23] + xor_out[84][3][23];
assign sum_out[17][3][23] = xor_out[85][3][23] + xor_out[86][3][23] + xor_out[87][3][23] + xor_out[88][3][23] + xor_out[89][3][23];
assign sum_out[18][3][23] = xor_out[90][3][23] + xor_out[91][3][23] + xor_out[92][3][23] + xor_out[93][3][23] + xor_out[94][3][23];
assign sum_out[19][3][23] = xor_out[95][3][23] + xor_out[96][3][23] + xor_out[97][3][23] + xor_out[98][3][23] + xor_out[99][3][23];

assign sum_out[0][4][0] = xor_out[0][4][0] + xor_out[1][4][0] + xor_out[2][4][0] + xor_out[3][4][0] + xor_out[4][4][0];
assign sum_out[1][4][0] = xor_out[5][4][0] + xor_out[6][4][0] + xor_out[7][4][0] + xor_out[8][4][0] + xor_out[9][4][0];
assign sum_out[2][4][0] = xor_out[10][4][0] + xor_out[11][4][0] + xor_out[12][4][0] + xor_out[13][4][0] + xor_out[14][4][0];
assign sum_out[3][4][0] = xor_out[15][4][0] + xor_out[16][4][0] + xor_out[17][4][0] + xor_out[18][4][0] + xor_out[19][4][0];
assign sum_out[4][4][0] = xor_out[20][4][0] + xor_out[21][4][0] + xor_out[22][4][0] + xor_out[23][4][0] + xor_out[24][4][0];
assign sum_out[5][4][0] = xor_out[25][4][0] + xor_out[26][4][0] + xor_out[27][4][0] + xor_out[28][4][0] + xor_out[29][4][0];
assign sum_out[6][4][0] = xor_out[30][4][0] + xor_out[31][4][0] + xor_out[32][4][0] + xor_out[33][4][0] + xor_out[34][4][0];
assign sum_out[7][4][0] = xor_out[35][4][0] + xor_out[36][4][0] + xor_out[37][4][0] + xor_out[38][4][0] + xor_out[39][4][0];
assign sum_out[8][4][0] = xor_out[40][4][0] + xor_out[41][4][0] + xor_out[42][4][0] + xor_out[43][4][0] + xor_out[44][4][0];
assign sum_out[9][4][0] = xor_out[45][4][0] + xor_out[46][4][0] + xor_out[47][4][0] + xor_out[48][4][0] + xor_out[49][4][0];
assign sum_out[10][4][0] = xor_out[50][4][0] + xor_out[51][4][0] + xor_out[52][4][0] + xor_out[53][4][0] + xor_out[54][4][0];
assign sum_out[11][4][0] = xor_out[55][4][0] + xor_out[56][4][0] + xor_out[57][4][0] + xor_out[58][4][0] + xor_out[59][4][0];
assign sum_out[12][4][0] = xor_out[60][4][0] + xor_out[61][4][0] + xor_out[62][4][0] + xor_out[63][4][0] + xor_out[64][4][0];
assign sum_out[13][4][0] = xor_out[65][4][0] + xor_out[66][4][0] + xor_out[67][4][0] + xor_out[68][4][0] + xor_out[69][4][0];
assign sum_out[14][4][0] = xor_out[70][4][0] + xor_out[71][4][0] + xor_out[72][4][0] + xor_out[73][4][0] + xor_out[74][4][0];
assign sum_out[15][4][0] = xor_out[75][4][0] + xor_out[76][4][0] + xor_out[77][4][0] + xor_out[78][4][0] + xor_out[79][4][0];
assign sum_out[16][4][0] = xor_out[80][4][0] + xor_out[81][4][0] + xor_out[82][4][0] + xor_out[83][4][0] + xor_out[84][4][0];
assign sum_out[17][4][0] = xor_out[85][4][0] + xor_out[86][4][0] + xor_out[87][4][0] + xor_out[88][4][0] + xor_out[89][4][0];
assign sum_out[18][4][0] = xor_out[90][4][0] + xor_out[91][4][0] + xor_out[92][4][0] + xor_out[93][4][0] + xor_out[94][4][0];
assign sum_out[19][4][0] = xor_out[95][4][0] + xor_out[96][4][0] + xor_out[97][4][0] + xor_out[98][4][0] + xor_out[99][4][0];

assign sum_out[0][4][1] = xor_out[0][4][1] + xor_out[1][4][1] + xor_out[2][4][1] + xor_out[3][4][1] + xor_out[4][4][1];
assign sum_out[1][4][1] = xor_out[5][4][1] + xor_out[6][4][1] + xor_out[7][4][1] + xor_out[8][4][1] + xor_out[9][4][1];
assign sum_out[2][4][1] = xor_out[10][4][1] + xor_out[11][4][1] + xor_out[12][4][1] + xor_out[13][4][1] + xor_out[14][4][1];
assign sum_out[3][4][1] = xor_out[15][4][1] + xor_out[16][4][1] + xor_out[17][4][1] + xor_out[18][4][1] + xor_out[19][4][1];
assign sum_out[4][4][1] = xor_out[20][4][1] + xor_out[21][4][1] + xor_out[22][4][1] + xor_out[23][4][1] + xor_out[24][4][1];
assign sum_out[5][4][1] = xor_out[25][4][1] + xor_out[26][4][1] + xor_out[27][4][1] + xor_out[28][4][1] + xor_out[29][4][1];
assign sum_out[6][4][1] = xor_out[30][4][1] + xor_out[31][4][1] + xor_out[32][4][1] + xor_out[33][4][1] + xor_out[34][4][1];
assign sum_out[7][4][1] = xor_out[35][4][1] + xor_out[36][4][1] + xor_out[37][4][1] + xor_out[38][4][1] + xor_out[39][4][1];
assign sum_out[8][4][1] = xor_out[40][4][1] + xor_out[41][4][1] + xor_out[42][4][1] + xor_out[43][4][1] + xor_out[44][4][1];
assign sum_out[9][4][1] = xor_out[45][4][1] + xor_out[46][4][1] + xor_out[47][4][1] + xor_out[48][4][1] + xor_out[49][4][1];
assign sum_out[10][4][1] = xor_out[50][4][1] + xor_out[51][4][1] + xor_out[52][4][1] + xor_out[53][4][1] + xor_out[54][4][1];
assign sum_out[11][4][1] = xor_out[55][4][1] + xor_out[56][4][1] + xor_out[57][4][1] + xor_out[58][4][1] + xor_out[59][4][1];
assign sum_out[12][4][1] = xor_out[60][4][1] + xor_out[61][4][1] + xor_out[62][4][1] + xor_out[63][4][1] + xor_out[64][4][1];
assign sum_out[13][4][1] = xor_out[65][4][1] + xor_out[66][4][1] + xor_out[67][4][1] + xor_out[68][4][1] + xor_out[69][4][1];
assign sum_out[14][4][1] = xor_out[70][4][1] + xor_out[71][4][1] + xor_out[72][4][1] + xor_out[73][4][1] + xor_out[74][4][1];
assign sum_out[15][4][1] = xor_out[75][4][1] + xor_out[76][4][1] + xor_out[77][4][1] + xor_out[78][4][1] + xor_out[79][4][1];
assign sum_out[16][4][1] = xor_out[80][4][1] + xor_out[81][4][1] + xor_out[82][4][1] + xor_out[83][4][1] + xor_out[84][4][1];
assign sum_out[17][4][1] = xor_out[85][4][1] + xor_out[86][4][1] + xor_out[87][4][1] + xor_out[88][4][1] + xor_out[89][4][1];
assign sum_out[18][4][1] = xor_out[90][4][1] + xor_out[91][4][1] + xor_out[92][4][1] + xor_out[93][4][1] + xor_out[94][4][1];
assign sum_out[19][4][1] = xor_out[95][4][1] + xor_out[96][4][1] + xor_out[97][4][1] + xor_out[98][4][1] + xor_out[99][4][1];

assign sum_out[0][4][2] = xor_out[0][4][2] + xor_out[1][4][2] + xor_out[2][4][2] + xor_out[3][4][2] + xor_out[4][4][2];
assign sum_out[1][4][2] = xor_out[5][4][2] + xor_out[6][4][2] + xor_out[7][4][2] + xor_out[8][4][2] + xor_out[9][4][2];
assign sum_out[2][4][2] = xor_out[10][4][2] + xor_out[11][4][2] + xor_out[12][4][2] + xor_out[13][4][2] + xor_out[14][4][2];
assign sum_out[3][4][2] = xor_out[15][4][2] + xor_out[16][4][2] + xor_out[17][4][2] + xor_out[18][4][2] + xor_out[19][4][2];
assign sum_out[4][4][2] = xor_out[20][4][2] + xor_out[21][4][2] + xor_out[22][4][2] + xor_out[23][4][2] + xor_out[24][4][2];
assign sum_out[5][4][2] = xor_out[25][4][2] + xor_out[26][4][2] + xor_out[27][4][2] + xor_out[28][4][2] + xor_out[29][4][2];
assign sum_out[6][4][2] = xor_out[30][4][2] + xor_out[31][4][2] + xor_out[32][4][2] + xor_out[33][4][2] + xor_out[34][4][2];
assign sum_out[7][4][2] = xor_out[35][4][2] + xor_out[36][4][2] + xor_out[37][4][2] + xor_out[38][4][2] + xor_out[39][4][2];
assign sum_out[8][4][2] = xor_out[40][4][2] + xor_out[41][4][2] + xor_out[42][4][2] + xor_out[43][4][2] + xor_out[44][4][2];
assign sum_out[9][4][2] = xor_out[45][4][2] + xor_out[46][4][2] + xor_out[47][4][2] + xor_out[48][4][2] + xor_out[49][4][2];
assign sum_out[10][4][2] = xor_out[50][4][2] + xor_out[51][4][2] + xor_out[52][4][2] + xor_out[53][4][2] + xor_out[54][4][2];
assign sum_out[11][4][2] = xor_out[55][4][2] + xor_out[56][4][2] + xor_out[57][4][2] + xor_out[58][4][2] + xor_out[59][4][2];
assign sum_out[12][4][2] = xor_out[60][4][2] + xor_out[61][4][2] + xor_out[62][4][2] + xor_out[63][4][2] + xor_out[64][4][2];
assign sum_out[13][4][2] = xor_out[65][4][2] + xor_out[66][4][2] + xor_out[67][4][2] + xor_out[68][4][2] + xor_out[69][4][2];
assign sum_out[14][4][2] = xor_out[70][4][2] + xor_out[71][4][2] + xor_out[72][4][2] + xor_out[73][4][2] + xor_out[74][4][2];
assign sum_out[15][4][2] = xor_out[75][4][2] + xor_out[76][4][2] + xor_out[77][4][2] + xor_out[78][4][2] + xor_out[79][4][2];
assign sum_out[16][4][2] = xor_out[80][4][2] + xor_out[81][4][2] + xor_out[82][4][2] + xor_out[83][4][2] + xor_out[84][4][2];
assign sum_out[17][4][2] = xor_out[85][4][2] + xor_out[86][4][2] + xor_out[87][4][2] + xor_out[88][4][2] + xor_out[89][4][2];
assign sum_out[18][4][2] = xor_out[90][4][2] + xor_out[91][4][2] + xor_out[92][4][2] + xor_out[93][4][2] + xor_out[94][4][2];
assign sum_out[19][4][2] = xor_out[95][4][2] + xor_out[96][4][2] + xor_out[97][4][2] + xor_out[98][4][2] + xor_out[99][4][2];

assign sum_out[0][4][3] = xor_out[0][4][3] + xor_out[1][4][3] + xor_out[2][4][3] + xor_out[3][4][3] + xor_out[4][4][3];
assign sum_out[1][4][3] = xor_out[5][4][3] + xor_out[6][4][3] + xor_out[7][4][3] + xor_out[8][4][3] + xor_out[9][4][3];
assign sum_out[2][4][3] = xor_out[10][4][3] + xor_out[11][4][3] + xor_out[12][4][3] + xor_out[13][4][3] + xor_out[14][4][3];
assign sum_out[3][4][3] = xor_out[15][4][3] + xor_out[16][4][3] + xor_out[17][4][3] + xor_out[18][4][3] + xor_out[19][4][3];
assign sum_out[4][4][3] = xor_out[20][4][3] + xor_out[21][4][3] + xor_out[22][4][3] + xor_out[23][4][3] + xor_out[24][4][3];
assign sum_out[5][4][3] = xor_out[25][4][3] + xor_out[26][4][3] + xor_out[27][4][3] + xor_out[28][4][3] + xor_out[29][4][3];
assign sum_out[6][4][3] = xor_out[30][4][3] + xor_out[31][4][3] + xor_out[32][4][3] + xor_out[33][4][3] + xor_out[34][4][3];
assign sum_out[7][4][3] = xor_out[35][4][3] + xor_out[36][4][3] + xor_out[37][4][3] + xor_out[38][4][3] + xor_out[39][4][3];
assign sum_out[8][4][3] = xor_out[40][4][3] + xor_out[41][4][3] + xor_out[42][4][3] + xor_out[43][4][3] + xor_out[44][4][3];
assign sum_out[9][4][3] = xor_out[45][4][3] + xor_out[46][4][3] + xor_out[47][4][3] + xor_out[48][4][3] + xor_out[49][4][3];
assign sum_out[10][4][3] = xor_out[50][4][3] + xor_out[51][4][3] + xor_out[52][4][3] + xor_out[53][4][3] + xor_out[54][4][3];
assign sum_out[11][4][3] = xor_out[55][4][3] + xor_out[56][4][3] + xor_out[57][4][3] + xor_out[58][4][3] + xor_out[59][4][3];
assign sum_out[12][4][3] = xor_out[60][4][3] + xor_out[61][4][3] + xor_out[62][4][3] + xor_out[63][4][3] + xor_out[64][4][3];
assign sum_out[13][4][3] = xor_out[65][4][3] + xor_out[66][4][3] + xor_out[67][4][3] + xor_out[68][4][3] + xor_out[69][4][3];
assign sum_out[14][4][3] = xor_out[70][4][3] + xor_out[71][4][3] + xor_out[72][4][3] + xor_out[73][4][3] + xor_out[74][4][3];
assign sum_out[15][4][3] = xor_out[75][4][3] + xor_out[76][4][3] + xor_out[77][4][3] + xor_out[78][4][3] + xor_out[79][4][3];
assign sum_out[16][4][3] = xor_out[80][4][3] + xor_out[81][4][3] + xor_out[82][4][3] + xor_out[83][4][3] + xor_out[84][4][3];
assign sum_out[17][4][3] = xor_out[85][4][3] + xor_out[86][4][3] + xor_out[87][4][3] + xor_out[88][4][3] + xor_out[89][4][3];
assign sum_out[18][4][3] = xor_out[90][4][3] + xor_out[91][4][3] + xor_out[92][4][3] + xor_out[93][4][3] + xor_out[94][4][3];
assign sum_out[19][4][3] = xor_out[95][4][3] + xor_out[96][4][3] + xor_out[97][4][3] + xor_out[98][4][3] + xor_out[99][4][3];

assign sum_out[0][4][4] = xor_out[0][4][4] + xor_out[1][4][4] + xor_out[2][4][4] + xor_out[3][4][4] + xor_out[4][4][4];
assign sum_out[1][4][4] = xor_out[5][4][4] + xor_out[6][4][4] + xor_out[7][4][4] + xor_out[8][4][4] + xor_out[9][4][4];
assign sum_out[2][4][4] = xor_out[10][4][4] + xor_out[11][4][4] + xor_out[12][4][4] + xor_out[13][4][4] + xor_out[14][4][4];
assign sum_out[3][4][4] = xor_out[15][4][4] + xor_out[16][4][4] + xor_out[17][4][4] + xor_out[18][4][4] + xor_out[19][4][4];
assign sum_out[4][4][4] = xor_out[20][4][4] + xor_out[21][4][4] + xor_out[22][4][4] + xor_out[23][4][4] + xor_out[24][4][4];
assign sum_out[5][4][4] = xor_out[25][4][4] + xor_out[26][4][4] + xor_out[27][4][4] + xor_out[28][4][4] + xor_out[29][4][4];
assign sum_out[6][4][4] = xor_out[30][4][4] + xor_out[31][4][4] + xor_out[32][4][4] + xor_out[33][4][4] + xor_out[34][4][4];
assign sum_out[7][4][4] = xor_out[35][4][4] + xor_out[36][4][4] + xor_out[37][4][4] + xor_out[38][4][4] + xor_out[39][4][4];
assign sum_out[8][4][4] = xor_out[40][4][4] + xor_out[41][4][4] + xor_out[42][4][4] + xor_out[43][4][4] + xor_out[44][4][4];
assign sum_out[9][4][4] = xor_out[45][4][4] + xor_out[46][4][4] + xor_out[47][4][4] + xor_out[48][4][4] + xor_out[49][4][4];
assign sum_out[10][4][4] = xor_out[50][4][4] + xor_out[51][4][4] + xor_out[52][4][4] + xor_out[53][4][4] + xor_out[54][4][4];
assign sum_out[11][4][4] = xor_out[55][4][4] + xor_out[56][4][4] + xor_out[57][4][4] + xor_out[58][4][4] + xor_out[59][4][4];
assign sum_out[12][4][4] = xor_out[60][4][4] + xor_out[61][4][4] + xor_out[62][4][4] + xor_out[63][4][4] + xor_out[64][4][4];
assign sum_out[13][4][4] = xor_out[65][4][4] + xor_out[66][4][4] + xor_out[67][4][4] + xor_out[68][4][4] + xor_out[69][4][4];
assign sum_out[14][4][4] = xor_out[70][4][4] + xor_out[71][4][4] + xor_out[72][4][4] + xor_out[73][4][4] + xor_out[74][4][4];
assign sum_out[15][4][4] = xor_out[75][4][4] + xor_out[76][4][4] + xor_out[77][4][4] + xor_out[78][4][4] + xor_out[79][4][4];
assign sum_out[16][4][4] = xor_out[80][4][4] + xor_out[81][4][4] + xor_out[82][4][4] + xor_out[83][4][4] + xor_out[84][4][4];
assign sum_out[17][4][4] = xor_out[85][4][4] + xor_out[86][4][4] + xor_out[87][4][4] + xor_out[88][4][4] + xor_out[89][4][4];
assign sum_out[18][4][4] = xor_out[90][4][4] + xor_out[91][4][4] + xor_out[92][4][4] + xor_out[93][4][4] + xor_out[94][4][4];
assign sum_out[19][4][4] = xor_out[95][4][4] + xor_out[96][4][4] + xor_out[97][4][4] + xor_out[98][4][4] + xor_out[99][4][4];

assign sum_out[0][4][5] = xor_out[0][4][5] + xor_out[1][4][5] + xor_out[2][4][5] + xor_out[3][4][5] + xor_out[4][4][5];
assign sum_out[1][4][5] = xor_out[5][4][5] + xor_out[6][4][5] + xor_out[7][4][5] + xor_out[8][4][5] + xor_out[9][4][5];
assign sum_out[2][4][5] = xor_out[10][4][5] + xor_out[11][4][5] + xor_out[12][4][5] + xor_out[13][4][5] + xor_out[14][4][5];
assign sum_out[3][4][5] = xor_out[15][4][5] + xor_out[16][4][5] + xor_out[17][4][5] + xor_out[18][4][5] + xor_out[19][4][5];
assign sum_out[4][4][5] = xor_out[20][4][5] + xor_out[21][4][5] + xor_out[22][4][5] + xor_out[23][4][5] + xor_out[24][4][5];
assign sum_out[5][4][5] = xor_out[25][4][5] + xor_out[26][4][5] + xor_out[27][4][5] + xor_out[28][4][5] + xor_out[29][4][5];
assign sum_out[6][4][5] = xor_out[30][4][5] + xor_out[31][4][5] + xor_out[32][4][5] + xor_out[33][4][5] + xor_out[34][4][5];
assign sum_out[7][4][5] = xor_out[35][4][5] + xor_out[36][4][5] + xor_out[37][4][5] + xor_out[38][4][5] + xor_out[39][4][5];
assign sum_out[8][4][5] = xor_out[40][4][5] + xor_out[41][4][5] + xor_out[42][4][5] + xor_out[43][4][5] + xor_out[44][4][5];
assign sum_out[9][4][5] = xor_out[45][4][5] + xor_out[46][4][5] + xor_out[47][4][5] + xor_out[48][4][5] + xor_out[49][4][5];
assign sum_out[10][4][5] = xor_out[50][4][5] + xor_out[51][4][5] + xor_out[52][4][5] + xor_out[53][4][5] + xor_out[54][4][5];
assign sum_out[11][4][5] = xor_out[55][4][5] + xor_out[56][4][5] + xor_out[57][4][5] + xor_out[58][4][5] + xor_out[59][4][5];
assign sum_out[12][4][5] = xor_out[60][4][5] + xor_out[61][4][5] + xor_out[62][4][5] + xor_out[63][4][5] + xor_out[64][4][5];
assign sum_out[13][4][5] = xor_out[65][4][5] + xor_out[66][4][5] + xor_out[67][4][5] + xor_out[68][4][5] + xor_out[69][4][5];
assign sum_out[14][4][5] = xor_out[70][4][5] + xor_out[71][4][5] + xor_out[72][4][5] + xor_out[73][4][5] + xor_out[74][4][5];
assign sum_out[15][4][5] = xor_out[75][4][5] + xor_out[76][4][5] + xor_out[77][4][5] + xor_out[78][4][5] + xor_out[79][4][5];
assign sum_out[16][4][5] = xor_out[80][4][5] + xor_out[81][4][5] + xor_out[82][4][5] + xor_out[83][4][5] + xor_out[84][4][5];
assign sum_out[17][4][5] = xor_out[85][4][5] + xor_out[86][4][5] + xor_out[87][4][5] + xor_out[88][4][5] + xor_out[89][4][5];
assign sum_out[18][4][5] = xor_out[90][4][5] + xor_out[91][4][5] + xor_out[92][4][5] + xor_out[93][4][5] + xor_out[94][4][5];
assign sum_out[19][4][5] = xor_out[95][4][5] + xor_out[96][4][5] + xor_out[97][4][5] + xor_out[98][4][5] + xor_out[99][4][5];

assign sum_out[0][4][6] = xor_out[0][4][6] + xor_out[1][4][6] + xor_out[2][4][6] + xor_out[3][4][6] + xor_out[4][4][6];
assign sum_out[1][4][6] = xor_out[5][4][6] + xor_out[6][4][6] + xor_out[7][4][6] + xor_out[8][4][6] + xor_out[9][4][6];
assign sum_out[2][4][6] = xor_out[10][4][6] + xor_out[11][4][6] + xor_out[12][4][6] + xor_out[13][4][6] + xor_out[14][4][6];
assign sum_out[3][4][6] = xor_out[15][4][6] + xor_out[16][4][6] + xor_out[17][4][6] + xor_out[18][4][6] + xor_out[19][4][6];
assign sum_out[4][4][6] = xor_out[20][4][6] + xor_out[21][4][6] + xor_out[22][4][6] + xor_out[23][4][6] + xor_out[24][4][6];
assign sum_out[5][4][6] = xor_out[25][4][6] + xor_out[26][4][6] + xor_out[27][4][6] + xor_out[28][4][6] + xor_out[29][4][6];
assign sum_out[6][4][6] = xor_out[30][4][6] + xor_out[31][4][6] + xor_out[32][4][6] + xor_out[33][4][6] + xor_out[34][4][6];
assign sum_out[7][4][6] = xor_out[35][4][6] + xor_out[36][4][6] + xor_out[37][4][6] + xor_out[38][4][6] + xor_out[39][4][6];
assign sum_out[8][4][6] = xor_out[40][4][6] + xor_out[41][4][6] + xor_out[42][4][6] + xor_out[43][4][6] + xor_out[44][4][6];
assign sum_out[9][4][6] = xor_out[45][4][6] + xor_out[46][4][6] + xor_out[47][4][6] + xor_out[48][4][6] + xor_out[49][4][6];
assign sum_out[10][4][6] = xor_out[50][4][6] + xor_out[51][4][6] + xor_out[52][4][6] + xor_out[53][4][6] + xor_out[54][4][6];
assign sum_out[11][4][6] = xor_out[55][4][6] + xor_out[56][4][6] + xor_out[57][4][6] + xor_out[58][4][6] + xor_out[59][4][6];
assign sum_out[12][4][6] = xor_out[60][4][6] + xor_out[61][4][6] + xor_out[62][4][6] + xor_out[63][4][6] + xor_out[64][4][6];
assign sum_out[13][4][6] = xor_out[65][4][6] + xor_out[66][4][6] + xor_out[67][4][6] + xor_out[68][4][6] + xor_out[69][4][6];
assign sum_out[14][4][6] = xor_out[70][4][6] + xor_out[71][4][6] + xor_out[72][4][6] + xor_out[73][4][6] + xor_out[74][4][6];
assign sum_out[15][4][6] = xor_out[75][4][6] + xor_out[76][4][6] + xor_out[77][4][6] + xor_out[78][4][6] + xor_out[79][4][6];
assign sum_out[16][4][6] = xor_out[80][4][6] + xor_out[81][4][6] + xor_out[82][4][6] + xor_out[83][4][6] + xor_out[84][4][6];
assign sum_out[17][4][6] = xor_out[85][4][6] + xor_out[86][4][6] + xor_out[87][4][6] + xor_out[88][4][6] + xor_out[89][4][6];
assign sum_out[18][4][6] = xor_out[90][4][6] + xor_out[91][4][6] + xor_out[92][4][6] + xor_out[93][4][6] + xor_out[94][4][6];
assign sum_out[19][4][6] = xor_out[95][4][6] + xor_out[96][4][6] + xor_out[97][4][6] + xor_out[98][4][6] + xor_out[99][4][6];

assign sum_out[0][4][7] = xor_out[0][4][7] + xor_out[1][4][7] + xor_out[2][4][7] + xor_out[3][4][7] + xor_out[4][4][7];
assign sum_out[1][4][7] = xor_out[5][4][7] + xor_out[6][4][7] + xor_out[7][4][7] + xor_out[8][4][7] + xor_out[9][4][7];
assign sum_out[2][4][7] = xor_out[10][4][7] + xor_out[11][4][7] + xor_out[12][4][7] + xor_out[13][4][7] + xor_out[14][4][7];
assign sum_out[3][4][7] = xor_out[15][4][7] + xor_out[16][4][7] + xor_out[17][4][7] + xor_out[18][4][7] + xor_out[19][4][7];
assign sum_out[4][4][7] = xor_out[20][4][7] + xor_out[21][4][7] + xor_out[22][4][7] + xor_out[23][4][7] + xor_out[24][4][7];
assign sum_out[5][4][7] = xor_out[25][4][7] + xor_out[26][4][7] + xor_out[27][4][7] + xor_out[28][4][7] + xor_out[29][4][7];
assign sum_out[6][4][7] = xor_out[30][4][7] + xor_out[31][4][7] + xor_out[32][4][7] + xor_out[33][4][7] + xor_out[34][4][7];
assign sum_out[7][4][7] = xor_out[35][4][7] + xor_out[36][4][7] + xor_out[37][4][7] + xor_out[38][4][7] + xor_out[39][4][7];
assign sum_out[8][4][7] = xor_out[40][4][7] + xor_out[41][4][7] + xor_out[42][4][7] + xor_out[43][4][7] + xor_out[44][4][7];
assign sum_out[9][4][7] = xor_out[45][4][7] + xor_out[46][4][7] + xor_out[47][4][7] + xor_out[48][4][7] + xor_out[49][4][7];
assign sum_out[10][4][7] = xor_out[50][4][7] + xor_out[51][4][7] + xor_out[52][4][7] + xor_out[53][4][7] + xor_out[54][4][7];
assign sum_out[11][4][7] = xor_out[55][4][7] + xor_out[56][4][7] + xor_out[57][4][7] + xor_out[58][4][7] + xor_out[59][4][7];
assign sum_out[12][4][7] = xor_out[60][4][7] + xor_out[61][4][7] + xor_out[62][4][7] + xor_out[63][4][7] + xor_out[64][4][7];
assign sum_out[13][4][7] = xor_out[65][4][7] + xor_out[66][4][7] + xor_out[67][4][7] + xor_out[68][4][7] + xor_out[69][4][7];
assign sum_out[14][4][7] = xor_out[70][4][7] + xor_out[71][4][7] + xor_out[72][4][7] + xor_out[73][4][7] + xor_out[74][4][7];
assign sum_out[15][4][7] = xor_out[75][4][7] + xor_out[76][4][7] + xor_out[77][4][7] + xor_out[78][4][7] + xor_out[79][4][7];
assign sum_out[16][4][7] = xor_out[80][4][7] + xor_out[81][4][7] + xor_out[82][4][7] + xor_out[83][4][7] + xor_out[84][4][7];
assign sum_out[17][4][7] = xor_out[85][4][7] + xor_out[86][4][7] + xor_out[87][4][7] + xor_out[88][4][7] + xor_out[89][4][7];
assign sum_out[18][4][7] = xor_out[90][4][7] + xor_out[91][4][7] + xor_out[92][4][7] + xor_out[93][4][7] + xor_out[94][4][7];
assign sum_out[19][4][7] = xor_out[95][4][7] + xor_out[96][4][7] + xor_out[97][4][7] + xor_out[98][4][7] + xor_out[99][4][7];

assign sum_out[0][4][8] = xor_out[0][4][8] + xor_out[1][4][8] + xor_out[2][4][8] + xor_out[3][4][8] + xor_out[4][4][8];
assign sum_out[1][4][8] = xor_out[5][4][8] + xor_out[6][4][8] + xor_out[7][4][8] + xor_out[8][4][8] + xor_out[9][4][8];
assign sum_out[2][4][8] = xor_out[10][4][8] + xor_out[11][4][8] + xor_out[12][4][8] + xor_out[13][4][8] + xor_out[14][4][8];
assign sum_out[3][4][8] = xor_out[15][4][8] + xor_out[16][4][8] + xor_out[17][4][8] + xor_out[18][4][8] + xor_out[19][4][8];
assign sum_out[4][4][8] = xor_out[20][4][8] + xor_out[21][4][8] + xor_out[22][4][8] + xor_out[23][4][8] + xor_out[24][4][8];
assign sum_out[5][4][8] = xor_out[25][4][8] + xor_out[26][4][8] + xor_out[27][4][8] + xor_out[28][4][8] + xor_out[29][4][8];
assign sum_out[6][4][8] = xor_out[30][4][8] + xor_out[31][4][8] + xor_out[32][4][8] + xor_out[33][4][8] + xor_out[34][4][8];
assign sum_out[7][4][8] = xor_out[35][4][8] + xor_out[36][4][8] + xor_out[37][4][8] + xor_out[38][4][8] + xor_out[39][4][8];
assign sum_out[8][4][8] = xor_out[40][4][8] + xor_out[41][4][8] + xor_out[42][4][8] + xor_out[43][4][8] + xor_out[44][4][8];
assign sum_out[9][4][8] = xor_out[45][4][8] + xor_out[46][4][8] + xor_out[47][4][8] + xor_out[48][4][8] + xor_out[49][4][8];
assign sum_out[10][4][8] = xor_out[50][4][8] + xor_out[51][4][8] + xor_out[52][4][8] + xor_out[53][4][8] + xor_out[54][4][8];
assign sum_out[11][4][8] = xor_out[55][4][8] + xor_out[56][4][8] + xor_out[57][4][8] + xor_out[58][4][8] + xor_out[59][4][8];
assign sum_out[12][4][8] = xor_out[60][4][8] + xor_out[61][4][8] + xor_out[62][4][8] + xor_out[63][4][8] + xor_out[64][4][8];
assign sum_out[13][4][8] = xor_out[65][4][8] + xor_out[66][4][8] + xor_out[67][4][8] + xor_out[68][4][8] + xor_out[69][4][8];
assign sum_out[14][4][8] = xor_out[70][4][8] + xor_out[71][4][8] + xor_out[72][4][8] + xor_out[73][4][8] + xor_out[74][4][8];
assign sum_out[15][4][8] = xor_out[75][4][8] + xor_out[76][4][8] + xor_out[77][4][8] + xor_out[78][4][8] + xor_out[79][4][8];
assign sum_out[16][4][8] = xor_out[80][4][8] + xor_out[81][4][8] + xor_out[82][4][8] + xor_out[83][4][8] + xor_out[84][4][8];
assign sum_out[17][4][8] = xor_out[85][4][8] + xor_out[86][4][8] + xor_out[87][4][8] + xor_out[88][4][8] + xor_out[89][4][8];
assign sum_out[18][4][8] = xor_out[90][4][8] + xor_out[91][4][8] + xor_out[92][4][8] + xor_out[93][4][8] + xor_out[94][4][8];
assign sum_out[19][4][8] = xor_out[95][4][8] + xor_out[96][4][8] + xor_out[97][4][8] + xor_out[98][4][8] + xor_out[99][4][8];

assign sum_out[0][4][9] = xor_out[0][4][9] + xor_out[1][4][9] + xor_out[2][4][9] + xor_out[3][4][9] + xor_out[4][4][9];
assign sum_out[1][4][9] = xor_out[5][4][9] + xor_out[6][4][9] + xor_out[7][4][9] + xor_out[8][4][9] + xor_out[9][4][9];
assign sum_out[2][4][9] = xor_out[10][4][9] + xor_out[11][4][9] + xor_out[12][4][9] + xor_out[13][4][9] + xor_out[14][4][9];
assign sum_out[3][4][9] = xor_out[15][4][9] + xor_out[16][4][9] + xor_out[17][4][9] + xor_out[18][4][9] + xor_out[19][4][9];
assign sum_out[4][4][9] = xor_out[20][4][9] + xor_out[21][4][9] + xor_out[22][4][9] + xor_out[23][4][9] + xor_out[24][4][9];
assign sum_out[5][4][9] = xor_out[25][4][9] + xor_out[26][4][9] + xor_out[27][4][9] + xor_out[28][4][9] + xor_out[29][4][9];
assign sum_out[6][4][9] = xor_out[30][4][9] + xor_out[31][4][9] + xor_out[32][4][9] + xor_out[33][4][9] + xor_out[34][4][9];
assign sum_out[7][4][9] = xor_out[35][4][9] + xor_out[36][4][9] + xor_out[37][4][9] + xor_out[38][4][9] + xor_out[39][4][9];
assign sum_out[8][4][9] = xor_out[40][4][9] + xor_out[41][4][9] + xor_out[42][4][9] + xor_out[43][4][9] + xor_out[44][4][9];
assign sum_out[9][4][9] = xor_out[45][4][9] + xor_out[46][4][9] + xor_out[47][4][9] + xor_out[48][4][9] + xor_out[49][4][9];
assign sum_out[10][4][9] = xor_out[50][4][9] + xor_out[51][4][9] + xor_out[52][4][9] + xor_out[53][4][9] + xor_out[54][4][9];
assign sum_out[11][4][9] = xor_out[55][4][9] + xor_out[56][4][9] + xor_out[57][4][9] + xor_out[58][4][9] + xor_out[59][4][9];
assign sum_out[12][4][9] = xor_out[60][4][9] + xor_out[61][4][9] + xor_out[62][4][9] + xor_out[63][4][9] + xor_out[64][4][9];
assign sum_out[13][4][9] = xor_out[65][4][9] + xor_out[66][4][9] + xor_out[67][4][9] + xor_out[68][4][9] + xor_out[69][4][9];
assign sum_out[14][4][9] = xor_out[70][4][9] + xor_out[71][4][9] + xor_out[72][4][9] + xor_out[73][4][9] + xor_out[74][4][9];
assign sum_out[15][4][9] = xor_out[75][4][9] + xor_out[76][4][9] + xor_out[77][4][9] + xor_out[78][4][9] + xor_out[79][4][9];
assign sum_out[16][4][9] = xor_out[80][4][9] + xor_out[81][4][9] + xor_out[82][4][9] + xor_out[83][4][9] + xor_out[84][4][9];
assign sum_out[17][4][9] = xor_out[85][4][9] + xor_out[86][4][9] + xor_out[87][4][9] + xor_out[88][4][9] + xor_out[89][4][9];
assign sum_out[18][4][9] = xor_out[90][4][9] + xor_out[91][4][9] + xor_out[92][4][9] + xor_out[93][4][9] + xor_out[94][4][9];
assign sum_out[19][4][9] = xor_out[95][4][9] + xor_out[96][4][9] + xor_out[97][4][9] + xor_out[98][4][9] + xor_out[99][4][9];

assign sum_out[0][4][10] = xor_out[0][4][10] + xor_out[1][4][10] + xor_out[2][4][10] + xor_out[3][4][10] + xor_out[4][4][10];
assign sum_out[1][4][10] = xor_out[5][4][10] + xor_out[6][4][10] + xor_out[7][4][10] + xor_out[8][4][10] + xor_out[9][4][10];
assign sum_out[2][4][10] = xor_out[10][4][10] + xor_out[11][4][10] + xor_out[12][4][10] + xor_out[13][4][10] + xor_out[14][4][10];
assign sum_out[3][4][10] = xor_out[15][4][10] + xor_out[16][4][10] + xor_out[17][4][10] + xor_out[18][4][10] + xor_out[19][4][10];
assign sum_out[4][4][10] = xor_out[20][4][10] + xor_out[21][4][10] + xor_out[22][4][10] + xor_out[23][4][10] + xor_out[24][4][10];
assign sum_out[5][4][10] = xor_out[25][4][10] + xor_out[26][4][10] + xor_out[27][4][10] + xor_out[28][4][10] + xor_out[29][4][10];
assign sum_out[6][4][10] = xor_out[30][4][10] + xor_out[31][4][10] + xor_out[32][4][10] + xor_out[33][4][10] + xor_out[34][4][10];
assign sum_out[7][4][10] = xor_out[35][4][10] + xor_out[36][4][10] + xor_out[37][4][10] + xor_out[38][4][10] + xor_out[39][4][10];
assign sum_out[8][4][10] = xor_out[40][4][10] + xor_out[41][4][10] + xor_out[42][4][10] + xor_out[43][4][10] + xor_out[44][4][10];
assign sum_out[9][4][10] = xor_out[45][4][10] + xor_out[46][4][10] + xor_out[47][4][10] + xor_out[48][4][10] + xor_out[49][4][10];
assign sum_out[10][4][10] = xor_out[50][4][10] + xor_out[51][4][10] + xor_out[52][4][10] + xor_out[53][4][10] + xor_out[54][4][10];
assign sum_out[11][4][10] = xor_out[55][4][10] + xor_out[56][4][10] + xor_out[57][4][10] + xor_out[58][4][10] + xor_out[59][4][10];
assign sum_out[12][4][10] = xor_out[60][4][10] + xor_out[61][4][10] + xor_out[62][4][10] + xor_out[63][4][10] + xor_out[64][4][10];
assign sum_out[13][4][10] = xor_out[65][4][10] + xor_out[66][4][10] + xor_out[67][4][10] + xor_out[68][4][10] + xor_out[69][4][10];
assign sum_out[14][4][10] = xor_out[70][4][10] + xor_out[71][4][10] + xor_out[72][4][10] + xor_out[73][4][10] + xor_out[74][4][10];
assign sum_out[15][4][10] = xor_out[75][4][10] + xor_out[76][4][10] + xor_out[77][4][10] + xor_out[78][4][10] + xor_out[79][4][10];
assign sum_out[16][4][10] = xor_out[80][4][10] + xor_out[81][4][10] + xor_out[82][4][10] + xor_out[83][4][10] + xor_out[84][4][10];
assign sum_out[17][4][10] = xor_out[85][4][10] + xor_out[86][4][10] + xor_out[87][4][10] + xor_out[88][4][10] + xor_out[89][4][10];
assign sum_out[18][4][10] = xor_out[90][4][10] + xor_out[91][4][10] + xor_out[92][4][10] + xor_out[93][4][10] + xor_out[94][4][10];
assign sum_out[19][4][10] = xor_out[95][4][10] + xor_out[96][4][10] + xor_out[97][4][10] + xor_out[98][4][10] + xor_out[99][4][10];

assign sum_out[0][4][11] = xor_out[0][4][11] + xor_out[1][4][11] + xor_out[2][4][11] + xor_out[3][4][11] + xor_out[4][4][11];
assign sum_out[1][4][11] = xor_out[5][4][11] + xor_out[6][4][11] + xor_out[7][4][11] + xor_out[8][4][11] + xor_out[9][4][11];
assign sum_out[2][4][11] = xor_out[10][4][11] + xor_out[11][4][11] + xor_out[12][4][11] + xor_out[13][4][11] + xor_out[14][4][11];
assign sum_out[3][4][11] = xor_out[15][4][11] + xor_out[16][4][11] + xor_out[17][4][11] + xor_out[18][4][11] + xor_out[19][4][11];
assign sum_out[4][4][11] = xor_out[20][4][11] + xor_out[21][4][11] + xor_out[22][4][11] + xor_out[23][4][11] + xor_out[24][4][11];
assign sum_out[5][4][11] = xor_out[25][4][11] + xor_out[26][4][11] + xor_out[27][4][11] + xor_out[28][4][11] + xor_out[29][4][11];
assign sum_out[6][4][11] = xor_out[30][4][11] + xor_out[31][4][11] + xor_out[32][4][11] + xor_out[33][4][11] + xor_out[34][4][11];
assign sum_out[7][4][11] = xor_out[35][4][11] + xor_out[36][4][11] + xor_out[37][4][11] + xor_out[38][4][11] + xor_out[39][4][11];
assign sum_out[8][4][11] = xor_out[40][4][11] + xor_out[41][4][11] + xor_out[42][4][11] + xor_out[43][4][11] + xor_out[44][4][11];
assign sum_out[9][4][11] = xor_out[45][4][11] + xor_out[46][4][11] + xor_out[47][4][11] + xor_out[48][4][11] + xor_out[49][4][11];
assign sum_out[10][4][11] = xor_out[50][4][11] + xor_out[51][4][11] + xor_out[52][4][11] + xor_out[53][4][11] + xor_out[54][4][11];
assign sum_out[11][4][11] = xor_out[55][4][11] + xor_out[56][4][11] + xor_out[57][4][11] + xor_out[58][4][11] + xor_out[59][4][11];
assign sum_out[12][4][11] = xor_out[60][4][11] + xor_out[61][4][11] + xor_out[62][4][11] + xor_out[63][4][11] + xor_out[64][4][11];
assign sum_out[13][4][11] = xor_out[65][4][11] + xor_out[66][4][11] + xor_out[67][4][11] + xor_out[68][4][11] + xor_out[69][4][11];
assign sum_out[14][4][11] = xor_out[70][4][11] + xor_out[71][4][11] + xor_out[72][4][11] + xor_out[73][4][11] + xor_out[74][4][11];
assign sum_out[15][4][11] = xor_out[75][4][11] + xor_out[76][4][11] + xor_out[77][4][11] + xor_out[78][4][11] + xor_out[79][4][11];
assign sum_out[16][4][11] = xor_out[80][4][11] + xor_out[81][4][11] + xor_out[82][4][11] + xor_out[83][4][11] + xor_out[84][4][11];
assign sum_out[17][4][11] = xor_out[85][4][11] + xor_out[86][4][11] + xor_out[87][4][11] + xor_out[88][4][11] + xor_out[89][4][11];
assign sum_out[18][4][11] = xor_out[90][4][11] + xor_out[91][4][11] + xor_out[92][4][11] + xor_out[93][4][11] + xor_out[94][4][11];
assign sum_out[19][4][11] = xor_out[95][4][11] + xor_out[96][4][11] + xor_out[97][4][11] + xor_out[98][4][11] + xor_out[99][4][11];

assign sum_out[0][4][12] = xor_out[0][4][12] + xor_out[1][4][12] + xor_out[2][4][12] + xor_out[3][4][12] + xor_out[4][4][12];
assign sum_out[1][4][12] = xor_out[5][4][12] + xor_out[6][4][12] + xor_out[7][4][12] + xor_out[8][4][12] + xor_out[9][4][12];
assign sum_out[2][4][12] = xor_out[10][4][12] + xor_out[11][4][12] + xor_out[12][4][12] + xor_out[13][4][12] + xor_out[14][4][12];
assign sum_out[3][4][12] = xor_out[15][4][12] + xor_out[16][4][12] + xor_out[17][4][12] + xor_out[18][4][12] + xor_out[19][4][12];
assign sum_out[4][4][12] = xor_out[20][4][12] + xor_out[21][4][12] + xor_out[22][4][12] + xor_out[23][4][12] + xor_out[24][4][12];
assign sum_out[5][4][12] = xor_out[25][4][12] + xor_out[26][4][12] + xor_out[27][4][12] + xor_out[28][4][12] + xor_out[29][4][12];
assign sum_out[6][4][12] = xor_out[30][4][12] + xor_out[31][4][12] + xor_out[32][4][12] + xor_out[33][4][12] + xor_out[34][4][12];
assign sum_out[7][4][12] = xor_out[35][4][12] + xor_out[36][4][12] + xor_out[37][4][12] + xor_out[38][4][12] + xor_out[39][4][12];
assign sum_out[8][4][12] = xor_out[40][4][12] + xor_out[41][4][12] + xor_out[42][4][12] + xor_out[43][4][12] + xor_out[44][4][12];
assign sum_out[9][4][12] = xor_out[45][4][12] + xor_out[46][4][12] + xor_out[47][4][12] + xor_out[48][4][12] + xor_out[49][4][12];
assign sum_out[10][4][12] = xor_out[50][4][12] + xor_out[51][4][12] + xor_out[52][4][12] + xor_out[53][4][12] + xor_out[54][4][12];
assign sum_out[11][4][12] = xor_out[55][4][12] + xor_out[56][4][12] + xor_out[57][4][12] + xor_out[58][4][12] + xor_out[59][4][12];
assign sum_out[12][4][12] = xor_out[60][4][12] + xor_out[61][4][12] + xor_out[62][4][12] + xor_out[63][4][12] + xor_out[64][4][12];
assign sum_out[13][4][12] = xor_out[65][4][12] + xor_out[66][4][12] + xor_out[67][4][12] + xor_out[68][4][12] + xor_out[69][4][12];
assign sum_out[14][4][12] = xor_out[70][4][12] + xor_out[71][4][12] + xor_out[72][4][12] + xor_out[73][4][12] + xor_out[74][4][12];
assign sum_out[15][4][12] = xor_out[75][4][12] + xor_out[76][4][12] + xor_out[77][4][12] + xor_out[78][4][12] + xor_out[79][4][12];
assign sum_out[16][4][12] = xor_out[80][4][12] + xor_out[81][4][12] + xor_out[82][4][12] + xor_out[83][4][12] + xor_out[84][4][12];
assign sum_out[17][4][12] = xor_out[85][4][12] + xor_out[86][4][12] + xor_out[87][4][12] + xor_out[88][4][12] + xor_out[89][4][12];
assign sum_out[18][4][12] = xor_out[90][4][12] + xor_out[91][4][12] + xor_out[92][4][12] + xor_out[93][4][12] + xor_out[94][4][12];
assign sum_out[19][4][12] = xor_out[95][4][12] + xor_out[96][4][12] + xor_out[97][4][12] + xor_out[98][4][12] + xor_out[99][4][12];

assign sum_out[0][4][13] = xor_out[0][4][13] + xor_out[1][4][13] + xor_out[2][4][13] + xor_out[3][4][13] + xor_out[4][4][13];
assign sum_out[1][4][13] = xor_out[5][4][13] + xor_out[6][4][13] + xor_out[7][4][13] + xor_out[8][4][13] + xor_out[9][4][13];
assign sum_out[2][4][13] = xor_out[10][4][13] + xor_out[11][4][13] + xor_out[12][4][13] + xor_out[13][4][13] + xor_out[14][4][13];
assign sum_out[3][4][13] = xor_out[15][4][13] + xor_out[16][4][13] + xor_out[17][4][13] + xor_out[18][4][13] + xor_out[19][4][13];
assign sum_out[4][4][13] = xor_out[20][4][13] + xor_out[21][4][13] + xor_out[22][4][13] + xor_out[23][4][13] + xor_out[24][4][13];
assign sum_out[5][4][13] = xor_out[25][4][13] + xor_out[26][4][13] + xor_out[27][4][13] + xor_out[28][4][13] + xor_out[29][4][13];
assign sum_out[6][4][13] = xor_out[30][4][13] + xor_out[31][4][13] + xor_out[32][4][13] + xor_out[33][4][13] + xor_out[34][4][13];
assign sum_out[7][4][13] = xor_out[35][4][13] + xor_out[36][4][13] + xor_out[37][4][13] + xor_out[38][4][13] + xor_out[39][4][13];
assign sum_out[8][4][13] = xor_out[40][4][13] + xor_out[41][4][13] + xor_out[42][4][13] + xor_out[43][4][13] + xor_out[44][4][13];
assign sum_out[9][4][13] = xor_out[45][4][13] + xor_out[46][4][13] + xor_out[47][4][13] + xor_out[48][4][13] + xor_out[49][4][13];
assign sum_out[10][4][13] = xor_out[50][4][13] + xor_out[51][4][13] + xor_out[52][4][13] + xor_out[53][4][13] + xor_out[54][4][13];
assign sum_out[11][4][13] = xor_out[55][4][13] + xor_out[56][4][13] + xor_out[57][4][13] + xor_out[58][4][13] + xor_out[59][4][13];
assign sum_out[12][4][13] = xor_out[60][4][13] + xor_out[61][4][13] + xor_out[62][4][13] + xor_out[63][4][13] + xor_out[64][4][13];
assign sum_out[13][4][13] = xor_out[65][4][13] + xor_out[66][4][13] + xor_out[67][4][13] + xor_out[68][4][13] + xor_out[69][4][13];
assign sum_out[14][4][13] = xor_out[70][4][13] + xor_out[71][4][13] + xor_out[72][4][13] + xor_out[73][4][13] + xor_out[74][4][13];
assign sum_out[15][4][13] = xor_out[75][4][13] + xor_out[76][4][13] + xor_out[77][4][13] + xor_out[78][4][13] + xor_out[79][4][13];
assign sum_out[16][4][13] = xor_out[80][4][13] + xor_out[81][4][13] + xor_out[82][4][13] + xor_out[83][4][13] + xor_out[84][4][13];
assign sum_out[17][4][13] = xor_out[85][4][13] + xor_out[86][4][13] + xor_out[87][4][13] + xor_out[88][4][13] + xor_out[89][4][13];
assign sum_out[18][4][13] = xor_out[90][4][13] + xor_out[91][4][13] + xor_out[92][4][13] + xor_out[93][4][13] + xor_out[94][4][13];
assign sum_out[19][4][13] = xor_out[95][4][13] + xor_out[96][4][13] + xor_out[97][4][13] + xor_out[98][4][13] + xor_out[99][4][13];

assign sum_out[0][4][14] = xor_out[0][4][14] + xor_out[1][4][14] + xor_out[2][4][14] + xor_out[3][4][14] + xor_out[4][4][14];
assign sum_out[1][4][14] = xor_out[5][4][14] + xor_out[6][4][14] + xor_out[7][4][14] + xor_out[8][4][14] + xor_out[9][4][14];
assign sum_out[2][4][14] = xor_out[10][4][14] + xor_out[11][4][14] + xor_out[12][4][14] + xor_out[13][4][14] + xor_out[14][4][14];
assign sum_out[3][4][14] = xor_out[15][4][14] + xor_out[16][4][14] + xor_out[17][4][14] + xor_out[18][4][14] + xor_out[19][4][14];
assign sum_out[4][4][14] = xor_out[20][4][14] + xor_out[21][4][14] + xor_out[22][4][14] + xor_out[23][4][14] + xor_out[24][4][14];
assign sum_out[5][4][14] = xor_out[25][4][14] + xor_out[26][4][14] + xor_out[27][4][14] + xor_out[28][4][14] + xor_out[29][4][14];
assign sum_out[6][4][14] = xor_out[30][4][14] + xor_out[31][4][14] + xor_out[32][4][14] + xor_out[33][4][14] + xor_out[34][4][14];
assign sum_out[7][4][14] = xor_out[35][4][14] + xor_out[36][4][14] + xor_out[37][4][14] + xor_out[38][4][14] + xor_out[39][4][14];
assign sum_out[8][4][14] = xor_out[40][4][14] + xor_out[41][4][14] + xor_out[42][4][14] + xor_out[43][4][14] + xor_out[44][4][14];
assign sum_out[9][4][14] = xor_out[45][4][14] + xor_out[46][4][14] + xor_out[47][4][14] + xor_out[48][4][14] + xor_out[49][4][14];
assign sum_out[10][4][14] = xor_out[50][4][14] + xor_out[51][4][14] + xor_out[52][4][14] + xor_out[53][4][14] + xor_out[54][4][14];
assign sum_out[11][4][14] = xor_out[55][4][14] + xor_out[56][4][14] + xor_out[57][4][14] + xor_out[58][4][14] + xor_out[59][4][14];
assign sum_out[12][4][14] = xor_out[60][4][14] + xor_out[61][4][14] + xor_out[62][4][14] + xor_out[63][4][14] + xor_out[64][4][14];
assign sum_out[13][4][14] = xor_out[65][4][14] + xor_out[66][4][14] + xor_out[67][4][14] + xor_out[68][4][14] + xor_out[69][4][14];
assign sum_out[14][4][14] = xor_out[70][4][14] + xor_out[71][4][14] + xor_out[72][4][14] + xor_out[73][4][14] + xor_out[74][4][14];
assign sum_out[15][4][14] = xor_out[75][4][14] + xor_out[76][4][14] + xor_out[77][4][14] + xor_out[78][4][14] + xor_out[79][4][14];
assign sum_out[16][4][14] = xor_out[80][4][14] + xor_out[81][4][14] + xor_out[82][4][14] + xor_out[83][4][14] + xor_out[84][4][14];
assign sum_out[17][4][14] = xor_out[85][4][14] + xor_out[86][4][14] + xor_out[87][4][14] + xor_out[88][4][14] + xor_out[89][4][14];
assign sum_out[18][4][14] = xor_out[90][4][14] + xor_out[91][4][14] + xor_out[92][4][14] + xor_out[93][4][14] + xor_out[94][4][14];
assign sum_out[19][4][14] = xor_out[95][4][14] + xor_out[96][4][14] + xor_out[97][4][14] + xor_out[98][4][14] + xor_out[99][4][14];

assign sum_out[0][4][15] = xor_out[0][4][15] + xor_out[1][4][15] + xor_out[2][4][15] + xor_out[3][4][15] + xor_out[4][4][15];
assign sum_out[1][4][15] = xor_out[5][4][15] + xor_out[6][4][15] + xor_out[7][4][15] + xor_out[8][4][15] + xor_out[9][4][15];
assign sum_out[2][4][15] = xor_out[10][4][15] + xor_out[11][4][15] + xor_out[12][4][15] + xor_out[13][4][15] + xor_out[14][4][15];
assign sum_out[3][4][15] = xor_out[15][4][15] + xor_out[16][4][15] + xor_out[17][4][15] + xor_out[18][4][15] + xor_out[19][4][15];
assign sum_out[4][4][15] = xor_out[20][4][15] + xor_out[21][4][15] + xor_out[22][4][15] + xor_out[23][4][15] + xor_out[24][4][15];
assign sum_out[5][4][15] = xor_out[25][4][15] + xor_out[26][4][15] + xor_out[27][4][15] + xor_out[28][4][15] + xor_out[29][4][15];
assign sum_out[6][4][15] = xor_out[30][4][15] + xor_out[31][4][15] + xor_out[32][4][15] + xor_out[33][4][15] + xor_out[34][4][15];
assign sum_out[7][4][15] = xor_out[35][4][15] + xor_out[36][4][15] + xor_out[37][4][15] + xor_out[38][4][15] + xor_out[39][4][15];
assign sum_out[8][4][15] = xor_out[40][4][15] + xor_out[41][4][15] + xor_out[42][4][15] + xor_out[43][4][15] + xor_out[44][4][15];
assign sum_out[9][4][15] = xor_out[45][4][15] + xor_out[46][4][15] + xor_out[47][4][15] + xor_out[48][4][15] + xor_out[49][4][15];
assign sum_out[10][4][15] = xor_out[50][4][15] + xor_out[51][4][15] + xor_out[52][4][15] + xor_out[53][4][15] + xor_out[54][4][15];
assign sum_out[11][4][15] = xor_out[55][4][15] + xor_out[56][4][15] + xor_out[57][4][15] + xor_out[58][4][15] + xor_out[59][4][15];
assign sum_out[12][4][15] = xor_out[60][4][15] + xor_out[61][4][15] + xor_out[62][4][15] + xor_out[63][4][15] + xor_out[64][4][15];
assign sum_out[13][4][15] = xor_out[65][4][15] + xor_out[66][4][15] + xor_out[67][4][15] + xor_out[68][4][15] + xor_out[69][4][15];
assign sum_out[14][4][15] = xor_out[70][4][15] + xor_out[71][4][15] + xor_out[72][4][15] + xor_out[73][4][15] + xor_out[74][4][15];
assign sum_out[15][4][15] = xor_out[75][4][15] + xor_out[76][4][15] + xor_out[77][4][15] + xor_out[78][4][15] + xor_out[79][4][15];
assign sum_out[16][4][15] = xor_out[80][4][15] + xor_out[81][4][15] + xor_out[82][4][15] + xor_out[83][4][15] + xor_out[84][4][15];
assign sum_out[17][4][15] = xor_out[85][4][15] + xor_out[86][4][15] + xor_out[87][4][15] + xor_out[88][4][15] + xor_out[89][4][15];
assign sum_out[18][4][15] = xor_out[90][4][15] + xor_out[91][4][15] + xor_out[92][4][15] + xor_out[93][4][15] + xor_out[94][4][15];
assign sum_out[19][4][15] = xor_out[95][4][15] + xor_out[96][4][15] + xor_out[97][4][15] + xor_out[98][4][15] + xor_out[99][4][15];

assign sum_out[0][4][16] = xor_out[0][4][16] + xor_out[1][4][16] + xor_out[2][4][16] + xor_out[3][4][16] + xor_out[4][4][16];
assign sum_out[1][4][16] = xor_out[5][4][16] + xor_out[6][4][16] + xor_out[7][4][16] + xor_out[8][4][16] + xor_out[9][4][16];
assign sum_out[2][4][16] = xor_out[10][4][16] + xor_out[11][4][16] + xor_out[12][4][16] + xor_out[13][4][16] + xor_out[14][4][16];
assign sum_out[3][4][16] = xor_out[15][4][16] + xor_out[16][4][16] + xor_out[17][4][16] + xor_out[18][4][16] + xor_out[19][4][16];
assign sum_out[4][4][16] = xor_out[20][4][16] + xor_out[21][4][16] + xor_out[22][4][16] + xor_out[23][4][16] + xor_out[24][4][16];
assign sum_out[5][4][16] = xor_out[25][4][16] + xor_out[26][4][16] + xor_out[27][4][16] + xor_out[28][4][16] + xor_out[29][4][16];
assign sum_out[6][4][16] = xor_out[30][4][16] + xor_out[31][4][16] + xor_out[32][4][16] + xor_out[33][4][16] + xor_out[34][4][16];
assign sum_out[7][4][16] = xor_out[35][4][16] + xor_out[36][4][16] + xor_out[37][4][16] + xor_out[38][4][16] + xor_out[39][4][16];
assign sum_out[8][4][16] = xor_out[40][4][16] + xor_out[41][4][16] + xor_out[42][4][16] + xor_out[43][4][16] + xor_out[44][4][16];
assign sum_out[9][4][16] = xor_out[45][4][16] + xor_out[46][4][16] + xor_out[47][4][16] + xor_out[48][4][16] + xor_out[49][4][16];
assign sum_out[10][4][16] = xor_out[50][4][16] + xor_out[51][4][16] + xor_out[52][4][16] + xor_out[53][4][16] + xor_out[54][4][16];
assign sum_out[11][4][16] = xor_out[55][4][16] + xor_out[56][4][16] + xor_out[57][4][16] + xor_out[58][4][16] + xor_out[59][4][16];
assign sum_out[12][4][16] = xor_out[60][4][16] + xor_out[61][4][16] + xor_out[62][4][16] + xor_out[63][4][16] + xor_out[64][4][16];
assign sum_out[13][4][16] = xor_out[65][4][16] + xor_out[66][4][16] + xor_out[67][4][16] + xor_out[68][4][16] + xor_out[69][4][16];
assign sum_out[14][4][16] = xor_out[70][4][16] + xor_out[71][4][16] + xor_out[72][4][16] + xor_out[73][4][16] + xor_out[74][4][16];
assign sum_out[15][4][16] = xor_out[75][4][16] + xor_out[76][4][16] + xor_out[77][4][16] + xor_out[78][4][16] + xor_out[79][4][16];
assign sum_out[16][4][16] = xor_out[80][4][16] + xor_out[81][4][16] + xor_out[82][4][16] + xor_out[83][4][16] + xor_out[84][4][16];
assign sum_out[17][4][16] = xor_out[85][4][16] + xor_out[86][4][16] + xor_out[87][4][16] + xor_out[88][4][16] + xor_out[89][4][16];
assign sum_out[18][4][16] = xor_out[90][4][16] + xor_out[91][4][16] + xor_out[92][4][16] + xor_out[93][4][16] + xor_out[94][4][16];
assign sum_out[19][4][16] = xor_out[95][4][16] + xor_out[96][4][16] + xor_out[97][4][16] + xor_out[98][4][16] + xor_out[99][4][16];

assign sum_out[0][4][17] = xor_out[0][4][17] + xor_out[1][4][17] + xor_out[2][4][17] + xor_out[3][4][17] + xor_out[4][4][17];
assign sum_out[1][4][17] = xor_out[5][4][17] + xor_out[6][4][17] + xor_out[7][4][17] + xor_out[8][4][17] + xor_out[9][4][17];
assign sum_out[2][4][17] = xor_out[10][4][17] + xor_out[11][4][17] + xor_out[12][4][17] + xor_out[13][4][17] + xor_out[14][4][17];
assign sum_out[3][4][17] = xor_out[15][4][17] + xor_out[16][4][17] + xor_out[17][4][17] + xor_out[18][4][17] + xor_out[19][4][17];
assign sum_out[4][4][17] = xor_out[20][4][17] + xor_out[21][4][17] + xor_out[22][4][17] + xor_out[23][4][17] + xor_out[24][4][17];
assign sum_out[5][4][17] = xor_out[25][4][17] + xor_out[26][4][17] + xor_out[27][4][17] + xor_out[28][4][17] + xor_out[29][4][17];
assign sum_out[6][4][17] = xor_out[30][4][17] + xor_out[31][4][17] + xor_out[32][4][17] + xor_out[33][4][17] + xor_out[34][4][17];
assign sum_out[7][4][17] = xor_out[35][4][17] + xor_out[36][4][17] + xor_out[37][4][17] + xor_out[38][4][17] + xor_out[39][4][17];
assign sum_out[8][4][17] = xor_out[40][4][17] + xor_out[41][4][17] + xor_out[42][4][17] + xor_out[43][4][17] + xor_out[44][4][17];
assign sum_out[9][4][17] = xor_out[45][4][17] + xor_out[46][4][17] + xor_out[47][4][17] + xor_out[48][4][17] + xor_out[49][4][17];
assign sum_out[10][4][17] = xor_out[50][4][17] + xor_out[51][4][17] + xor_out[52][4][17] + xor_out[53][4][17] + xor_out[54][4][17];
assign sum_out[11][4][17] = xor_out[55][4][17] + xor_out[56][4][17] + xor_out[57][4][17] + xor_out[58][4][17] + xor_out[59][4][17];
assign sum_out[12][4][17] = xor_out[60][4][17] + xor_out[61][4][17] + xor_out[62][4][17] + xor_out[63][4][17] + xor_out[64][4][17];
assign sum_out[13][4][17] = xor_out[65][4][17] + xor_out[66][4][17] + xor_out[67][4][17] + xor_out[68][4][17] + xor_out[69][4][17];
assign sum_out[14][4][17] = xor_out[70][4][17] + xor_out[71][4][17] + xor_out[72][4][17] + xor_out[73][4][17] + xor_out[74][4][17];
assign sum_out[15][4][17] = xor_out[75][4][17] + xor_out[76][4][17] + xor_out[77][4][17] + xor_out[78][4][17] + xor_out[79][4][17];
assign sum_out[16][4][17] = xor_out[80][4][17] + xor_out[81][4][17] + xor_out[82][4][17] + xor_out[83][4][17] + xor_out[84][4][17];
assign sum_out[17][4][17] = xor_out[85][4][17] + xor_out[86][4][17] + xor_out[87][4][17] + xor_out[88][4][17] + xor_out[89][4][17];
assign sum_out[18][4][17] = xor_out[90][4][17] + xor_out[91][4][17] + xor_out[92][4][17] + xor_out[93][4][17] + xor_out[94][4][17];
assign sum_out[19][4][17] = xor_out[95][4][17] + xor_out[96][4][17] + xor_out[97][4][17] + xor_out[98][4][17] + xor_out[99][4][17];

assign sum_out[0][4][18] = xor_out[0][4][18] + xor_out[1][4][18] + xor_out[2][4][18] + xor_out[3][4][18] + xor_out[4][4][18];
assign sum_out[1][4][18] = xor_out[5][4][18] + xor_out[6][4][18] + xor_out[7][4][18] + xor_out[8][4][18] + xor_out[9][4][18];
assign sum_out[2][4][18] = xor_out[10][4][18] + xor_out[11][4][18] + xor_out[12][4][18] + xor_out[13][4][18] + xor_out[14][4][18];
assign sum_out[3][4][18] = xor_out[15][4][18] + xor_out[16][4][18] + xor_out[17][4][18] + xor_out[18][4][18] + xor_out[19][4][18];
assign sum_out[4][4][18] = xor_out[20][4][18] + xor_out[21][4][18] + xor_out[22][4][18] + xor_out[23][4][18] + xor_out[24][4][18];
assign sum_out[5][4][18] = xor_out[25][4][18] + xor_out[26][4][18] + xor_out[27][4][18] + xor_out[28][4][18] + xor_out[29][4][18];
assign sum_out[6][4][18] = xor_out[30][4][18] + xor_out[31][4][18] + xor_out[32][4][18] + xor_out[33][4][18] + xor_out[34][4][18];
assign sum_out[7][4][18] = xor_out[35][4][18] + xor_out[36][4][18] + xor_out[37][4][18] + xor_out[38][4][18] + xor_out[39][4][18];
assign sum_out[8][4][18] = xor_out[40][4][18] + xor_out[41][4][18] + xor_out[42][4][18] + xor_out[43][4][18] + xor_out[44][4][18];
assign sum_out[9][4][18] = xor_out[45][4][18] + xor_out[46][4][18] + xor_out[47][4][18] + xor_out[48][4][18] + xor_out[49][4][18];
assign sum_out[10][4][18] = xor_out[50][4][18] + xor_out[51][4][18] + xor_out[52][4][18] + xor_out[53][4][18] + xor_out[54][4][18];
assign sum_out[11][4][18] = xor_out[55][4][18] + xor_out[56][4][18] + xor_out[57][4][18] + xor_out[58][4][18] + xor_out[59][4][18];
assign sum_out[12][4][18] = xor_out[60][4][18] + xor_out[61][4][18] + xor_out[62][4][18] + xor_out[63][4][18] + xor_out[64][4][18];
assign sum_out[13][4][18] = xor_out[65][4][18] + xor_out[66][4][18] + xor_out[67][4][18] + xor_out[68][4][18] + xor_out[69][4][18];
assign sum_out[14][4][18] = xor_out[70][4][18] + xor_out[71][4][18] + xor_out[72][4][18] + xor_out[73][4][18] + xor_out[74][4][18];
assign sum_out[15][4][18] = xor_out[75][4][18] + xor_out[76][4][18] + xor_out[77][4][18] + xor_out[78][4][18] + xor_out[79][4][18];
assign sum_out[16][4][18] = xor_out[80][4][18] + xor_out[81][4][18] + xor_out[82][4][18] + xor_out[83][4][18] + xor_out[84][4][18];
assign sum_out[17][4][18] = xor_out[85][4][18] + xor_out[86][4][18] + xor_out[87][4][18] + xor_out[88][4][18] + xor_out[89][4][18];
assign sum_out[18][4][18] = xor_out[90][4][18] + xor_out[91][4][18] + xor_out[92][4][18] + xor_out[93][4][18] + xor_out[94][4][18];
assign sum_out[19][4][18] = xor_out[95][4][18] + xor_out[96][4][18] + xor_out[97][4][18] + xor_out[98][4][18] + xor_out[99][4][18];

assign sum_out[0][4][19] = xor_out[0][4][19] + xor_out[1][4][19] + xor_out[2][4][19] + xor_out[3][4][19] + xor_out[4][4][19];
assign sum_out[1][4][19] = xor_out[5][4][19] + xor_out[6][4][19] + xor_out[7][4][19] + xor_out[8][4][19] + xor_out[9][4][19];
assign sum_out[2][4][19] = xor_out[10][4][19] + xor_out[11][4][19] + xor_out[12][4][19] + xor_out[13][4][19] + xor_out[14][4][19];
assign sum_out[3][4][19] = xor_out[15][4][19] + xor_out[16][4][19] + xor_out[17][4][19] + xor_out[18][4][19] + xor_out[19][4][19];
assign sum_out[4][4][19] = xor_out[20][4][19] + xor_out[21][4][19] + xor_out[22][4][19] + xor_out[23][4][19] + xor_out[24][4][19];
assign sum_out[5][4][19] = xor_out[25][4][19] + xor_out[26][4][19] + xor_out[27][4][19] + xor_out[28][4][19] + xor_out[29][4][19];
assign sum_out[6][4][19] = xor_out[30][4][19] + xor_out[31][4][19] + xor_out[32][4][19] + xor_out[33][4][19] + xor_out[34][4][19];
assign sum_out[7][4][19] = xor_out[35][4][19] + xor_out[36][4][19] + xor_out[37][4][19] + xor_out[38][4][19] + xor_out[39][4][19];
assign sum_out[8][4][19] = xor_out[40][4][19] + xor_out[41][4][19] + xor_out[42][4][19] + xor_out[43][4][19] + xor_out[44][4][19];
assign sum_out[9][4][19] = xor_out[45][4][19] + xor_out[46][4][19] + xor_out[47][4][19] + xor_out[48][4][19] + xor_out[49][4][19];
assign sum_out[10][4][19] = xor_out[50][4][19] + xor_out[51][4][19] + xor_out[52][4][19] + xor_out[53][4][19] + xor_out[54][4][19];
assign sum_out[11][4][19] = xor_out[55][4][19] + xor_out[56][4][19] + xor_out[57][4][19] + xor_out[58][4][19] + xor_out[59][4][19];
assign sum_out[12][4][19] = xor_out[60][4][19] + xor_out[61][4][19] + xor_out[62][4][19] + xor_out[63][4][19] + xor_out[64][4][19];
assign sum_out[13][4][19] = xor_out[65][4][19] + xor_out[66][4][19] + xor_out[67][4][19] + xor_out[68][4][19] + xor_out[69][4][19];
assign sum_out[14][4][19] = xor_out[70][4][19] + xor_out[71][4][19] + xor_out[72][4][19] + xor_out[73][4][19] + xor_out[74][4][19];
assign sum_out[15][4][19] = xor_out[75][4][19] + xor_out[76][4][19] + xor_out[77][4][19] + xor_out[78][4][19] + xor_out[79][4][19];
assign sum_out[16][4][19] = xor_out[80][4][19] + xor_out[81][4][19] + xor_out[82][4][19] + xor_out[83][4][19] + xor_out[84][4][19];
assign sum_out[17][4][19] = xor_out[85][4][19] + xor_out[86][4][19] + xor_out[87][4][19] + xor_out[88][4][19] + xor_out[89][4][19];
assign sum_out[18][4][19] = xor_out[90][4][19] + xor_out[91][4][19] + xor_out[92][4][19] + xor_out[93][4][19] + xor_out[94][4][19];
assign sum_out[19][4][19] = xor_out[95][4][19] + xor_out[96][4][19] + xor_out[97][4][19] + xor_out[98][4][19] + xor_out[99][4][19];

assign sum_out[0][4][20] = xor_out[0][4][20] + xor_out[1][4][20] + xor_out[2][4][20] + xor_out[3][4][20] + xor_out[4][4][20];
assign sum_out[1][4][20] = xor_out[5][4][20] + xor_out[6][4][20] + xor_out[7][4][20] + xor_out[8][4][20] + xor_out[9][4][20];
assign sum_out[2][4][20] = xor_out[10][4][20] + xor_out[11][4][20] + xor_out[12][4][20] + xor_out[13][4][20] + xor_out[14][4][20];
assign sum_out[3][4][20] = xor_out[15][4][20] + xor_out[16][4][20] + xor_out[17][4][20] + xor_out[18][4][20] + xor_out[19][4][20];
assign sum_out[4][4][20] = xor_out[20][4][20] + xor_out[21][4][20] + xor_out[22][4][20] + xor_out[23][4][20] + xor_out[24][4][20];
assign sum_out[5][4][20] = xor_out[25][4][20] + xor_out[26][4][20] + xor_out[27][4][20] + xor_out[28][4][20] + xor_out[29][4][20];
assign sum_out[6][4][20] = xor_out[30][4][20] + xor_out[31][4][20] + xor_out[32][4][20] + xor_out[33][4][20] + xor_out[34][4][20];
assign sum_out[7][4][20] = xor_out[35][4][20] + xor_out[36][4][20] + xor_out[37][4][20] + xor_out[38][4][20] + xor_out[39][4][20];
assign sum_out[8][4][20] = xor_out[40][4][20] + xor_out[41][4][20] + xor_out[42][4][20] + xor_out[43][4][20] + xor_out[44][4][20];
assign sum_out[9][4][20] = xor_out[45][4][20] + xor_out[46][4][20] + xor_out[47][4][20] + xor_out[48][4][20] + xor_out[49][4][20];
assign sum_out[10][4][20] = xor_out[50][4][20] + xor_out[51][4][20] + xor_out[52][4][20] + xor_out[53][4][20] + xor_out[54][4][20];
assign sum_out[11][4][20] = xor_out[55][4][20] + xor_out[56][4][20] + xor_out[57][4][20] + xor_out[58][4][20] + xor_out[59][4][20];
assign sum_out[12][4][20] = xor_out[60][4][20] + xor_out[61][4][20] + xor_out[62][4][20] + xor_out[63][4][20] + xor_out[64][4][20];
assign sum_out[13][4][20] = xor_out[65][4][20] + xor_out[66][4][20] + xor_out[67][4][20] + xor_out[68][4][20] + xor_out[69][4][20];
assign sum_out[14][4][20] = xor_out[70][4][20] + xor_out[71][4][20] + xor_out[72][4][20] + xor_out[73][4][20] + xor_out[74][4][20];
assign sum_out[15][4][20] = xor_out[75][4][20] + xor_out[76][4][20] + xor_out[77][4][20] + xor_out[78][4][20] + xor_out[79][4][20];
assign sum_out[16][4][20] = xor_out[80][4][20] + xor_out[81][4][20] + xor_out[82][4][20] + xor_out[83][4][20] + xor_out[84][4][20];
assign sum_out[17][4][20] = xor_out[85][4][20] + xor_out[86][4][20] + xor_out[87][4][20] + xor_out[88][4][20] + xor_out[89][4][20];
assign sum_out[18][4][20] = xor_out[90][4][20] + xor_out[91][4][20] + xor_out[92][4][20] + xor_out[93][4][20] + xor_out[94][4][20];
assign sum_out[19][4][20] = xor_out[95][4][20] + xor_out[96][4][20] + xor_out[97][4][20] + xor_out[98][4][20] + xor_out[99][4][20];

assign sum_out[0][4][21] = xor_out[0][4][21] + xor_out[1][4][21] + xor_out[2][4][21] + xor_out[3][4][21] + xor_out[4][4][21];
assign sum_out[1][4][21] = xor_out[5][4][21] + xor_out[6][4][21] + xor_out[7][4][21] + xor_out[8][4][21] + xor_out[9][4][21];
assign sum_out[2][4][21] = xor_out[10][4][21] + xor_out[11][4][21] + xor_out[12][4][21] + xor_out[13][4][21] + xor_out[14][4][21];
assign sum_out[3][4][21] = xor_out[15][4][21] + xor_out[16][4][21] + xor_out[17][4][21] + xor_out[18][4][21] + xor_out[19][4][21];
assign sum_out[4][4][21] = xor_out[20][4][21] + xor_out[21][4][21] + xor_out[22][4][21] + xor_out[23][4][21] + xor_out[24][4][21];
assign sum_out[5][4][21] = xor_out[25][4][21] + xor_out[26][4][21] + xor_out[27][4][21] + xor_out[28][4][21] + xor_out[29][4][21];
assign sum_out[6][4][21] = xor_out[30][4][21] + xor_out[31][4][21] + xor_out[32][4][21] + xor_out[33][4][21] + xor_out[34][4][21];
assign sum_out[7][4][21] = xor_out[35][4][21] + xor_out[36][4][21] + xor_out[37][4][21] + xor_out[38][4][21] + xor_out[39][4][21];
assign sum_out[8][4][21] = xor_out[40][4][21] + xor_out[41][4][21] + xor_out[42][4][21] + xor_out[43][4][21] + xor_out[44][4][21];
assign sum_out[9][4][21] = xor_out[45][4][21] + xor_out[46][4][21] + xor_out[47][4][21] + xor_out[48][4][21] + xor_out[49][4][21];
assign sum_out[10][4][21] = xor_out[50][4][21] + xor_out[51][4][21] + xor_out[52][4][21] + xor_out[53][4][21] + xor_out[54][4][21];
assign sum_out[11][4][21] = xor_out[55][4][21] + xor_out[56][4][21] + xor_out[57][4][21] + xor_out[58][4][21] + xor_out[59][4][21];
assign sum_out[12][4][21] = xor_out[60][4][21] + xor_out[61][4][21] + xor_out[62][4][21] + xor_out[63][4][21] + xor_out[64][4][21];
assign sum_out[13][4][21] = xor_out[65][4][21] + xor_out[66][4][21] + xor_out[67][4][21] + xor_out[68][4][21] + xor_out[69][4][21];
assign sum_out[14][4][21] = xor_out[70][4][21] + xor_out[71][4][21] + xor_out[72][4][21] + xor_out[73][4][21] + xor_out[74][4][21];
assign sum_out[15][4][21] = xor_out[75][4][21] + xor_out[76][4][21] + xor_out[77][4][21] + xor_out[78][4][21] + xor_out[79][4][21];
assign sum_out[16][4][21] = xor_out[80][4][21] + xor_out[81][4][21] + xor_out[82][4][21] + xor_out[83][4][21] + xor_out[84][4][21];
assign sum_out[17][4][21] = xor_out[85][4][21] + xor_out[86][4][21] + xor_out[87][4][21] + xor_out[88][4][21] + xor_out[89][4][21];
assign sum_out[18][4][21] = xor_out[90][4][21] + xor_out[91][4][21] + xor_out[92][4][21] + xor_out[93][4][21] + xor_out[94][4][21];
assign sum_out[19][4][21] = xor_out[95][4][21] + xor_out[96][4][21] + xor_out[97][4][21] + xor_out[98][4][21] + xor_out[99][4][21];

assign sum_out[0][4][22] = xor_out[0][4][22] + xor_out[1][4][22] + xor_out[2][4][22] + xor_out[3][4][22] + xor_out[4][4][22];
assign sum_out[1][4][22] = xor_out[5][4][22] + xor_out[6][4][22] + xor_out[7][4][22] + xor_out[8][4][22] + xor_out[9][4][22];
assign sum_out[2][4][22] = xor_out[10][4][22] + xor_out[11][4][22] + xor_out[12][4][22] + xor_out[13][4][22] + xor_out[14][4][22];
assign sum_out[3][4][22] = xor_out[15][4][22] + xor_out[16][4][22] + xor_out[17][4][22] + xor_out[18][4][22] + xor_out[19][4][22];
assign sum_out[4][4][22] = xor_out[20][4][22] + xor_out[21][4][22] + xor_out[22][4][22] + xor_out[23][4][22] + xor_out[24][4][22];
assign sum_out[5][4][22] = xor_out[25][4][22] + xor_out[26][4][22] + xor_out[27][4][22] + xor_out[28][4][22] + xor_out[29][4][22];
assign sum_out[6][4][22] = xor_out[30][4][22] + xor_out[31][4][22] + xor_out[32][4][22] + xor_out[33][4][22] + xor_out[34][4][22];
assign sum_out[7][4][22] = xor_out[35][4][22] + xor_out[36][4][22] + xor_out[37][4][22] + xor_out[38][4][22] + xor_out[39][4][22];
assign sum_out[8][4][22] = xor_out[40][4][22] + xor_out[41][4][22] + xor_out[42][4][22] + xor_out[43][4][22] + xor_out[44][4][22];
assign sum_out[9][4][22] = xor_out[45][4][22] + xor_out[46][4][22] + xor_out[47][4][22] + xor_out[48][4][22] + xor_out[49][4][22];
assign sum_out[10][4][22] = xor_out[50][4][22] + xor_out[51][4][22] + xor_out[52][4][22] + xor_out[53][4][22] + xor_out[54][4][22];
assign sum_out[11][4][22] = xor_out[55][4][22] + xor_out[56][4][22] + xor_out[57][4][22] + xor_out[58][4][22] + xor_out[59][4][22];
assign sum_out[12][4][22] = xor_out[60][4][22] + xor_out[61][4][22] + xor_out[62][4][22] + xor_out[63][4][22] + xor_out[64][4][22];
assign sum_out[13][4][22] = xor_out[65][4][22] + xor_out[66][4][22] + xor_out[67][4][22] + xor_out[68][4][22] + xor_out[69][4][22];
assign sum_out[14][4][22] = xor_out[70][4][22] + xor_out[71][4][22] + xor_out[72][4][22] + xor_out[73][4][22] + xor_out[74][4][22];
assign sum_out[15][4][22] = xor_out[75][4][22] + xor_out[76][4][22] + xor_out[77][4][22] + xor_out[78][4][22] + xor_out[79][4][22];
assign sum_out[16][4][22] = xor_out[80][4][22] + xor_out[81][4][22] + xor_out[82][4][22] + xor_out[83][4][22] + xor_out[84][4][22];
assign sum_out[17][4][22] = xor_out[85][4][22] + xor_out[86][4][22] + xor_out[87][4][22] + xor_out[88][4][22] + xor_out[89][4][22];
assign sum_out[18][4][22] = xor_out[90][4][22] + xor_out[91][4][22] + xor_out[92][4][22] + xor_out[93][4][22] + xor_out[94][4][22];
assign sum_out[19][4][22] = xor_out[95][4][22] + xor_out[96][4][22] + xor_out[97][4][22] + xor_out[98][4][22] + xor_out[99][4][22];

assign sum_out[0][4][23] = xor_out[0][4][23] + xor_out[1][4][23] + xor_out[2][4][23] + xor_out[3][4][23] + xor_out[4][4][23];
assign sum_out[1][4][23] = xor_out[5][4][23] + xor_out[6][4][23] + xor_out[7][4][23] + xor_out[8][4][23] + xor_out[9][4][23];
assign sum_out[2][4][23] = xor_out[10][4][23] + xor_out[11][4][23] + xor_out[12][4][23] + xor_out[13][4][23] + xor_out[14][4][23];
assign sum_out[3][4][23] = xor_out[15][4][23] + xor_out[16][4][23] + xor_out[17][4][23] + xor_out[18][4][23] + xor_out[19][4][23];
assign sum_out[4][4][23] = xor_out[20][4][23] + xor_out[21][4][23] + xor_out[22][4][23] + xor_out[23][4][23] + xor_out[24][4][23];
assign sum_out[5][4][23] = xor_out[25][4][23] + xor_out[26][4][23] + xor_out[27][4][23] + xor_out[28][4][23] + xor_out[29][4][23];
assign sum_out[6][4][23] = xor_out[30][4][23] + xor_out[31][4][23] + xor_out[32][4][23] + xor_out[33][4][23] + xor_out[34][4][23];
assign sum_out[7][4][23] = xor_out[35][4][23] + xor_out[36][4][23] + xor_out[37][4][23] + xor_out[38][4][23] + xor_out[39][4][23];
assign sum_out[8][4][23] = xor_out[40][4][23] + xor_out[41][4][23] + xor_out[42][4][23] + xor_out[43][4][23] + xor_out[44][4][23];
assign sum_out[9][4][23] = xor_out[45][4][23] + xor_out[46][4][23] + xor_out[47][4][23] + xor_out[48][4][23] + xor_out[49][4][23];
assign sum_out[10][4][23] = xor_out[50][4][23] + xor_out[51][4][23] + xor_out[52][4][23] + xor_out[53][4][23] + xor_out[54][4][23];
assign sum_out[11][4][23] = xor_out[55][4][23] + xor_out[56][4][23] + xor_out[57][4][23] + xor_out[58][4][23] + xor_out[59][4][23];
assign sum_out[12][4][23] = xor_out[60][4][23] + xor_out[61][4][23] + xor_out[62][4][23] + xor_out[63][4][23] + xor_out[64][4][23];
assign sum_out[13][4][23] = xor_out[65][4][23] + xor_out[66][4][23] + xor_out[67][4][23] + xor_out[68][4][23] + xor_out[69][4][23];
assign sum_out[14][4][23] = xor_out[70][4][23] + xor_out[71][4][23] + xor_out[72][4][23] + xor_out[73][4][23] + xor_out[74][4][23];
assign sum_out[15][4][23] = xor_out[75][4][23] + xor_out[76][4][23] + xor_out[77][4][23] + xor_out[78][4][23] + xor_out[79][4][23];
assign sum_out[16][4][23] = xor_out[80][4][23] + xor_out[81][4][23] + xor_out[82][4][23] + xor_out[83][4][23] + xor_out[84][4][23];
assign sum_out[17][4][23] = xor_out[85][4][23] + xor_out[86][4][23] + xor_out[87][4][23] + xor_out[88][4][23] + xor_out[89][4][23];
assign sum_out[18][4][23] = xor_out[90][4][23] + xor_out[91][4][23] + xor_out[92][4][23] + xor_out[93][4][23] + xor_out[94][4][23];
assign sum_out[19][4][23] = xor_out[95][4][23] + xor_out[96][4][23] + xor_out[97][4][23] + xor_out[98][4][23] + xor_out[99][4][23];

assign sum_out[0][5][0] = xor_out[0][5][0] + xor_out[1][5][0] + xor_out[2][5][0] + xor_out[3][5][0] + xor_out[4][5][0];
assign sum_out[1][5][0] = xor_out[5][5][0] + xor_out[6][5][0] + xor_out[7][5][0] + xor_out[8][5][0] + xor_out[9][5][0];
assign sum_out[2][5][0] = xor_out[10][5][0] + xor_out[11][5][0] + xor_out[12][5][0] + xor_out[13][5][0] + xor_out[14][5][0];
assign sum_out[3][5][0] = xor_out[15][5][0] + xor_out[16][5][0] + xor_out[17][5][0] + xor_out[18][5][0] + xor_out[19][5][0];
assign sum_out[4][5][0] = xor_out[20][5][0] + xor_out[21][5][0] + xor_out[22][5][0] + xor_out[23][5][0] + xor_out[24][5][0];
assign sum_out[5][5][0] = xor_out[25][5][0] + xor_out[26][5][0] + xor_out[27][5][0] + xor_out[28][5][0] + xor_out[29][5][0];
assign sum_out[6][5][0] = xor_out[30][5][0] + xor_out[31][5][0] + xor_out[32][5][0] + xor_out[33][5][0] + xor_out[34][5][0];
assign sum_out[7][5][0] = xor_out[35][5][0] + xor_out[36][5][0] + xor_out[37][5][0] + xor_out[38][5][0] + xor_out[39][5][0];
assign sum_out[8][5][0] = xor_out[40][5][0] + xor_out[41][5][0] + xor_out[42][5][0] + xor_out[43][5][0] + xor_out[44][5][0];
assign sum_out[9][5][0] = xor_out[45][5][0] + xor_out[46][5][0] + xor_out[47][5][0] + xor_out[48][5][0] + xor_out[49][5][0];
assign sum_out[10][5][0] = xor_out[50][5][0] + xor_out[51][5][0] + xor_out[52][5][0] + xor_out[53][5][0] + xor_out[54][5][0];
assign sum_out[11][5][0] = xor_out[55][5][0] + xor_out[56][5][0] + xor_out[57][5][0] + xor_out[58][5][0] + xor_out[59][5][0];
assign sum_out[12][5][0] = xor_out[60][5][0] + xor_out[61][5][0] + xor_out[62][5][0] + xor_out[63][5][0] + xor_out[64][5][0];
assign sum_out[13][5][0] = xor_out[65][5][0] + xor_out[66][5][0] + xor_out[67][5][0] + xor_out[68][5][0] + xor_out[69][5][0];
assign sum_out[14][5][0] = xor_out[70][5][0] + xor_out[71][5][0] + xor_out[72][5][0] + xor_out[73][5][0] + xor_out[74][5][0];
assign sum_out[15][5][0] = xor_out[75][5][0] + xor_out[76][5][0] + xor_out[77][5][0] + xor_out[78][5][0] + xor_out[79][5][0];
assign sum_out[16][5][0] = xor_out[80][5][0] + xor_out[81][5][0] + xor_out[82][5][0] + xor_out[83][5][0] + xor_out[84][5][0];
assign sum_out[17][5][0] = xor_out[85][5][0] + xor_out[86][5][0] + xor_out[87][5][0] + xor_out[88][5][0] + xor_out[89][5][0];
assign sum_out[18][5][0] = xor_out[90][5][0] + xor_out[91][5][0] + xor_out[92][5][0] + xor_out[93][5][0] + xor_out[94][5][0];
assign sum_out[19][5][0] = xor_out[95][5][0] + xor_out[96][5][0] + xor_out[97][5][0] + xor_out[98][5][0] + xor_out[99][5][0];

assign sum_out[0][5][1] = xor_out[0][5][1] + xor_out[1][5][1] + xor_out[2][5][1] + xor_out[3][5][1] + xor_out[4][5][1];
assign sum_out[1][5][1] = xor_out[5][5][1] + xor_out[6][5][1] + xor_out[7][5][1] + xor_out[8][5][1] + xor_out[9][5][1];
assign sum_out[2][5][1] = xor_out[10][5][1] + xor_out[11][5][1] + xor_out[12][5][1] + xor_out[13][5][1] + xor_out[14][5][1];
assign sum_out[3][5][1] = xor_out[15][5][1] + xor_out[16][5][1] + xor_out[17][5][1] + xor_out[18][5][1] + xor_out[19][5][1];
assign sum_out[4][5][1] = xor_out[20][5][1] + xor_out[21][5][1] + xor_out[22][5][1] + xor_out[23][5][1] + xor_out[24][5][1];
assign sum_out[5][5][1] = xor_out[25][5][1] + xor_out[26][5][1] + xor_out[27][5][1] + xor_out[28][5][1] + xor_out[29][5][1];
assign sum_out[6][5][1] = xor_out[30][5][1] + xor_out[31][5][1] + xor_out[32][5][1] + xor_out[33][5][1] + xor_out[34][5][1];
assign sum_out[7][5][1] = xor_out[35][5][1] + xor_out[36][5][1] + xor_out[37][5][1] + xor_out[38][5][1] + xor_out[39][5][1];
assign sum_out[8][5][1] = xor_out[40][5][1] + xor_out[41][5][1] + xor_out[42][5][1] + xor_out[43][5][1] + xor_out[44][5][1];
assign sum_out[9][5][1] = xor_out[45][5][1] + xor_out[46][5][1] + xor_out[47][5][1] + xor_out[48][5][1] + xor_out[49][5][1];
assign sum_out[10][5][1] = xor_out[50][5][1] + xor_out[51][5][1] + xor_out[52][5][1] + xor_out[53][5][1] + xor_out[54][5][1];
assign sum_out[11][5][1] = xor_out[55][5][1] + xor_out[56][5][1] + xor_out[57][5][1] + xor_out[58][5][1] + xor_out[59][5][1];
assign sum_out[12][5][1] = xor_out[60][5][1] + xor_out[61][5][1] + xor_out[62][5][1] + xor_out[63][5][1] + xor_out[64][5][1];
assign sum_out[13][5][1] = xor_out[65][5][1] + xor_out[66][5][1] + xor_out[67][5][1] + xor_out[68][5][1] + xor_out[69][5][1];
assign sum_out[14][5][1] = xor_out[70][5][1] + xor_out[71][5][1] + xor_out[72][5][1] + xor_out[73][5][1] + xor_out[74][5][1];
assign sum_out[15][5][1] = xor_out[75][5][1] + xor_out[76][5][1] + xor_out[77][5][1] + xor_out[78][5][1] + xor_out[79][5][1];
assign sum_out[16][5][1] = xor_out[80][5][1] + xor_out[81][5][1] + xor_out[82][5][1] + xor_out[83][5][1] + xor_out[84][5][1];
assign sum_out[17][5][1] = xor_out[85][5][1] + xor_out[86][5][1] + xor_out[87][5][1] + xor_out[88][5][1] + xor_out[89][5][1];
assign sum_out[18][5][1] = xor_out[90][5][1] + xor_out[91][5][1] + xor_out[92][5][1] + xor_out[93][5][1] + xor_out[94][5][1];
assign sum_out[19][5][1] = xor_out[95][5][1] + xor_out[96][5][1] + xor_out[97][5][1] + xor_out[98][5][1] + xor_out[99][5][1];

assign sum_out[0][5][2] = xor_out[0][5][2] + xor_out[1][5][2] + xor_out[2][5][2] + xor_out[3][5][2] + xor_out[4][5][2];
assign sum_out[1][5][2] = xor_out[5][5][2] + xor_out[6][5][2] + xor_out[7][5][2] + xor_out[8][5][2] + xor_out[9][5][2];
assign sum_out[2][5][2] = xor_out[10][5][2] + xor_out[11][5][2] + xor_out[12][5][2] + xor_out[13][5][2] + xor_out[14][5][2];
assign sum_out[3][5][2] = xor_out[15][5][2] + xor_out[16][5][2] + xor_out[17][5][2] + xor_out[18][5][2] + xor_out[19][5][2];
assign sum_out[4][5][2] = xor_out[20][5][2] + xor_out[21][5][2] + xor_out[22][5][2] + xor_out[23][5][2] + xor_out[24][5][2];
assign sum_out[5][5][2] = xor_out[25][5][2] + xor_out[26][5][2] + xor_out[27][5][2] + xor_out[28][5][2] + xor_out[29][5][2];
assign sum_out[6][5][2] = xor_out[30][5][2] + xor_out[31][5][2] + xor_out[32][5][2] + xor_out[33][5][2] + xor_out[34][5][2];
assign sum_out[7][5][2] = xor_out[35][5][2] + xor_out[36][5][2] + xor_out[37][5][2] + xor_out[38][5][2] + xor_out[39][5][2];
assign sum_out[8][5][2] = xor_out[40][5][2] + xor_out[41][5][2] + xor_out[42][5][2] + xor_out[43][5][2] + xor_out[44][5][2];
assign sum_out[9][5][2] = xor_out[45][5][2] + xor_out[46][5][2] + xor_out[47][5][2] + xor_out[48][5][2] + xor_out[49][5][2];
assign sum_out[10][5][2] = xor_out[50][5][2] + xor_out[51][5][2] + xor_out[52][5][2] + xor_out[53][5][2] + xor_out[54][5][2];
assign sum_out[11][5][2] = xor_out[55][5][2] + xor_out[56][5][2] + xor_out[57][5][2] + xor_out[58][5][2] + xor_out[59][5][2];
assign sum_out[12][5][2] = xor_out[60][5][2] + xor_out[61][5][2] + xor_out[62][5][2] + xor_out[63][5][2] + xor_out[64][5][2];
assign sum_out[13][5][2] = xor_out[65][5][2] + xor_out[66][5][2] + xor_out[67][5][2] + xor_out[68][5][2] + xor_out[69][5][2];
assign sum_out[14][5][2] = xor_out[70][5][2] + xor_out[71][5][2] + xor_out[72][5][2] + xor_out[73][5][2] + xor_out[74][5][2];
assign sum_out[15][5][2] = xor_out[75][5][2] + xor_out[76][5][2] + xor_out[77][5][2] + xor_out[78][5][2] + xor_out[79][5][2];
assign sum_out[16][5][2] = xor_out[80][5][2] + xor_out[81][5][2] + xor_out[82][5][2] + xor_out[83][5][2] + xor_out[84][5][2];
assign sum_out[17][5][2] = xor_out[85][5][2] + xor_out[86][5][2] + xor_out[87][5][2] + xor_out[88][5][2] + xor_out[89][5][2];
assign sum_out[18][5][2] = xor_out[90][5][2] + xor_out[91][5][2] + xor_out[92][5][2] + xor_out[93][5][2] + xor_out[94][5][2];
assign sum_out[19][5][2] = xor_out[95][5][2] + xor_out[96][5][2] + xor_out[97][5][2] + xor_out[98][5][2] + xor_out[99][5][2];

assign sum_out[0][5][3] = xor_out[0][5][3] + xor_out[1][5][3] + xor_out[2][5][3] + xor_out[3][5][3] + xor_out[4][5][3];
assign sum_out[1][5][3] = xor_out[5][5][3] + xor_out[6][5][3] + xor_out[7][5][3] + xor_out[8][5][3] + xor_out[9][5][3];
assign sum_out[2][5][3] = xor_out[10][5][3] + xor_out[11][5][3] + xor_out[12][5][3] + xor_out[13][5][3] + xor_out[14][5][3];
assign sum_out[3][5][3] = xor_out[15][5][3] + xor_out[16][5][3] + xor_out[17][5][3] + xor_out[18][5][3] + xor_out[19][5][3];
assign sum_out[4][5][3] = xor_out[20][5][3] + xor_out[21][5][3] + xor_out[22][5][3] + xor_out[23][5][3] + xor_out[24][5][3];
assign sum_out[5][5][3] = xor_out[25][5][3] + xor_out[26][5][3] + xor_out[27][5][3] + xor_out[28][5][3] + xor_out[29][5][3];
assign sum_out[6][5][3] = xor_out[30][5][3] + xor_out[31][5][3] + xor_out[32][5][3] + xor_out[33][5][3] + xor_out[34][5][3];
assign sum_out[7][5][3] = xor_out[35][5][3] + xor_out[36][5][3] + xor_out[37][5][3] + xor_out[38][5][3] + xor_out[39][5][3];
assign sum_out[8][5][3] = xor_out[40][5][3] + xor_out[41][5][3] + xor_out[42][5][3] + xor_out[43][5][3] + xor_out[44][5][3];
assign sum_out[9][5][3] = xor_out[45][5][3] + xor_out[46][5][3] + xor_out[47][5][3] + xor_out[48][5][3] + xor_out[49][5][3];
assign sum_out[10][5][3] = xor_out[50][5][3] + xor_out[51][5][3] + xor_out[52][5][3] + xor_out[53][5][3] + xor_out[54][5][3];
assign sum_out[11][5][3] = xor_out[55][5][3] + xor_out[56][5][3] + xor_out[57][5][3] + xor_out[58][5][3] + xor_out[59][5][3];
assign sum_out[12][5][3] = xor_out[60][5][3] + xor_out[61][5][3] + xor_out[62][5][3] + xor_out[63][5][3] + xor_out[64][5][3];
assign sum_out[13][5][3] = xor_out[65][5][3] + xor_out[66][5][3] + xor_out[67][5][3] + xor_out[68][5][3] + xor_out[69][5][3];
assign sum_out[14][5][3] = xor_out[70][5][3] + xor_out[71][5][3] + xor_out[72][5][3] + xor_out[73][5][3] + xor_out[74][5][3];
assign sum_out[15][5][3] = xor_out[75][5][3] + xor_out[76][5][3] + xor_out[77][5][3] + xor_out[78][5][3] + xor_out[79][5][3];
assign sum_out[16][5][3] = xor_out[80][5][3] + xor_out[81][5][3] + xor_out[82][5][3] + xor_out[83][5][3] + xor_out[84][5][3];
assign sum_out[17][5][3] = xor_out[85][5][3] + xor_out[86][5][3] + xor_out[87][5][3] + xor_out[88][5][3] + xor_out[89][5][3];
assign sum_out[18][5][3] = xor_out[90][5][3] + xor_out[91][5][3] + xor_out[92][5][3] + xor_out[93][5][3] + xor_out[94][5][3];
assign sum_out[19][5][3] = xor_out[95][5][3] + xor_out[96][5][3] + xor_out[97][5][3] + xor_out[98][5][3] + xor_out[99][5][3];

assign sum_out[0][5][4] = xor_out[0][5][4] + xor_out[1][5][4] + xor_out[2][5][4] + xor_out[3][5][4] + xor_out[4][5][4];
assign sum_out[1][5][4] = xor_out[5][5][4] + xor_out[6][5][4] + xor_out[7][5][4] + xor_out[8][5][4] + xor_out[9][5][4];
assign sum_out[2][5][4] = xor_out[10][5][4] + xor_out[11][5][4] + xor_out[12][5][4] + xor_out[13][5][4] + xor_out[14][5][4];
assign sum_out[3][5][4] = xor_out[15][5][4] + xor_out[16][5][4] + xor_out[17][5][4] + xor_out[18][5][4] + xor_out[19][5][4];
assign sum_out[4][5][4] = xor_out[20][5][4] + xor_out[21][5][4] + xor_out[22][5][4] + xor_out[23][5][4] + xor_out[24][5][4];
assign sum_out[5][5][4] = xor_out[25][5][4] + xor_out[26][5][4] + xor_out[27][5][4] + xor_out[28][5][4] + xor_out[29][5][4];
assign sum_out[6][5][4] = xor_out[30][5][4] + xor_out[31][5][4] + xor_out[32][5][4] + xor_out[33][5][4] + xor_out[34][5][4];
assign sum_out[7][5][4] = xor_out[35][5][4] + xor_out[36][5][4] + xor_out[37][5][4] + xor_out[38][5][4] + xor_out[39][5][4];
assign sum_out[8][5][4] = xor_out[40][5][4] + xor_out[41][5][4] + xor_out[42][5][4] + xor_out[43][5][4] + xor_out[44][5][4];
assign sum_out[9][5][4] = xor_out[45][5][4] + xor_out[46][5][4] + xor_out[47][5][4] + xor_out[48][5][4] + xor_out[49][5][4];
assign sum_out[10][5][4] = xor_out[50][5][4] + xor_out[51][5][4] + xor_out[52][5][4] + xor_out[53][5][4] + xor_out[54][5][4];
assign sum_out[11][5][4] = xor_out[55][5][4] + xor_out[56][5][4] + xor_out[57][5][4] + xor_out[58][5][4] + xor_out[59][5][4];
assign sum_out[12][5][4] = xor_out[60][5][4] + xor_out[61][5][4] + xor_out[62][5][4] + xor_out[63][5][4] + xor_out[64][5][4];
assign sum_out[13][5][4] = xor_out[65][5][4] + xor_out[66][5][4] + xor_out[67][5][4] + xor_out[68][5][4] + xor_out[69][5][4];
assign sum_out[14][5][4] = xor_out[70][5][4] + xor_out[71][5][4] + xor_out[72][5][4] + xor_out[73][5][4] + xor_out[74][5][4];
assign sum_out[15][5][4] = xor_out[75][5][4] + xor_out[76][5][4] + xor_out[77][5][4] + xor_out[78][5][4] + xor_out[79][5][4];
assign sum_out[16][5][4] = xor_out[80][5][4] + xor_out[81][5][4] + xor_out[82][5][4] + xor_out[83][5][4] + xor_out[84][5][4];
assign sum_out[17][5][4] = xor_out[85][5][4] + xor_out[86][5][4] + xor_out[87][5][4] + xor_out[88][5][4] + xor_out[89][5][4];
assign sum_out[18][5][4] = xor_out[90][5][4] + xor_out[91][5][4] + xor_out[92][5][4] + xor_out[93][5][4] + xor_out[94][5][4];
assign sum_out[19][5][4] = xor_out[95][5][4] + xor_out[96][5][4] + xor_out[97][5][4] + xor_out[98][5][4] + xor_out[99][5][4];

assign sum_out[0][5][5] = xor_out[0][5][5] + xor_out[1][5][5] + xor_out[2][5][5] + xor_out[3][5][5] + xor_out[4][5][5];
assign sum_out[1][5][5] = xor_out[5][5][5] + xor_out[6][5][5] + xor_out[7][5][5] + xor_out[8][5][5] + xor_out[9][5][5];
assign sum_out[2][5][5] = xor_out[10][5][5] + xor_out[11][5][5] + xor_out[12][5][5] + xor_out[13][5][5] + xor_out[14][5][5];
assign sum_out[3][5][5] = xor_out[15][5][5] + xor_out[16][5][5] + xor_out[17][5][5] + xor_out[18][5][5] + xor_out[19][5][5];
assign sum_out[4][5][5] = xor_out[20][5][5] + xor_out[21][5][5] + xor_out[22][5][5] + xor_out[23][5][5] + xor_out[24][5][5];
assign sum_out[5][5][5] = xor_out[25][5][5] + xor_out[26][5][5] + xor_out[27][5][5] + xor_out[28][5][5] + xor_out[29][5][5];
assign sum_out[6][5][5] = xor_out[30][5][5] + xor_out[31][5][5] + xor_out[32][5][5] + xor_out[33][5][5] + xor_out[34][5][5];
assign sum_out[7][5][5] = xor_out[35][5][5] + xor_out[36][5][5] + xor_out[37][5][5] + xor_out[38][5][5] + xor_out[39][5][5];
assign sum_out[8][5][5] = xor_out[40][5][5] + xor_out[41][5][5] + xor_out[42][5][5] + xor_out[43][5][5] + xor_out[44][5][5];
assign sum_out[9][5][5] = xor_out[45][5][5] + xor_out[46][5][5] + xor_out[47][5][5] + xor_out[48][5][5] + xor_out[49][5][5];
assign sum_out[10][5][5] = xor_out[50][5][5] + xor_out[51][5][5] + xor_out[52][5][5] + xor_out[53][5][5] + xor_out[54][5][5];
assign sum_out[11][5][5] = xor_out[55][5][5] + xor_out[56][5][5] + xor_out[57][5][5] + xor_out[58][5][5] + xor_out[59][5][5];
assign sum_out[12][5][5] = xor_out[60][5][5] + xor_out[61][5][5] + xor_out[62][5][5] + xor_out[63][5][5] + xor_out[64][5][5];
assign sum_out[13][5][5] = xor_out[65][5][5] + xor_out[66][5][5] + xor_out[67][5][5] + xor_out[68][5][5] + xor_out[69][5][5];
assign sum_out[14][5][5] = xor_out[70][5][5] + xor_out[71][5][5] + xor_out[72][5][5] + xor_out[73][5][5] + xor_out[74][5][5];
assign sum_out[15][5][5] = xor_out[75][5][5] + xor_out[76][5][5] + xor_out[77][5][5] + xor_out[78][5][5] + xor_out[79][5][5];
assign sum_out[16][5][5] = xor_out[80][5][5] + xor_out[81][5][5] + xor_out[82][5][5] + xor_out[83][5][5] + xor_out[84][5][5];
assign sum_out[17][5][5] = xor_out[85][5][5] + xor_out[86][5][5] + xor_out[87][5][5] + xor_out[88][5][5] + xor_out[89][5][5];
assign sum_out[18][5][5] = xor_out[90][5][5] + xor_out[91][5][5] + xor_out[92][5][5] + xor_out[93][5][5] + xor_out[94][5][5];
assign sum_out[19][5][5] = xor_out[95][5][5] + xor_out[96][5][5] + xor_out[97][5][5] + xor_out[98][5][5] + xor_out[99][5][5];

assign sum_out[0][5][6] = xor_out[0][5][6] + xor_out[1][5][6] + xor_out[2][5][6] + xor_out[3][5][6] + xor_out[4][5][6];
assign sum_out[1][5][6] = xor_out[5][5][6] + xor_out[6][5][6] + xor_out[7][5][6] + xor_out[8][5][6] + xor_out[9][5][6];
assign sum_out[2][5][6] = xor_out[10][5][6] + xor_out[11][5][6] + xor_out[12][5][6] + xor_out[13][5][6] + xor_out[14][5][6];
assign sum_out[3][5][6] = xor_out[15][5][6] + xor_out[16][5][6] + xor_out[17][5][6] + xor_out[18][5][6] + xor_out[19][5][6];
assign sum_out[4][5][6] = xor_out[20][5][6] + xor_out[21][5][6] + xor_out[22][5][6] + xor_out[23][5][6] + xor_out[24][5][6];
assign sum_out[5][5][6] = xor_out[25][5][6] + xor_out[26][5][6] + xor_out[27][5][6] + xor_out[28][5][6] + xor_out[29][5][6];
assign sum_out[6][5][6] = xor_out[30][5][6] + xor_out[31][5][6] + xor_out[32][5][6] + xor_out[33][5][6] + xor_out[34][5][6];
assign sum_out[7][5][6] = xor_out[35][5][6] + xor_out[36][5][6] + xor_out[37][5][6] + xor_out[38][5][6] + xor_out[39][5][6];
assign sum_out[8][5][6] = xor_out[40][5][6] + xor_out[41][5][6] + xor_out[42][5][6] + xor_out[43][5][6] + xor_out[44][5][6];
assign sum_out[9][5][6] = xor_out[45][5][6] + xor_out[46][5][6] + xor_out[47][5][6] + xor_out[48][5][6] + xor_out[49][5][6];
assign sum_out[10][5][6] = xor_out[50][5][6] + xor_out[51][5][6] + xor_out[52][5][6] + xor_out[53][5][6] + xor_out[54][5][6];
assign sum_out[11][5][6] = xor_out[55][5][6] + xor_out[56][5][6] + xor_out[57][5][6] + xor_out[58][5][6] + xor_out[59][5][6];
assign sum_out[12][5][6] = xor_out[60][5][6] + xor_out[61][5][6] + xor_out[62][5][6] + xor_out[63][5][6] + xor_out[64][5][6];
assign sum_out[13][5][6] = xor_out[65][5][6] + xor_out[66][5][6] + xor_out[67][5][6] + xor_out[68][5][6] + xor_out[69][5][6];
assign sum_out[14][5][6] = xor_out[70][5][6] + xor_out[71][5][6] + xor_out[72][5][6] + xor_out[73][5][6] + xor_out[74][5][6];
assign sum_out[15][5][6] = xor_out[75][5][6] + xor_out[76][5][6] + xor_out[77][5][6] + xor_out[78][5][6] + xor_out[79][5][6];
assign sum_out[16][5][6] = xor_out[80][5][6] + xor_out[81][5][6] + xor_out[82][5][6] + xor_out[83][5][6] + xor_out[84][5][6];
assign sum_out[17][5][6] = xor_out[85][5][6] + xor_out[86][5][6] + xor_out[87][5][6] + xor_out[88][5][6] + xor_out[89][5][6];
assign sum_out[18][5][6] = xor_out[90][5][6] + xor_out[91][5][6] + xor_out[92][5][6] + xor_out[93][5][6] + xor_out[94][5][6];
assign sum_out[19][5][6] = xor_out[95][5][6] + xor_out[96][5][6] + xor_out[97][5][6] + xor_out[98][5][6] + xor_out[99][5][6];

assign sum_out[0][5][7] = xor_out[0][5][7] + xor_out[1][5][7] + xor_out[2][5][7] + xor_out[3][5][7] + xor_out[4][5][7];
assign sum_out[1][5][7] = xor_out[5][5][7] + xor_out[6][5][7] + xor_out[7][5][7] + xor_out[8][5][7] + xor_out[9][5][7];
assign sum_out[2][5][7] = xor_out[10][5][7] + xor_out[11][5][7] + xor_out[12][5][7] + xor_out[13][5][7] + xor_out[14][5][7];
assign sum_out[3][5][7] = xor_out[15][5][7] + xor_out[16][5][7] + xor_out[17][5][7] + xor_out[18][5][7] + xor_out[19][5][7];
assign sum_out[4][5][7] = xor_out[20][5][7] + xor_out[21][5][7] + xor_out[22][5][7] + xor_out[23][5][7] + xor_out[24][5][7];
assign sum_out[5][5][7] = xor_out[25][5][7] + xor_out[26][5][7] + xor_out[27][5][7] + xor_out[28][5][7] + xor_out[29][5][7];
assign sum_out[6][5][7] = xor_out[30][5][7] + xor_out[31][5][7] + xor_out[32][5][7] + xor_out[33][5][7] + xor_out[34][5][7];
assign sum_out[7][5][7] = xor_out[35][5][7] + xor_out[36][5][7] + xor_out[37][5][7] + xor_out[38][5][7] + xor_out[39][5][7];
assign sum_out[8][5][7] = xor_out[40][5][7] + xor_out[41][5][7] + xor_out[42][5][7] + xor_out[43][5][7] + xor_out[44][5][7];
assign sum_out[9][5][7] = xor_out[45][5][7] + xor_out[46][5][7] + xor_out[47][5][7] + xor_out[48][5][7] + xor_out[49][5][7];
assign sum_out[10][5][7] = xor_out[50][5][7] + xor_out[51][5][7] + xor_out[52][5][7] + xor_out[53][5][7] + xor_out[54][5][7];
assign sum_out[11][5][7] = xor_out[55][5][7] + xor_out[56][5][7] + xor_out[57][5][7] + xor_out[58][5][7] + xor_out[59][5][7];
assign sum_out[12][5][7] = xor_out[60][5][7] + xor_out[61][5][7] + xor_out[62][5][7] + xor_out[63][5][7] + xor_out[64][5][7];
assign sum_out[13][5][7] = xor_out[65][5][7] + xor_out[66][5][7] + xor_out[67][5][7] + xor_out[68][5][7] + xor_out[69][5][7];
assign sum_out[14][5][7] = xor_out[70][5][7] + xor_out[71][5][7] + xor_out[72][5][7] + xor_out[73][5][7] + xor_out[74][5][7];
assign sum_out[15][5][7] = xor_out[75][5][7] + xor_out[76][5][7] + xor_out[77][5][7] + xor_out[78][5][7] + xor_out[79][5][7];
assign sum_out[16][5][7] = xor_out[80][5][7] + xor_out[81][5][7] + xor_out[82][5][7] + xor_out[83][5][7] + xor_out[84][5][7];
assign sum_out[17][5][7] = xor_out[85][5][7] + xor_out[86][5][7] + xor_out[87][5][7] + xor_out[88][5][7] + xor_out[89][5][7];
assign sum_out[18][5][7] = xor_out[90][5][7] + xor_out[91][5][7] + xor_out[92][5][7] + xor_out[93][5][7] + xor_out[94][5][7];
assign sum_out[19][5][7] = xor_out[95][5][7] + xor_out[96][5][7] + xor_out[97][5][7] + xor_out[98][5][7] + xor_out[99][5][7];

assign sum_out[0][5][8] = xor_out[0][5][8] + xor_out[1][5][8] + xor_out[2][5][8] + xor_out[3][5][8] + xor_out[4][5][8];
assign sum_out[1][5][8] = xor_out[5][5][8] + xor_out[6][5][8] + xor_out[7][5][8] + xor_out[8][5][8] + xor_out[9][5][8];
assign sum_out[2][5][8] = xor_out[10][5][8] + xor_out[11][5][8] + xor_out[12][5][8] + xor_out[13][5][8] + xor_out[14][5][8];
assign sum_out[3][5][8] = xor_out[15][5][8] + xor_out[16][5][8] + xor_out[17][5][8] + xor_out[18][5][8] + xor_out[19][5][8];
assign sum_out[4][5][8] = xor_out[20][5][8] + xor_out[21][5][8] + xor_out[22][5][8] + xor_out[23][5][8] + xor_out[24][5][8];
assign sum_out[5][5][8] = xor_out[25][5][8] + xor_out[26][5][8] + xor_out[27][5][8] + xor_out[28][5][8] + xor_out[29][5][8];
assign sum_out[6][5][8] = xor_out[30][5][8] + xor_out[31][5][8] + xor_out[32][5][8] + xor_out[33][5][8] + xor_out[34][5][8];
assign sum_out[7][5][8] = xor_out[35][5][8] + xor_out[36][5][8] + xor_out[37][5][8] + xor_out[38][5][8] + xor_out[39][5][8];
assign sum_out[8][5][8] = xor_out[40][5][8] + xor_out[41][5][8] + xor_out[42][5][8] + xor_out[43][5][8] + xor_out[44][5][8];
assign sum_out[9][5][8] = xor_out[45][5][8] + xor_out[46][5][8] + xor_out[47][5][8] + xor_out[48][5][8] + xor_out[49][5][8];
assign sum_out[10][5][8] = xor_out[50][5][8] + xor_out[51][5][8] + xor_out[52][5][8] + xor_out[53][5][8] + xor_out[54][5][8];
assign sum_out[11][5][8] = xor_out[55][5][8] + xor_out[56][5][8] + xor_out[57][5][8] + xor_out[58][5][8] + xor_out[59][5][8];
assign sum_out[12][5][8] = xor_out[60][5][8] + xor_out[61][5][8] + xor_out[62][5][8] + xor_out[63][5][8] + xor_out[64][5][8];
assign sum_out[13][5][8] = xor_out[65][5][8] + xor_out[66][5][8] + xor_out[67][5][8] + xor_out[68][5][8] + xor_out[69][5][8];
assign sum_out[14][5][8] = xor_out[70][5][8] + xor_out[71][5][8] + xor_out[72][5][8] + xor_out[73][5][8] + xor_out[74][5][8];
assign sum_out[15][5][8] = xor_out[75][5][8] + xor_out[76][5][8] + xor_out[77][5][8] + xor_out[78][5][8] + xor_out[79][5][8];
assign sum_out[16][5][8] = xor_out[80][5][8] + xor_out[81][5][8] + xor_out[82][5][8] + xor_out[83][5][8] + xor_out[84][5][8];
assign sum_out[17][5][8] = xor_out[85][5][8] + xor_out[86][5][8] + xor_out[87][5][8] + xor_out[88][5][8] + xor_out[89][5][8];
assign sum_out[18][5][8] = xor_out[90][5][8] + xor_out[91][5][8] + xor_out[92][5][8] + xor_out[93][5][8] + xor_out[94][5][8];
assign sum_out[19][5][8] = xor_out[95][5][8] + xor_out[96][5][8] + xor_out[97][5][8] + xor_out[98][5][8] + xor_out[99][5][8];

assign sum_out[0][5][9] = xor_out[0][5][9] + xor_out[1][5][9] + xor_out[2][5][9] + xor_out[3][5][9] + xor_out[4][5][9];
assign sum_out[1][5][9] = xor_out[5][5][9] + xor_out[6][5][9] + xor_out[7][5][9] + xor_out[8][5][9] + xor_out[9][5][9];
assign sum_out[2][5][9] = xor_out[10][5][9] + xor_out[11][5][9] + xor_out[12][5][9] + xor_out[13][5][9] + xor_out[14][5][9];
assign sum_out[3][5][9] = xor_out[15][5][9] + xor_out[16][5][9] + xor_out[17][5][9] + xor_out[18][5][9] + xor_out[19][5][9];
assign sum_out[4][5][9] = xor_out[20][5][9] + xor_out[21][5][9] + xor_out[22][5][9] + xor_out[23][5][9] + xor_out[24][5][9];
assign sum_out[5][5][9] = xor_out[25][5][9] + xor_out[26][5][9] + xor_out[27][5][9] + xor_out[28][5][9] + xor_out[29][5][9];
assign sum_out[6][5][9] = xor_out[30][5][9] + xor_out[31][5][9] + xor_out[32][5][9] + xor_out[33][5][9] + xor_out[34][5][9];
assign sum_out[7][5][9] = xor_out[35][5][9] + xor_out[36][5][9] + xor_out[37][5][9] + xor_out[38][5][9] + xor_out[39][5][9];
assign sum_out[8][5][9] = xor_out[40][5][9] + xor_out[41][5][9] + xor_out[42][5][9] + xor_out[43][5][9] + xor_out[44][5][9];
assign sum_out[9][5][9] = xor_out[45][5][9] + xor_out[46][5][9] + xor_out[47][5][9] + xor_out[48][5][9] + xor_out[49][5][9];
assign sum_out[10][5][9] = xor_out[50][5][9] + xor_out[51][5][9] + xor_out[52][5][9] + xor_out[53][5][9] + xor_out[54][5][9];
assign sum_out[11][5][9] = xor_out[55][5][9] + xor_out[56][5][9] + xor_out[57][5][9] + xor_out[58][5][9] + xor_out[59][5][9];
assign sum_out[12][5][9] = xor_out[60][5][9] + xor_out[61][5][9] + xor_out[62][5][9] + xor_out[63][5][9] + xor_out[64][5][9];
assign sum_out[13][5][9] = xor_out[65][5][9] + xor_out[66][5][9] + xor_out[67][5][9] + xor_out[68][5][9] + xor_out[69][5][9];
assign sum_out[14][5][9] = xor_out[70][5][9] + xor_out[71][5][9] + xor_out[72][5][9] + xor_out[73][5][9] + xor_out[74][5][9];
assign sum_out[15][5][9] = xor_out[75][5][9] + xor_out[76][5][9] + xor_out[77][5][9] + xor_out[78][5][9] + xor_out[79][5][9];
assign sum_out[16][5][9] = xor_out[80][5][9] + xor_out[81][5][9] + xor_out[82][5][9] + xor_out[83][5][9] + xor_out[84][5][9];
assign sum_out[17][5][9] = xor_out[85][5][9] + xor_out[86][5][9] + xor_out[87][5][9] + xor_out[88][5][9] + xor_out[89][5][9];
assign sum_out[18][5][9] = xor_out[90][5][9] + xor_out[91][5][9] + xor_out[92][5][9] + xor_out[93][5][9] + xor_out[94][5][9];
assign sum_out[19][5][9] = xor_out[95][5][9] + xor_out[96][5][9] + xor_out[97][5][9] + xor_out[98][5][9] + xor_out[99][5][9];

assign sum_out[0][5][10] = xor_out[0][5][10] + xor_out[1][5][10] + xor_out[2][5][10] + xor_out[3][5][10] + xor_out[4][5][10];
assign sum_out[1][5][10] = xor_out[5][5][10] + xor_out[6][5][10] + xor_out[7][5][10] + xor_out[8][5][10] + xor_out[9][5][10];
assign sum_out[2][5][10] = xor_out[10][5][10] + xor_out[11][5][10] + xor_out[12][5][10] + xor_out[13][5][10] + xor_out[14][5][10];
assign sum_out[3][5][10] = xor_out[15][5][10] + xor_out[16][5][10] + xor_out[17][5][10] + xor_out[18][5][10] + xor_out[19][5][10];
assign sum_out[4][5][10] = xor_out[20][5][10] + xor_out[21][5][10] + xor_out[22][5][10] + xor_out[23][5][10] + xor_out[24][5][10];
assign sum_out[5][5][10] = xor_out[25][5][10] + xor_out[26][5][10] + xor_out[27][5][10] + xor_out[28][5][10] + xor_out[29][5][10];
assign sum_out[6][5][10] = xor_out[30][5][10] + xor_out[31][5][10] + xor_out[32][5][10] + xor_out[33][5][10] + xor_out[34][5][10];
assign sum_out[7][5][10] = xor_out[35][5][10] + xor_out[36][5][10] + xor_out[37][5][10] + xor_out[38][5][10] + xor_out[39][5][10];
assign sum_out[8][5][10] = xor_out[40][5][10] + xor_out[41][5][10] + xor_out[42][5][10] + xor_out[43][5][10] + xor_out[44][5][10];
assign sum_out[9][5][10] = xor_out[45][5][10] + xor_out[46][5][10] + xor_out[47][5][10] + xor_out[48][5][10] + xor_out[49][5][10];
assign sum_out[10][5][10] = xor_out[50][5][10] + xor_out[51][5][10] + xor_out[52][5][10] + xor_out[53][5][10] + xor_out[54][5][10];
assign sum_out[11][5][10] = xor_out[55][5][10] + xor_out[56][5][10] + xor_out[57][5][10] + xor_out[58][5][10] + xor_out[59][5][10];
assign sum_out[12][5][10] = xor_out[60][5][10] + xor_out[61][5][10] + xor_out[62][5][10] + xor_out[63][5][10] + xor_out[64][5][10];
assign sum_out[13][5][10] = xor_out[65][5][10] + xor_out[66][5][10] + xor_out[67][5][10] + xor_out[68][5][10] + xor_out[69][5][10];
assign sum_out[14][5][10] = xor_out[70][5][10] + xor_out[71][5][10] + xor_out[72][5][10] + xor_out[73][5][10] + xor_out[74][5][10];
assign sum_out[15][5][10] = xor_out[75][5][10] + xor_out[76][5][10] + xor_out[77][5][10] + xor_out[78][5][10] + xor_out[79][5][10];
assign sum_out[16][5][10] = xor_out[80][5][10] + xor_out[81][5][10] + xor_out[82][5][10] + xor_out[83][5][10] + xor_out[84][5][10];
assign sum_out[17][5][10] = xor_out[85][5][10] + xor_out[86][5][10] + xor_out[87][5][10] + xor_out[88][5][10] + xor_out[89][5][10];
assign sum_out[18][5][10] = xor_out[90][5][10] + xor_out[91][5][10] + xor_out[92][5][10] + xor_out[93][5][10] + xor_out[94][5][10];
assign sum_out[19][5][10] = xor_out[95][5][10] + xor_out[96][5][10] + xor_out[97][5][10] + xor_out[98][5][10] + xor_out[99][5][10];

assign sum_out[0][5][11] = xor_out[0][5][11] + xor_out[1][5][11] + xor_out[2][5][11] + xor_out[3][5][11] + xor_out[4][5][11];
assign sum_out[1][5][11] = xor_out[5][5][11] + xor_out[6][5][11] + xor_out[7][5][11] + xor_out[8][5][11] + xor_out[9][5][11];
assign sum_out[2][5][11] = xor_out[10][5][11] + xor_out[11][5][11] + xor_out[12][5][11] + xor_out[13][5][11] + xor_out[14][5][11];
assign sum_out[3][5][11] = xor_out[15][5][11] + xor_out[16][5][11] + xor_out[17][5][11] + xor_out[18][5][11] + xor_out[19][5][11];
assign sum_out[4][5][11] = xor_out[20][5][11] + xor_out[21][5][11] + xor_out[22][5][11] + xor_out[23][5][11] + xor_out[24][5][11];
assign sum_out[5][5][11] = xor_out[25][5][11] + xor_out[26][5][11] + xor_out[27][5][11] + xor_out[28][5][11] + xor_out[29][5][11];
assign sum_out[6][5][11] = xor_out[30][5][11] + xor_out[31][5][11] + xor_out[32][5][11] + xor_out[33][5][11] + xor_out[34][5][11];
assign sum_out[7][5][11] = xor_out[35][5][11] + xor_out[36][5][11] + xor_out[37][5][11] + xor_out[38][5][11] + xor_out[39][5][11];
assign sum_out[8][5][11] = xor_out[40][5][11] + xor_out[41][5][11] + xor_out[42][5][11] + xor_out[43][5][11] + xor_out[44][5][11];
assign sum_out[9][5][11] = xor_out[45][5][11] + xor_out[46][5][11] + xor_out[47][5][11] + xor_out[48][5][11] + xor_out[49][5][11];
assign sum_out[10][5][11] = xor_out[50][5][11] + xor_out[51][5][11] + xor_out[52][5][11] + xor_out[53][5][11] + xor_out[54][5][11];
assign sum_out[11][5][11] = xor_out[55][5][11] + xor_out[56][5][11] + xor_out[57][5][11] + xor_out[58][5][11] + xor_out[59][5][11];
assign sum_out[12][5][11] = xor_out[60][5][11] + xor_out[61][5][11] + xor_out[62][5][11] + xor_out[63][5][11] + xor_out[64][5][11];
assign sum_out[13][5][11] = xor_out[65][5][11] + xor_out[66][5][11] + xor_out[67][5][11] + xor_out[68][5][11] + xor_out[69][5][11];
assign sum_out[14][5][11] = xor_out[70][5][11] + xor_out[71][5][11] + xor_out[72][5][11] + xor_out[73][5][11] + xor_out[74][5][11];
assign sum_out[15][5][11] = xor_out[75][5][11] + xor_out[76][5][11] + xor_out[77][5][11] + xor_out[78][5][11] + xor_out[79][5][11];
assign sum_out[16][5][11] = xor_out[80][5][11] + xor_out[81][5][11] + xor_out[82][5][11] + xor_out[83][5][11] + xor_out[84][5][11];
assign sum_out[17][5][11] = xor_out[85][5][11] + xor_out[86][5][11] + xor_out[87][5][11] + xor_out[88][5][11] + xor_out[89][5][11];
assign sum_out[18][5][11] = xor_out[90][5][11] + xor_out[91][5][11] + xor_out[92][5][11] + xor_out[93][5][11] + xor_out[94][5][11];
assign sum_out[19][5][11] = xor_out[95][5][11] + xor_out[96][5][11] + xor_out[97][5][11] + xor_out[98][5][11] + xor_out[99][5][11];

assign sum_out[0][5][12] = xor_out[0][5][12] + xor_out[1][5][12] + xor_out[2][5][12] + xor_out[3][5][12] + xor_out[4][5][12];
assign sum_out[1][5][12] = xor_out[5][5][12] + xor_out[6][5][12] + xor_out[7][5][12] + xor_out[8][5][12] + xor_out[9][5][12];
assign sum_out[2][5][12] = xor_out[10][5][12] + xor_out[11][5][12] + xor_out[12][5][12] + xor_out[13][5][12] + xor_out[14][5][12];
assign sum_out[3][5][12] = xor_out[15][5][12] + xor_out[16][5][12] + xor_out[17][5][12] + xor_out[18][5][12] + xor_out[19][5][12];
assign sum_out[4][5][12] = xor_out[20][5][12] + xor_out[21][5][12] + xor_out[22][5][12] + xor_out[23][5][12] + xor_out[24][5][12];
assign sum_out[5][5][12] = xor_out[25][5][12] + xor_out[26][5][12] + xor_out[27][5][12] + xor_out[28][5][12] + xor_out[29][5][12];
assign sum_out[6][5][12] = xor_out[30][5][12] + xor_out[31][5][12] + xor_out[32][5][12] + xor_out[33][5][12] + xor_out[34][5][12];
assign sum_out[7][5][12] = xor_out[35][5][12] + xor_out[36][5][12] + xor_out[37][5][12] + xor_out[38][5][12] + xor_out[39][5][12];
assign sum_out[8][5][12] = xor_out[40][5][12] + xor_out[41][5][12] + xor_out[42][5][12] + xor_out[43][5][12] + xor_out[44][5][12];
assign sum_out[9][5][12] = xor_out[45][5][12] + xor_out[46][5][12] + xor_out[47][5][12] + xor_out[48][5][12] + xor_out[49][5][12];
assign sum_out[10][5][12] = xor_out[50][5][12] + xor_out[51][5][12] + xor_out[52][5][12] + xor_out[53][5][12] + xor_out[54][5][12];
assign sum_out[11][5][12] = xor_out[55][5][12] + xor_out[56][5][12] + xor_out[57][5][12] + xor_out[58][5][12] + xor_out[59][5][12];
assign sum_out[12][5][12] = xor_out[60][5][12] + xor_out[61][5][12] + xor_out[62][5][12] + xor_out[63][5][12] + xor_out[64][5][12];
assign sum_out[13][5][12] = xor_out[65][5][12] + xor_out[66][5][12] + xor_out[67][5][12] + xor_out[68][5][12] + xor_out[69][5][12];
assign sum_out[14][5][12] = xor_out[70][5][12] + xor_out[71][5][12] + xor_out[72][5][12] + xor_out[73][5][12] + xor_out[74][5][12];
assign sum_out[15][5][12] = xor_out[75][5][12] + xor_out[76][5][12] + xor_out[77][5][12] + xor_out[78][5][12] + xor_out[79][5][12];
assign sum_out[16][5][12] = xor_out[80][5][12] + xor_out[81][5][12] + xor_out[82][5][12] + xor_out[83][5][12] + xor_out[84][5][12];
assign sum_out[17][5][12] = xor_out[85][5][12] + xor_out[86][5][12] + xor_out[87][5][12] + xor_out[88][5][12] + xor_out[89][5][12];
assign sum_out[18][5][12] = xor_out[90][5][12] + xor_out[91][5][12] + xor_out[92][5][12] + xor_out[93][5][12] + xor_out[94][5][12];
assign sum_out[19][5][12] = xor_out[95][5][12] + xor_out[96][5][12] + xor_out[97][5][12] + xor_out[98][5][12] + xor_out[99][5][12];

assign sum_out[0][5][13] = xor_out[0][5][13] + xor_out[1][5][13] + xor_out[2][5][13] + xor_out[3][5][13] + xor_out[4][5][13];
assign sum_out[1][5][13] = xor_out[5][5][13] + xor_out[6][5][13] + xor_out[7][5][13] + xor_out[8][5][13] + xor_out[9][5][13];
assign sum_out[2][5][13] = xor_out[10][5][13] + xor_out[11][5][13] + xor_out[12][5][13] + xor_out[13][5][13] + xor_out[14][5][13];
assign sum_out[3][5][13] = xor_out[15][5][13] + xor_out[16][5][13] + xor_out[17][5][13] + xor_out[18][5][13] + xor_out[19][5][13];
assign sum_out[4][5][13] = xor_out[20][5][13] + xor_out[21][5][13] + xor_out[22][5][13] + xor_out[23][5][13] + xor_out[24][5][13];
assign sum_out[5][5][13] = xor_out[25][5][13] + xor_out[26][5][13] + xor_out[27][5][13] + xor_out[28][5][13] + xor_out[29][5][13];
assign sum_out[6][5][13] = xor_out[30][5][13] + xor_out[31][5][13] + xor_out[32][5][13] + xor_out[33][5][13] + xor_out[34][5][13];
assign sum_out[7][5][13] = xor_out[35][5][13] + xor_out[36][5][13] + xor_out[37][5][13] + xor_out[38][5][13] + xor_out[39][5][13];
assign sum_out[8][5][13] = xor_out[40][5][13] + xor_out[41][5][13] + xor_out[42][5][13] + xor_out[43][5][13] + xor_out[44][5][13];
assign sum_out[9][5][13] = xor_out[45][5][13] + xor_out[46][5][13] + xor_out[47][5][13] + xor_out[48][5][13] + xor_out[49][5][13];
assign sum_out[10][5][13] = xor_out[50][5][13] + xor_out[51][5][13] + xor_out[52][5][13] + xor_out[53][5][13] + xor_out[54][5][13];
assign sum_out[11][5][13] = xor_out[55][5][13] + xor_out[56][5][13] + xor_out[57][5][13] + xor_out[58][5][13] + xor_out[59][5][13];
assign sum_out[12][5][13] = xor_out[60][5][13] + xor_out[61][5][13] + xor_out[62][5][13] + xor_out[63][5][13] + xor_out[64][5][13];
assign sum_out[13][5][13] = xor_out[65][5][13] + xor_out[66][5][13] + xor_out[67][5][13] + xor_out[68][5][13] + xor_out[69][5][13];
assign sum_out[14][5][13] = xor_out[70][5][13] + xor_out[71][5][13] + xor_out[72][5][13] + xor_out[73][5][13] + xor_out[74][5][13];
assign sum_out[15][5][13] = xor_out[75][5][13] + xor_out[76][5][13] + xor_out[77][5][13] + xor_out[78][5][13] + xor_out[79][5][13];
assign sum_out[16][5][13] = xor_out[80][5][13] + xor_out[81][5][13] + xor_out[82][5][13] + xor_out[83][5][13] + xor_out[84][5][13];
assign sum_out[17][5][13] = xor_out[85][5][13] + xor_out[86][5][13] + xor_out[87][5][13] + xor_out[88][5][13] + xor_out[89][5][13];
assign sum_out[18][5][13] = xor_out[90][5][13] + xor_out[91][5][13] + xor_out[92][5][13] + xor_out[93][5][13] + xor_out[94][5][13];
assign sum_out[19][5][13] = xor_out[95][5][13] + xor_out[96][5][13] + xor_out[97][5][13] + xor_out[98][5][13] + xor_out[99][5][13];

assign sum_out[0][5][14] = xor_out[0][5][14] + xor_out[1][5][14] + xor_out[2][5][14] + xor_out[3][5][14] + xor_out[4][5][14];
assign sum_out[1][5][14] = xor_out[5][5][14] + xor_out[6][5][14] + xor_out[7][5][14] + xor_out[8][5][14] + xor_out[9][5][14];
assign sum_out[2][5][14] = xor_out[10][5][14] + xor_out[11][5][14] + xor_out[12][5][14] + xor_out[13][5][14] + xor_out[14][5][14];
assign sum_out[3][5][14] = xor_out[15][5][14] + xor_out[16][5][14] + xor_out[17][5][14] + xor_out[18][5][14] + xor_out[19][5][14];
assign sum_out[4][5][14] = xor_out[20][5][14] + xor_out[21][5][14] + xor_out[22][5][14] + xor_out[23][5][14] + xor_out[24][5][14];
assign sum_out[5][5][14] = xor_out[25][5][14] + xor_out[26][5][14] + xor_out[27][5][14] + xor_out[28][5][14] + xor_out[29][5][14];
assign sum_out[6][5][14] = xor_out[30][5][14] + xor_out[31][5][14] + xor_out[32][5][14] + xor_out[33][5][14] + xor_out[34][5][14];
assign sum_out[7][5][14] = xor_out[35][5][14] + xor_out[36][5][14] + xor_out[37][5][14] + xor_out[38][5][14] + xor_out[39][5][14];
assign sum_out[8][5][14] = xor_out[40][5][14] + xor_out[41][5][14] + xor_out[42][5][14] + xor_out[43][5][14] + xor_out[44][5][14];
assign sum_out[9][5][14] = xor_out[45][5][14] + xor_out[46][5][14] + xor_out[47][5][14] + xor_out[48][5][14] + xor_out[49][5][14];
assign sum_out[10][5][14] = xor_out[50][5][14] + xor_out[51][5][14] + xor_out[52][5][14] + xor_out[53][5][14] + xor_out[54][5][14];
assign sum_out[11][5][14] = xor_out[55][5][14] + xor_out[56][5][14] + xor_out[57][5][14] + xor_out[58][5][14] + xor_out[59][5][14];
assign sum_out[12][5][14] = xor_out[60][5][14] + xor_out[61][5][14] + xor_out[62][5][14] + xor_out[63][5][14] + xor_out[64][5][14];
assign sum_out[13][5][14] = xor_out[65][5][14] + xor_out[66][5][14] + xor_out[67][5][14] + xor_out[68][5][14] + xor_out[69][5][14];
assign sum_out[14][5][14] = xor_out[70][5][14] + xor_out[71][5][14] + xor_out[72][5][14] + xor_out[73][5][14] + xor_out[74][5][14];
assign sum_out[15][5][14] = xor_out[75][5][14] + xor_out[76][5][14] + xor_out[77][5][14] + xor_out[78][5][14] + xor_out[79][5][14];
assign sum_out[16][5][14] = xor_out[80][5][14] + xor_out[81][5][14] + xor_out[82][5][14] + xor_out[83][5][14] + xor_out[84][5][14];
assign sum_out[17][5][14] = xor_out[85][5][14] + xor_out[86][5][14] + xor_out[87][5][14] + xor_out[88][5][14] + xor_out[89][5][14];
assign sum_out[18][5][14] = xor_out[90][5][14] + xor_out[91][5][14] + xor_out[92][5][14] + xor_out[93][5][14] + xor_out[94][5][14];
assign sum_out[19][5][14] = xor_out[95][5][14] + xor_out[96][5][14] + xor_out[97][5][14] + xor_out[98][5][14] + xor_out[99][5][14];

assign sum_out[0][5][15] = xor_out[0][5][15] + xor_out[1][5][15] + xor_out[2][5][15] + xor_out[3][5][15] + xor_out[4][5][15];
assign sum_out[1][5][15] = xor_out[5][5][15] + xor_out[6][5][15] + xor_out[7][5][15] + xor_out[8][5][15] + xor_out[9][5][15];
assign sum_out[2][5][15] = xor_out[10][5][15] + xor_out[11][5][15] + xor_out[12][5][15] + xor_out[13][5][15] + xor_out[14][5][15];
assign sum_out[3][5][15] = xor_out[15][5][15] + xor_out[16][5][15] + xor_out[17][5][15] + xor_out[18][5][15] + xor_out[19][5][15];
assign sum_out[4][5][15] = xor_out[20][5][15] + xor_out[21][5][15] + xor_out[22][5][15] + xor_out[23][5][15] + xor_out[24][5][15];
assign sum_out[5][5][15] = xor_out[25][5][15] + xor_out[26][5][15] + xor_out[27][5][15] + xor_out[28][5][15] + xor_out[29][5][15];
assign sum_out[6][5][15] = xor_out[30][5][15] + xor_out[31][5][15] + xor_out[32][5][15] + xor_out[33][5][15] + xor_out[34][5][15];
assign sum_out[7][5][15] = xor_out[35][5][15] + xor_out[36][5][15] + xor_out[37][5][15] + xor_out[38][5][15] + xor_out[39][5][15];
assign sum_out[8][5][15] = xor_out[40][5][15] + xor_out[41][5][15] + xor_out[42][5][15] + xor_out[43][5][15] + xor_out[44][5][15];
assign sum_out[9][5][15] = xor_out[45][5][15] + xor_out[46][5][15] + xor_out[47][5][15] + xor_out[48][5][15] + xor_out[49][5][15];
assign sum_out[10][5][15] = xor_out[50][5][15] + xor_out[51][5][15] + xor_out[52][5][15] + xor_out[53][5][15] + xor_out[54][5][15];
assign sum_out[11][5][15] = xor_out[55][5][15] + xor_out[56][5][15] + xor_out[57][5][15] + xor_out[58][5][15] + xor_out[59][5][15];
assign sum_out[12][5][15] = xor_out[60][5][15] + xor_out[61][5][15] + xor_out[62][5][15] + xor_out[63][5][15] + xor_out[64][5][15];
assign sum_out[13][5][15] = xor_out[65][5][15] + xor_out[66][5][15] + xor_out[67][5][15] + xor_out[68][5][15] + xor_out[69][5][15];
assign sum_out[14][5][15] = xor_out[70][5][15] + xor_out[71][5][15] + xor_out[72][5][15] + xor_out[73][5][15] + xor_out[74][5][15];
assign sum_out[15][5][15] = xor_out[75][5][15] + xor_out[76][5][15] + xor_out[77][5][15] + xor_out[78][5][15] + xor_out[79][5][15];
assign sum_out[16][5][15] = xor_out[80][5][15] + xor_out[81][5][15] + xor_out[82][5][15] + xor_out[83][5][15] + xor_out[84][5][15];
assign sum_out[17][5][15] = xor_out[85][5][15] + xor_out[86][5][15] + xor_out[87][5][15] + xor_out[88][5][15] + xor_out[89][5][15];
assign sum_out[18][5][15] = xor_out[90][5][15] + xor_out[91][5][15] + xor_out[92][5][15] + xor_out[93][5][15] + xor_out[94][5][15];
assign sum_out[19][5][15] = xor_out[95][5][15] + xor_out[96][5][15] + xor_out[97][5][15] + xor_out[98][5][15] + xor_out[99][5][15];

assign sum_out[0][5][16] = xor_out[0][5][16] + xor_out[1][5][16] + xor_out[2][5][16] + xor_out[3][5][16] + xor_out[4][5][16];
assign sum_out[1][5][16] = xor_out[5][5][16] + xor_out[6][5][16] + xor_out[7][5][16] + xor_out[8][5][16] + xor_out[9][5][16];
assign sum_out[2][5][16] = xor_out[10][5][16] + xor_out[11][5][16] + xor_out[12][5][16] + xor_out[13][5][16] + xor_out[14][5][16];
assign sum_out[3][5][16] = xor_out[15][5][16] + xor_out[16][5][16] + xor_out[17][5][16] + xor_out[18][5][16] + xor_out[19][5][16];
assign sum_out[4][5][16] = xor_out[20][5][16] + xor_out[21][5][16] + xor_out[22][5][16] + xor_out[23][5][16] + xor_out[24][5][16];
assign sum_out[5][5][16] = xor_out[25][5][16] + xor_out[26][5][16] + xor_out[27][5][16] + xor_out[28][5][16] + xor_out[29][5][16];
assign sum_out[6][5][16] = xor_out[30][5][16] + xor_out[31][5][16] + xor_out[32][5][16] + xor_out[33][5][16] + xor_out[34][5][16];
assign sum_out[7][5][16] = xor_out[35][5][16] + xor_out[36][5][16] + xor_out[37][5][16] + xor_out[38][5][16] + xor_out[39][5][16];
assign sum_out[8][5][16] = xor_out[40][5][16] + xor_out[41][5][16] + xor_out[42][5][16] + xor_out[43][5][16] + xor_out[44][5][16];
assign sum_out[9][5][16] = xor_out[45][5][16] + xor_out[46][5][16] + xor_out[47][5][16] + xor_out[48][5][16] + xor_out[49][5][16];
assign sum_out[10][5][16] = xor_out[50][5][16] + xor_out[51][5][16] + xor_out[52][5][16] + xor_out[53][5][16] + xor_out[54][5][16];
assign sum_out[11][5][16] = xor_out[55][5][16] + xor_out[56][5][16] + xor_out[57][5][16] + xor_out[58][5][16] + xor_out[59][5][16];
assign sum_out[12][5][16] = xor_out[60][5][16] + xor_out[61][5][16] + xor_out[62][5][16] + xor_out[63][5][16] + xor_out[64][5][16];
assign sum_out[13][5][16] = xor_out[65][5][16] + xor_out[66][5][16] + xor_out[67][5][16] + xor_out[68][5][16] + xor_out[69][5][16];
assign sum_out[14][5][16] = xor_out[70][5][16] + xor_out[71][5][16] + xor_out[72][5][16] + xor_out[73][5][16] + xor_out[74][5][16];
assign sum_out[15][5][16] = xor_out[75][5][16] + xor_out[76][5][16] + xor_out[77][5][16] + xor_out[78][5][16] + xor_out[79][5][16];
assign sum_out[16][5][16] = xor_out[80][5][16] + xor_out[81][5][16] + xor_out[82][5][16] + xor_out[83][5][16] + xor_out[84][5][16];
assign sum_out[17][5][16] = xor_out[85][5][16] + xor_out[86][5][16] + xor_out[87][5][16] + xor_out[88][5][16] + xor_out[89][5][16];
assign sum_out[18][5][16] = xor_out[90][5][16] + xor_out[91][5][16] + xor_out[92][5][16] + xor_out[93][5][16] + xor_out[94][5][16];
assign sum_out[19][5][16] = xor_out[95][5][16] + xor_out[96][5][16] + xor_out[97][5][16] + xor_out[98][5][16] + xor_out[99][5][16];

assign sum_out[0][5][17] = xor_out[0][5][17] + xor_out[1][5][17] + xor_out[2][5][17] + xor_out[3][5][17] + xor_out[4][5][17];
assign sum_out[1][5][17] = xor_out[5][5][17] + xor_out[6][5][17] + xor_out[7][5][17] + xor_out[8][5][17] + xor_out[9][5][17];
assign sum_out[2][5][17] = xor_out[10][5][17] + xor_out[11][5][17] + xor_out[12][5][17] + xor_out[13][5][17] + xor_out[14][5][17];
assign sum_out[3][5][17] = xor_out[15][5][17] + xor_out[16][5][17] + xor_out[17][5][17] + xor_out[18][5][17] + xor_out[19][5][17];
assign sum_out[4][5][17] = xor_out[20][5][17] + xor_out[21][5][17] + xor_out[22][5][17] + xor_out[23][5][17] + xor_out[24][5][17];
assign sum_out[5][5][17] = xor_out[25][5][17] + xor_out[26][5][17] + xor_out[27][5][17] + xor_out[28][5][17] + xor_out[29][5][17];
assign sum_out[6][5][17] = xor_out[30][5][17] + xor_out[31][5][17] + xor_out[32][5][17] + xor_out[33][5][17] + xor_out[34][5][17];
assign sum_out[7][5][17] = xor_out[35][5][17] + xor_out[36][5][17] + xor_out[37][5][17] + xor_out[38][5][17] + xor_out[39][5][17];
assign sum_out[8][5][17] = xor_out[40][5][17] + xor_out[41][5][17] + xor_out[42][5][17] + xor_out[43][5][17] + xor_out[44][5][17];
assign sum_out[9][5][17] = xor_out[45][5][17] + xor_out[46][5][17] + xor_out[47][5][17] + xor_out[48][5][17] + xor_out[49][5][17];
assign sum_out[10][5][17] = xor_out[50][5][17] + xor_out[51][5][17] + xor_out[52][5][17] + xor_out[53][5][17] + xor_out[54][5][17];
assign sum_out[11][5][17] = xor_out[55][5][17] + xor_out[56][5][17] + xor_out[57][5][17] + xor_out[58][5][17] + xor_out[59][5][17];
assign sum_out[12][5][17] = xor_out[60][5][17] + xor_out[61][5][17] + xor_out[62][5][17] + xor_out[63][5][17] + xor_out[64][5][17];
assign sum_out[13][5][17] = xor_out[65][5][17] + xor_out[66][5][17] + xor_out[67][5][17] + xor_out[68][5][17] + xor_out[69][5][17];
assign sum_out[14][5][17] = xor_out[70][5][17] + xor_out[71][5][17] + xor_out[72][5][17] + xor_out[73][5][17] + xor_out[74][5][17];
assign sum_out[15][5][17] = xor_out[75][5][17] + xor_out[76][5][17] + xor_out[77][5][17] + xor_out[78][5][17] + xor_out[79][5][17];
assign sum_out[16][5][17] = xor_out[80][5][17] + xor_out[81][5][17] + xor_out[82][5][17] + xor_out[83][5][17] + xor_out[84][5][17];
assign sum_out[17][5][17] = xor_out[85][5][17] + xor_out[86][5][17] + xor_out[87][5][17] + xor_out[88][5][17] + xor_out[89][5][17];
assign sum_out[18][5][17] = xor_out[90][5][17] + xor_out[91][5][17] + xor_out[92][5][17] + xor_out[93][5][17] + xor_out[94][5][17];
assign sum_out[19][5][17] = xor_out[95][5][17] + xor_out[96][5][17] + xor_out[97][5][17] + xor_out[98][5][17] + xor_out[99][5][17];

assign sum_out[0][5][18] = xor_out[0][5][18] + xor_out[1][5][18] + xor_out[2][5][18] + xor_out[3][5][18] + xor_out[4][5][18];
assign sum_out[1][5][18] = xor_out[5][5][18] + xor_out[6][5][18] + xor_out[7][5][18] + xor_out[8][5][18] + xor_out[9][5][18];
assign sum_out[2][5][18] = xor_out[10][5][18] + xor_out[11][5][18] + xor_out[12][5][18] + xor_out[13][5][18] + xor_out[14][5][18];
assign sum_out[3][5][18] = xor_out[15][5][18] + xor_out[16][5][18] + xor_out[17][5][18] + xor_out[18][5][18] + xor_out[19][5][18];
assign sum_out[4][5][18] = xor_out[20][5][18] + xor_out[21][5][18] + xor_out[22][5][18] + xor_out[23][5][18] + xor_out[24][5][18];
assign sum_out[5][5][18] = xor_out[25][5][18] + xor_out[26][5][18] + xor_out[27][5][18] + xor_out[28][5][18] + xor_out[29][5][18];
assign sum_out[6][5][18] = xor_out[30][5][18] + xor_out[31][5][18] + xor_out[32][5][18] + xor_out[33][5][18] + xor_out[34][5][18];
assign sum_out[7][5][18] = xor_out[35][5][18] + xor_out[36][5][18] + xor_out[37][5][18] + xor_out[38][5][18] + xor_out[39][5][18];
assign sum_out[8][5][18] = xor_out[40][5][18] + xor_out[41][5][18] + xor_out[42][5][18] + xor_out[43][5][18] + xor_out[44][5][18];
assign sum_out[9][5][18] = xor_out[45][5][18] + xor_out[46][5][18] + xor_out[47][5][18] + xor_out[48][5][18] + xor_out[49][5][18];
assign sum_out[10][5][18] = xor_out[50][5][18] + xor_out[51][5][18] + xor_out[52][5][18] + xor_out[53][5][18] + xor_out[54][5][18];
assign sum_out[11][5][18] = xor_out[55][5][18] + xor_out[56][5][18] + xor_out[57][5][18] + xor_out[58][5][18] + xor_out[59][5][18];
assign sum_out[12][5][18] = xor_out[60][5][18] + xor_out[61][5][18] + xor_out[62][5][18] + xor_out[63][5][18] + xor_out[64][5][18];
assign sum_out[13][5][18] = xor_out[65][5][18] + xor_out[66][5][18] + xor_out[67][5][18] + xor_out[68][5][18] + xor_out[69][5][18];
assign sum_out[14][5][18] = xor_out[70][5][18] + xor_out[71][5][18] + xor_out[72][5][18] + xor_out[73][5][18] + xor_out[74][5][18];
assign sum_out[15][5][18] = xor_out[75][5][18] + xor_out[76][5][18] + xor_out[77][5][18] + xor_out[78][5][18] + xor_out[79][5][18];
assign sum_out[16][5][18] = xor_out[80][5][18] + xor_out[81][5][18] + xor_out[82][5][18] + xor_out[83][5][18] + xor_out[84][5][18];
assign sum_out[17][5][18] = xor_out[85][5][18] + xor_out[86][5][18] + xor_out[87][5][18] + xor_out[88][5][18] + xor_out[89][5][18];
assign sum_out[18][5][18] = xor_out[90][5][18] + xor_out[91][5][18] + xor_out[92][5][18] + xor_out[93][5][18] + xor_out[94][5][18];
assign sum_out[19][5][18] = xor_out[95][5][18] + xor_out[96][5][18] + xor_out[97][5][18] + xor_out[98][5][18] + xor_out[99][5][18];

assign sum_out[0][5][19] = xor_out[0][5][19] + xor_out[1][5][19] + xor_out[2][5][19] + xor_out[3][5][19] + xor_out[4][5][19];
assign sum_out[1][5][19] = xor_out[5][5][19] + xor_out[6][5][19] + xor_out[7][5][19] + xor_out[8][5][19] + xor_out[9][5][19];
assign sum_out[2][5][19] = xor_out[10][5][19] + xor_out[11][5][19] + xor_out[12][5][19] + xor_out[13][5][19] + xor_out[14][5][19];
assign sum_out[3][5][19] = xor_out[15][5][19] + xor_out[16][5][19] + xor_out[17][5][19] + xor_out[18][5][19] + xor_out[19][5][19];
assign sum_out[4][5][19] = xor_out[20][5][19] + xor_out[21][5][19] + xor_out[22][5][19] + xor_out[23][5][19] + xor_out[24][5][19];
assign sum_out[5][5][19] = xor_out[25][5][19] + xor_out[26][5][19] + xor_out[27][5][19] + xor_out[28][5][19] + xor_out[29][5][19];
assign sum_out[6][5][19] = xor_out[30][5][19] + xor_out[31][5][19] + xor_out[32][5][19] + xor_out[33][5][19] + xor_out[34][5][19];
assign sum_out[7][5][19] = xor_out[35][5][19] + xor_out[36][5][19] + xor_out[37][5][19] + xor_out[38][5][19] + xor_out[39][5][19];
assign sum_out[8][5][19] = xor_out[40][5][19] + xor_out[41][5][19] + xor_out[42][5][19] + xor_out[43][5][19] + xor_out[44][5][19];
assign sum_out[9][5][19] = xor_out[45][5][19] + xor_out[46][5][19] + xor_out[47][5][19] + xor_out[48][5][19] + xor_out[49][5][19];
assign sum_out[10][5][19] = xor_out[50][5][19] + xor_out[51][5][19] + xor_out[52][5][19] + xor_out[53][5][19] + xor_out[54][5][19];
assign sum_out[11][5][19] = xor_out[55][5][19] + xor_out[56][5][19] + xor_out[57][5][19] + xor_out[58][5][19] + xor_out[59][5][19];
assign sum_out[12][5][19] = xor_out[60][5][19] + xor_out[61][5][19] + xor_out[62][5][19] + xor_out[63][5][19] + xor_out[64][5][19];
assign sum_out[13][5][19] = xor_out[65][5][19] + xor_out[66][5][19] + xor_out[67][5][19] + xor_out[68][5][19] + xor_out[69][5][19];
assign sum_out[14][5][19] = xor_out[70][5][19] + xor_out[71][5][19] + xor_out[72][5][19] + xor_out[73][5][19] + xor_out[74][5][19];
assign sum_out[15][5][19] = xor_out[75][5][19] + xor_out[76][5][19] + xor_out[77][5][19] + xor_out[78][5][19] + xor_out[79][5][19];
assign sum_out[16][5][19] = xor_out[80][5][19] + xor_out[81][5][19] + xor_out[82][5][19] + xor_out[83][5][19] + xor_out[84][5][19];
assign sum_out[17][5][19] = xor_out[85][5][19] + xor_out[86][5][19] + xor_out[87][5][19] + xor_out[88][5][19] + xor_out[89][5][19];
assign sum_out[18][5][19] = xor_out[90][5][19] + xor_out[91][5][19] + xor_out[92][5][19] + xor_out[93][5][19] + xor_out[94][5][19];
assign sum_out[19][5][19] = xor_out[95][5][19] + xor_out[96][5][19] + xor_out[97][5][19] + xor_out[98][5][19] + xor_out[99][5][19];

assign sum_out[0][5][20] = xor_out[0][5][20] + xor_out[1][5][20] + xor_out[2][5][20] + xor_out[3][5][20] + xor_out[4][5][20];
assign sum_out[1][5][20] = xor_out[5][5][20] + xor_out[6][5][20] + xor_out[7][5][20] + xor_out[8][5][20] + xor_out[9][5][20];
assign sum_out[2][5][20] = xor_out[10][5][20] + xor_out[11][5][20] + xor_out[12][5][20] + xor_out[13][5][20] + xor_out[14][5][20];
assign sum_out[3][5][20] = xor_out[15][5][20] + xor_out[16][5][20] + xor_out[17][5][20] + xor_out[18][5][20] + xor_out[19][5][20];
assign sum_out[4][5][20] = xor_out[20][5][20] + xor_out[21][5][20] + xor_out[22][5][20] + xor_out[23][5][20] + xor_out[24][5][20];
assign sum_out[5][5][20] = xor_out[25][5][20] + xor_out[26][5][20] + xor_out[27][5][20] + xor_out[28][5][20] + xor_out[29][5][20];
assign sum_out[6][5][20] = xor_out[30][5][20] + xor_out[31][5][20] + xor_out[32][5][20] + xor_out[33][5][20] + xor_out[34][5][20];
assign sum_out[7][5][20] = xor_out[35][5][20] + xor_out[36][5][20] + xor_out[37][5][20] + xor_out[38][5][20] + xor_out[39][5][20];
assign sum_out[8][5][20] = xor_out[40][5][20] + xor_out[41][5][20] + xor_out[42][5][20] + xor_out[43][5][20] + xor_out[44][5][20];
assign sum_out[9][5][20] = xor_out[45][5][20] + xor_out[46][5][20] + xor_out[47][5][20] + xor_out[48][5][20] + xor_out[49][5][20];
assign sum_out[10][5][20] = xor_out[50][5][20] + xor_out[51][5][20] + xor_out[52][5][20] + xor_out[53][5][20] + xor_out[54][5][20];
assign sum_out[11][5][20] = xor_out[55][5][20] + xor_out[56][5][20] + xor_out[57][5][20] + xor_out[58][5][20] + xor_out[59][5][20];
assign sum_out[12][5][20] = xor_out[60][5][20] + xor_out[61][5][20] + xor_out[62][5][20] + xor_out[63][5][20] + xor_out[64][5][20];
assign sum_out[13][5][20] = xor_out[65][5][20] + xor_out[66][5][20] + xor_out[67][5][20] + xor_out[68][5][20] + xor_out[69][5][20];
assign sum_out[14][5][20] = xor_out[70][5][20] + xor_out[71][5][20] + xor_out[72][5][20] + xor_out[73][5][20] + xor_out[74][5][20];
assign sum_out[15][5][20] = xor_out[75][5][20] + xor_out[76][5][20] + xor_out[77][5][20] + xor_out[78][5][20] + xor_out[79][5][20];
assign sum_out[16][5][20] = xor_out[80][5][20] + xor_out[81][5][20] + xor_out[82][5][20] + xor_out[83][5][20] + xor_out[84][5][20];
assign sum_out[17][5][20] = xor_out[85][5][20] + xor_out[86][5][20] + xor_out[87][5][20] + xor_out[88][5][20] + xor_out[89][5][20];
assign sum_out[18][5][20] = xor_out[90][5][20] + xor_out[91][5][20] + xor_out[92][5][20] + xor_out[93][5][20] + xor_out[94][5][20];
assign sum_out[19][5][20] = xor_out[95][5][20] + xor_out[96][5][20] + xor_out[97][5][20] + xor_out[98][5][20] + xor_out[99][5][20];

assign sum_out[0][5][21] = xor_out[0][5][21] + xor_out[1][5][21] + xor_out[2][5][21] + xor_out[3][5][21] + xor_out[4][5][21];
assign sum_out[1][5][21] = xor_out[5][5][21] + xor_out[6][5][21] + xor_out[7][5][21] + xor_out[8][5][21] + xor_out[9][5][21];
assign sum_out[2][5][21] = xor_out[10][5][21] + xor_out[11][5][21] + xor_out[12][5][21] + xor_out[13][5][21] + xor_out[14][5][21];
assign sum_out[3][5][21] = xor_out[15][5][21] + xor_out[16][5][21] + xor_out[17][5][21] + xor_out[18][5][21] + xor_out[19][5][21];
assign sum_out[4][5][21] = xor_out[20][5][21] + xor_out[21][5][21] + xor_out[22][5][21] + xor_out[23][5][21] + xor_out[24][5][21];
assign sum_out[5][5][21] = xor_out[25][5][21] + xor_out[26][5][21] + xor_out[27][5][21] + xor_out[28][5][21] + xor_out[29][5][21];
assign sum_out[6][5][21] = xor_out[30][5][21] + xor_out[31][5][21] + xor_out[32][5][21] + xor_out[33][5][21] + xor_out[34][5][21];
assign sum_out[7][5][21] = xor_out[35][5][21] + xor_out[36][5][21] + xor_out[37][5][21] + xor_out[38][5][21] + xor_out[39][5][21];
assign sum_out[8][5][21] = xor_out[40][5][21] + xor_out[41][5][21] + xor_out[42][5][21] + xor_out[43][5][21] + xor_out[44][5][21];
assign sum_out[9][5][21] = xor_out[45][5][21] + xor_out[46][5][21] + xor_out[47][5][21] + xor_out[48][5][21] + xor_out[49][5][21];
assign sum_out[10][5][21] = xor_out[50][5][21] + xor_out[51][5][21] + xor_out[52][5][21] + xor_out[53][5][21] + xor_out[54][5][21];
assign sum_out[11][5][21] = xor_out[55][5][21] + xor_out[56][5][21] + xor_out[57][5][21] + xor_out[58][5][21] + xor_out[59][5][21];
assign sum_out[12][5][21] = xor_out[60][5][21] + xor_out[61][5][21] + xor_out[62][5][21] + xor_out[63][5][21] + xor_out[64][5][21];
assign sum_out[13][5][21] = xor_out[65][5][21] + xor_out[66][5][21] + xor_out[67][5][21] + xor_out[68][5][21] + xor_out[69][5][21];
assign sum_out[14][5][21] = xor_out[70][5][21] + xor_out[71][5][21] + xor_out[72][5][21] + xor_out[73][5][21] + xor_out[74][5][21];
assign sum_out[15][5][21] = xor_out[75][5][21] + xor_out[76][5][21] + xor_out[77][5][21] + xor_out[78][5][21] + xor_out[79][5][21];
assign sum_out[16][5][21] = xor_out[80][5][21] + xor_out[81][5][21] + xor_out[82][5][21] + xor_out[83][5][21] + xor_out[84][5][21];
assign sum_out[17][5][21] = xor_out[85][5][21] + xor_out[86][5][21] + xor_out[87][5][21] + xor_out[88][5][21] + xor_out[89][5][21];
assign sum_out[18][5][21] = xor_out[90][5][21] + xor_out[91][5][21] + xor_out[92][5][21] + xor_out[93][5][21] + xor_out[94][5][21];
assign sum_out[19][5][21] = xor_out[95][5][21] + xor_out[96][5][21] + xor_out[97][5][21] + xor_out[98][5][21] + xor_out[99][5][21];

assign sum_out[0][5][22] = xor_out[0][5][22] + xor_out[1][5][22] + xor_out[2][5][22] + xor_out[3][5][22] + xor_out[4][5][22];
assign sum_out[1][5][22] = xor_out[5][5][22] + xor_out[6][5][22] + xor_out[7][5][22] + xor_out[8][5][22] + xor_out[9][5][22];
assign sum_out[2][5][22] = xor_out[10][5][22] + xor_out[11][5][22] + xor_out[12][5][22] + xor_out[13][5][22] + xor_out[14][5][22];
assign sum_out[3][5][22] = xor_out[15][5][22] + xor_out[16][5][22] + xor_out[17][5][22] + xor_out[18][5][22] + xor_out[19][5][22];
assign sum_out[4][5][22] = xor_out[20][5][22] + xor_out[21][5][22] + xor_out[22][5][22] + xor_out[23][5][22] + xor_out[24][5][22];
assign sum_out[5][5][22] = xor_out[25][5][22] + xor_out[26][5][22] + xor_out[27][5][22] + xor_out[28][5][22] + xor_out[29][5][22];
assign sum_out[6][5][22] = xor_out[30][5][22] + xor_out[31][5][22] + xor_out[32][5][22] + xor_out[33][5][22] + xor_out[34][5][22];
assign sum_out[7][5][22] = xor_out[35][5][22] + xor_out[36][5][22] + xor_out[37][5][22] + xor_out[38][5][22] + xor_out[39][5][22];
assign sum_out[8][5][22] = xor_out[40][5][22] + xor_out[41][5][22] + xor_out[42][5][22] + xor_out[43][5][22] + xor_out[44][5][22];
assign sum_out[9][5][22] = xor_out[45][5][22] + xor_out[46][5][22] + xor_out[47][5][22] + xor_out[48][5][22] + xor_out[49][5][22];
assign sum_out[10][5][22] = xor_out[50][5][22] + xor_out[51][5][22] + xor_out[52][5][22] + xor_out[53][5][22] + xor_out[54][5][22];
assign sum_out[11][5][22] = xor_out[55][5][22] + xor_out[56][5][22] + xor_out[57][5][22] + xor_out[58][5][22] + xor_out[59][5][22];
assign sum_out[12][5][22] = xor_out[60][5][22] + xor_out[61][5][22] + xor_out[62][5][22] + xor_out[63][5][22] + xor_out[64][5][22];
assign sum_out[13][5][22] = xor_out[65][5][22] + xor_out[66][5][22] + xor_out[67][5][22] + xor_out[68][5][22] + xor_out[69][5][22];
assign sum_out[14][5][22] = xor_out[70][5][22] + xor_out[71][5][22] + xor_out[72][5][22] + xor_out[73][5][22] + xor_out[74][5][22];
assign sum_out[15][5][22] = xor_out[75][5][22] + xor_out[76][5][22] + xor_out[77][5][22] + xor_out[78][5][22] + xor_out[79][5][22];
assign sum_out[16][5][22] = xor_out[80][5][22] + xor_out[81][5][22] + xor_out[82][5][22] + xor_out[83][5][22] + xor_out[84][5][22];
assign sum_out[17][5][22] = xor_out[85][5][22] + xor_out[86][5][22] + xor_out[87][5][22] + xor_out[88][5][22] + xor_out[89][5][22];
assign sum_out[18][5][22] = xor_out[90][5][22] + xor_out[91][5][22] + xor_out[92][5][22] + xor_out[93][5][22] + xor_out[94][5][22];
assign sum_out[19][5][22] = xor_out[95][5][22] + xor_out[96][5][22] + xor_out[97][5][22] + xor_out[98][5][22] + xor_out[99][5][22];

assign sum_out[0][5][23] = xor_out[0][5][23] + xor_out[1][5][23] + xor_out[2][5][23] + xor_out[3][5][23] + xor_out[4][5][23];
assign sum_out[1][5][23] = xor_out[5][5][23] + xor_out[6][5][23] + xor_out[7][5][23] + xor_out[8][5][23] + xor_out[9][5][23];
assign sum_out[2][5][23] = xor_out[10][5][23] + xor_out[11][5][23] + xor_out[12][5][23] + xor_out[13][5][23] + xor_out[14][5][23];
assign sum_out[3][5][23] = xor_out[15][5][23] + xor_out[16][5][23] + xor_out[17][5][23] + xor_out[18][5][23] + xor_out[19][5][23];
assign sum_out[4][5][23] = xor_out[20][5][23] + xor_out[21][5][23] + xor_out[22][5][23] + xor_out[23][5][23] + xor_out[24][5][23];
assign sum_out[5][5][23] = xor_out[25][5][23] + xor_out[26][5][23] + xor_out[27][5][23] + xor_out[28][5][23] + xor_out[29][5][23];
assign sum_out[6][5][23] = xor_out[30][5][23] + xor_out[31][5][23] + xor_out[32][5][23] + xor_out[33][5][23] + xor_out[34][5][23];
assign sum_out[7][5][23] = xor_out[35][5][23] + xor_out[36][5][23] + xor_out[37][5][23] + xor_out[38][5][23] + xor_out[39][5][23];
assign sum_out[8][5][23] = xor_out[40][5][23] + xor_out[41][5][23] + xor_out[42][5][23] + xor_out[43][5][23] + xor_out[44][5][23];
assign sum_out[9][5][23] = xor_out[45][5][23] + xor_out[46][5][23] + xor_out[47][5][23] + xor_out[48][5][23] + xor_out[49][5][23];
assign sum_out[10][5][23] = xor_out[50][5][23] + xor_out[51][5][23] + xor_out[52][5][23] + xor_out[53][5][23] + xor_out[54][5][23];
assign sum_out[11][5][23] = xor_out[55][5][23] + xor_out[56][5][23] + xor_out[57][5][23] + xor_out[58][5][23] + xor_out[59][5][23];
assign sum_out[12][5][23] = xor_out[60][5][23] + xor_out[61][5][23] + xor_out[62][5][23] + xor_out[63][5][23] + xor_out[64][5][23];
assign sum_out[13][5][23] = xor_out[65][5][23] + xor_out[66][5][23] + xor_out[67][5][23] + xor_out[68][5][23] + xor_out[69][5][23];
assign sum_out[14][5][23] = xor_out[70][5][23] + xor_out[71][5][23] + xor_out[72][5][23] + xor_out[73][5][23] + xor_out[74][5][23];
assign sum_out[15][5][23] = xor_out[75][5][23] + xor_out[76][5][23] + xor_out[77][5][23] + xor_out[78][5][23] + xor_out[79][5][23];
assign sum_out[16][5][23] = xor_out[80][5][23] + xor_out[81][5][23] + xor_out[82][5][23] + xor_out[83][5][23] + xor_out[84][5][23];
assign sum_out[17][5][23] = xor_out[85][5][23] + xor_out[86][5][23] + xor_out[87][5][23] + xor_out[88][5][23] + xor_out[89][5][23];
assign sum_out[18][5][23] = xor_out[90][5][23] + xor_out[91][5][23] + xor_out[92][5][23] + xor_out[93][5][23] + xor_out[94][5][23];
assign sum_out[19][5][23] = xor_out[95][5][23] + xor_out[96][5][23] + xor_out[97][5][23] + xor_out[98][5][23] + xor_out[99][5][23];

assign sum_out[0][6][0] = xor_out[0][6][0] + xor_out[1][6][0] + xor_out[2][6][0] + xor_out[3][6][0] + xor_out[4][6][0];
assign sum_out[1][6][0] = xor_out[5][6][0] + xor_out[6][6][0] + xor_out[7][6][0] + xor_out[8][6][0] + xor_out[9][6][0];
assign sum_out[2][6][0] = xor_out[10][6][0] + xor_out[11][6][0] + xor_out[12][6][0] + xor_out[13][6][0] + xor_out[14][6][0];
assign sum_out[3][6][0] = xor_out[15][6][0] + xor_out[16][6][0] + xor_out[17][6][0] + xor_out[18][6][0] + xor_out[19][6][0];
assign sum_out[4][6][0] = xor_out[20][6][0] + xor_out[21][6][0] + xor_out[22][6][0] + xor_out[23][6][0] + xor_out[24][6][0];
assign sum_out[5][6][0] = xor_out[25][6][0] + xor_out[26][6][0] + xor_out[27][6][0] + xor_out[28][6][0] + xor_out[29][6][0];
assign sum_out[6][6][0] = xor_out[30][6][0] + xor_out[31][6][0] + xor_out[32][6][0] + xor_out[33][6][0] + xor_out[34][6][0];
assign sum_out[7][6][0] = xor_out[35][6][0] + xor_out[36][6][0] + xor_out[37][6][0] + xor_out[38][6][0] + xor_out[39][6][0];
assign sum_out[8][6][0] = xor_out[40][6][0] + xor_out[41][6][0] + xor_out[42][6][0] + xor_out[43][6][0] + xor_out[44][6][0];
assign sum_out[9][6][0] = xor_out[45][6][0] + xor_out[46][6][0] + xor_out[47][6][0] + xor_out[48][6][0] + xor_out[49][6][0];
assign sum_out[10][6][0] = xor_out[50][6][0] + xor_out[51][6][0] + xor_out[52][6][0] + xor_out[53][6][0] + xor_out[54][6][0];
assign sum_out[11][6][0] = xor_out[55][6][0] + xor_out[56][6][0] + xor_out[57][6][0] + xor_out[58][6][0] + xor_out[59][6][0];
assign sum_out[12][6][0] = xor_out[60][6][0] + xor_out[61][6][0] + xor_out[62][6][0] + xor_out[63][6][0] + xor_out[64][6][0];
assign sum_out[13][6][0] = xor_out[65][6][0] + xor_out[66][6][0] + xor_out[67][6][0] + xor_out[68][6][0] + xor_out[69][6][0];
assign sum_out[14][6][0] = xor_out[70][6][0] + xor_out[71][6][0] + xor_out[72][6][0] + xor_out[73][6][0] + xor_out[74][6][0];
assign sum_out[15][6][0] = xor_out[75][6][0] + xor_out[76][6][0] + xor_out[77][6][0] + xor_out[78][6][0] + xor_out[79][6][0];
assign sum_out[16][6][0] = xor_out[80][6][0] + xor_out[81][6][0] + xor_out[82][6][0] + xor_out[83][6][0] + xor_out[84][6][0];
assign sum_out[17][6][0] = xor_out[85][6][0] + xor_out[86][6][0] + xor_out[87][6][0] + xor_out[88][6][0] + xor_out[89][6][0];
assign sum_out[18][6][0] = xor_out[90][6][0] + xor_out[91][6][0] + xor_out[92][6][0] + xor_out[93][6][0] + xor_out[94][6][0];
assign sum_out[19][6][0] = xor_out[95][6][0] + xor_out[96][6][0] + xor_out[97][6][0] + xor_out[98][6][0] + xor_out[99][6][0];

assign sum_out[0][6][1] = xor_out[0][6][1] + xor_out[1][6][1] + xor_out[2][6][1] + xor_out[3][6][1] + xor_out[4][6][1];
assign sum_out[1][6][1] = xor_out[5][6][1] + xor_out[6][6][1] + xor_out[7][6][1] + xor_out[8][6][1] + xor_out[9][6][1];
assign sum_out[2][6][1] = xor_out[10][6][1] + xor_out[11][6][1] + xor_out[12][6][1] + xor_out[13][6][1] + xor_out[14][6][1];
assign sum_out[3][6][1] = xor_out[15][6][1] + xor_out[16][6][1] + xor_out[17][6][1] + xor_out[18][6][1] + xor_out[19][6][1];
assign sum_out[4][6][1] = xor_out[20][6][1] + xor_out[21][6][1] + xor_out[22][6][1] + xor_out[23][6][1] + xor_out[24][6][1];
assign sum_out[5][6][1] = xor_out[25][6][1] + xor_out[26][6][1] + xor_out[27][6][1] + xor_out[28][6][1] + xor_out[29][6][1];
assign sum_out[6][6][1] = xor_out[30][6][1] + xor_out[31][6][1] + xor_out[32][6][1] + xor_out[33][6][1] + xor_out[34][6][1];
assign sum_out[7][6][1] = xor_out[35][6][1] + xor_out[36][6][1] + xor_out[37][6][1] + xor_out[38][6][1] + xor_out[39][6][1];
assign sum_out[8][6][1] = xor_out[40][6][1] + xor_out[41][6][1] + xor_out[42][6][1] + xor_out[43][6][1] + xor_out[44][6][1];
assign sum_out[9][6][1] = xor_out[45][6][1] + xor_out[46][6][1] + xor_out[47][6][1] + xor_out[48][6][1] + xor_out[49][6][1];
assign sum_out[10][6][1] = xor_out[50][6][1] + xor_out[51][6][1] + xor_out[52][6][1] + xor_out[53][6][1] + xor_out[54][6][1];
assign sum_out[11][6][1] = xor_out[55][6][1] + xor_out[56][6][1] + xor_out[57][6][1] + xor_out[58][6][1] + xor_out[59][6][1];
assign sum_out[12][6][1] = xor_out[60][6][1] + xor_out[61][6][1] + xor_out[62][6][1] + xor_out[63][6][1] + xor_out[64][6][1];
assign sum_out[13][6][1] = xor_out[65][6][1] + xor_out[66][6][1] + xor_out[67][6][1] + xor_out[68][6][1] + xor_out[69][6][1];
assign sum_out[14][6][1] = xor_out[70][6][1] + xor_out[71][6][1] + xor_out[72][6][1] + xor_out[73][6][1] + xor_out[74][6][1];
assign sum_out[15][6][1] = xor_out[75][6][1] + xor_out[76][6][1] + xor_out[77][6][1] + xor_out[78][6][1] + xor_out[79][6][1];
assign sum_out[16][6][1] = xor_out[80][6][1] + xor_out[81][6][1] + xor_out[82][6][1] + xor_out[83][6][1] + xor_out[84][6][1];
assign sum_out[17][6][1] = xor_out[85][6][1] + xor_out[86][6][1] + xor_out[87][6][1] + xor_out[88][6][1] + xor_out[89][6][1];
assign sum_out[18][6][1] = xor_out[90][6][1] + xor_out[91][6][1] + xor_out[92][6][1] + xor_out[93][6][1] + xor_out[94][6][1];
assign sum_out[19][6][1] = xor_out[95][6][1] + xor_out[96][6][1] + xor_out[97][6][1] + xor_out[98][6][1] + xor_out[99][6][1];

assign sum_out[0][6][2] = xor_out[0][6][2] + xor_out[1][6][2] + xor_out[2][6][2] + xor_out[3][6][2] + xor_out[4][6][2];
assign sum_out[1][6][2] = xor_out[5][6][2] + xor_out[6][6][2] + xor_out[7][6][2] + xor_out[8][6][2] + xor_out[9][6][2];
assign sum_out[2][6][2] = xor_out[10][6][2] + xor_out[11][6][2] + xor_out[12][6][2] + xor_out[13][6][2] + xor_out[14][6][2];
assign sum_out[3][6][2] = xor_out[15][6][2] + xor_out[16][6][2] + xor_out[17][6][2] + xor_out[18][6][2] + xor_out[19][6][2];
assign sum_out[4][6][2] = xor_out[20][6][2] + xor_out[21][6][2] + xor_out[22][6][2] + xor_out[23][6][2] + xor_out[24][6][2];
assign sum_out[5][6][2] = xor_out[25][6][2] + xor_out[26][6][2] + xor_out[27][6][2] + xor_out[28][6][2] + xor_out[29][6][2];
assign sum_out[6][6][2] = xor_out[30][6][2] + xor_out[31][6][2] + xor_out[32][6][2] + xor_out[33][6][2] + xor_out[34][6][2];
assign sum_out[7][6][2] = xor_out[35][6][2] + xor_out[36][6][2] + xor_out[37][6][2] + xor_out[38][6][2] + xor_out[39][6][2];
assign sum_out[8][6][2] = xor_out[40][6][2] + xor_out[41][6][2] + xor_out[42][6][2] + xor_out[43][6][2] + xor_out[44][6][2];
assign sum_out[9][6][2] = xor_out[45][6][2] + xor_out[46][6][2] + xor_out[47][6][2] + xor_out[48][6][2] + xor_out[49][6][2];
assign sum_out[10][6][2] = xor_out[50][6][2] + xor_out[51][6][2] + xor_out[52][6][2] + xor_out[53][6][2] + xor_out[54][6][2];
assign sum_out[11][6][2] = xor_out[55][6][2] + xor_out[56][6][2] + xor_out[57][6][2] + xor_out[58][6][2] + xor_out[59][6][2];
assign sum_out[12][6][2] = xor_out[60][6][2] + xor_out[61][6][2] + xor_out[62][6][2] + xor_out[63][6][2] + xor_out[64][6][2];
assign sum_out[13][6][2] = xor_out[65][6][2] + xor_out[66][6][2] + xor_out[67][6][2] + xor_out[68][6][2] + xor_out[69][6][2];
assign sum_out[14][6][2] = xor_out[70][6][2] + xor_out[71][6][2] + xor_out[72][6][2] + xor_out[73][6][2] + xor_out[74][6][2];
assign sum_out[15][6][2] = xor_out[75][6][2] + xor_out[76][6][2] + xor_out[77][6][2] + xor_out[78][6][2] + xor_out[79][6][2];
assign sum_out[16][6][2] = xor_out[80][6][2] + xor_out[81][6][2] + xor_out[82][6][2] + xor_out[83][6][2] + xor_out[84][6][2];
assign sum_out[17][6][2] = xor_out[85][6][2] + xor_out[86][6][2] + xor_out[87][6][2] + xor_out[88][6][2] + xor_out[89][6][2];
assign sum_out[18][6][2] = xor_out[90][6][2] + xor_out[91][6][2] + xor_out[92][6][2] + xor_out[93][6][2] + xor_out[94][6][2];
assign sum_out[19][6][2] = xor_out[95][6][2] + xor_out[96][6][2] + xor_out[97][6][2] + xor_out[98][6][2] + xor_out[99][6][2];

assign sum_out[0][6][3] = xor_out[0][6][3] + xor_out[1][6][3] + xor_out[2][6][3] + xor_out[3][6][3] + xor_out[4][6][3];
assign sum_out[1][6][3] = xor_out[5][6][3] + xor_out[6][6][3] + xor_out[7][6][3] + xor_out[8][6][3] + xor_out[9][6][3];
assign sum_out[2][6][3] = xor_out[10][6][3] + xor_out[11][6][3] + xor_out[12][6][3] + xor_out[13][6][3] + xor_out[14][6][3];
assign sum_out[3][6][3] = xor_out[15][6][3] + xor_out[16][6][3] + xor_out[17][6][3] + xor_out[18][6][3] + xor_out[19][6][3];
assign sum_out[4][6][3] = xor_out[20][6][3] + xor_out[21][6][3] + xor_out[22][6][3] + xor_out[23][6][3] + xor_out[24][6][3];
assign sum_out[5][6][3] = xor_out[25][6][3] + xor_out[26][6][3] + xor_out[27][6][3] + xor_out[28][6][3] + xor_out[29][6][3];
assign sum_out[6][6][3] = xor_out[30][6][3] + xor_out[31][6][3] + xor_out[32][6][3] + xor_out[33][6][3] + xor_out[34][6][3];
assign sum_out[7][6][3] = xor_out[35][6][3] + xor_out[36][6][3] + xor_out[37][6][3] + xor_out[38][6][3] + xor_out[39][6][3];
assign sum_out[8][6][3] = xor_out[40][6][3] + xor_out[41][6][3] + xor_out[42][6][3] + xor_out[43][6][3] + xor_out[44][6][3];
assign sum_out[9][6][3] = xor_out[45][6][3] + xor_out[46][6][3] + xor_out[47][6][3] + xor_out[48][6][3] + xor_out[49][6][3];
assign sum_out[10][6][3] = xor_out[50][6][3] + xor_out[51][6][3] + xor_out[52][6][3] + xor_out[53][6][3] + xor_out[54][6][3];
assign sum_out[11][6][3] = xor_out[55][6][3] + xor_out[56][6][3] + xor_out[57][6][3] + xor_out[58][6][3] + xor_out[59][6][3];
assign sum_out[12][6][3] = xor_out[60][6][3] + xor_out[61][6][3] + xor_out[62][6][3] + xor_out[63][6][3] + xor_out[64][6][3];
assign sum_out[13][6][3] = xor_out[65][6][3] + xor_out[66][6][3] + xor_out[67][6][3] + xor_out[68][6][3] + xor_out[69][6][3];
assign sum_out[14][6][3] = xor_out[70][6][3] + xor_out[71][6][3] + xor_out[72][6][3] + xor_out[73][6][3] + xor_out[74][6][3];
assign sum_out[15][6][3] = xor_out[75][6][3] + xor_out[76][6][3] + xor_out[77][6][3] + xor_out[78][6][3] + xor_out[79][6][3];
assign sum_out[16][6][3] = xor_out[80][6][3] + xor_out[81][6][3] + xor_out[82][6][3] + xor_out[83][6][3] + xor_out[84][6][3];
assign sum_out[17][6][3] = xor_out[85][6][3] + xor_out[86][6][3] + xor_out[87][6][3] + xor_out[88][6][3] + xor_out[89][6][3];
assign sum_out[18][6][3] = xor_out[90][6][3] + xor_out[91][6][3] + xor_out[92][6][3] + xor_out[93][6][3] + xor_out[94][6][3];
assign sum_out[19][6][3] = xor_out[95][6][3] + xor_out[96][6][3] + xor_out[97][6][3] + xor_out[98][6][3] + xor_out[99][6][3];

assign sum_out[0][6][4] = xor_out[0][6][4] + xor_out[1][6][4] + xor_out[2][6][4] + xor_out[3][6][4] + xor_out[4][6][4];
assign sum_out[1][6][4] = xor_out[5][6][4] + xor_out[6][6][4] + xor_out[7][6][4] + xor_out[8][6][4] + xor_out[9][6][4];
assign sum_out[2][6][4] = xor_out[10][6][4] + xor_out[11][6][4] + xor_out[12][6][4] + xor_out[13][6][4] + xor_out[14][6][4];
assign sum_out[3][6][4] = xor_out[15][6][4] + xor_out[16][6][4] + xor_out[17][6][4] + xor_out[18][6][4] + xor_out[19][6][4];
assign sum_out[4][6][4] = xor_out[20][6][4] + xor_out[21][6][4] + xor_out[22][6][4] + xor_out[23][6][4] + xor_out[24][6][4];
assign sum_out[5][6][4] = xor_out[25][6][4] + xor_out[26][6][4] + xor_out[27][6][4] + xor_out[28][6][4] + xor_out[29][6][4];
assign sum_out[6][6][4] = xor_out[30][6][4] + xor_out[31][6][4] + xor_out[32][6][4] + xor_out[33][6][4] + xor_out[34][6][4];
assign sum_out[7][6][4] = xor_out[35][6][4] + xor_out[36][6][4] + xor_out[37][6][4] + xor_out[38][6][4] + xor_out[39][6][4];
assign sum_out[8][6][4] = xor_out[40][6][4] + xor_out[41][6][4] + xor_out[42][6][4] + xor_out[43][6][4] + xor_out[44][6][4];
assign sum_out[9][6][4] = xor_out[45][6][4] + xor_out[46][6][4] + xor_out[47][6][4] + xor_out[48][6][4] + xor_out[49][6][4];
assign sum_out[10][6][4] = xor_out[50][6][4] + xor_out[51][6][4] + xor_out[52][6][4] + xor_out[53][6][4] + xor_out[54][6][4];
assign sum_out[11][6][4] = xor_out[55][6][4] + xor_out[56][6][4] + xor_out[57][6][4] + xor_out[58][6][4] + xor_out[59][6][4];
assign sum_out[12][6][4] = xor_out[60][6][4] + xor_out[61][6][4] + xor_out[62][6][4] + xor_out[63][6][4] + xor_out[64][6][4];
assign sum_out[13][6][4] = xor_out[65][6][4] + xor_out[66][6][4] + xor_out[67][6][4] + xor_out[68][6][4] + xor_out[69][6][4];
assign sum_out[14][6][4] = xor_out[70][6][4] + xor_out[71][6][4] + xor_out[72][6][4] + xor_out[73][6][4] + xor_out[74][6][4];
assign sum_out[15][6][4] = xor_out[75][6][4] + xor_out[76][6][4] + xor_out[77][6][4] + xor_out[78][6][4] + xor_out[79][6][4];
assign sum_out[16][6][4] = xor_out[80][6][4] + xor_out[81][6][4] + xor_out[82][6][4] + xor_out[83][6][4] + xor_out[84][6][4];
assign sum_out[17][6][4] = xor_out[85][6][4] + xor_out[86][6][4] + xor_out[87][6][4] + xor_out[88][6][4] + xor_out[89][6][4];
assign sum_out[18][6][4] = xor_out[90][6][4] + xor_out[91][6][4] + xor_out[92][6][4] + xor_out[93][6][4] + xor_out[94][6][4];
assign sum_out[19][6][4] = xor_out[95][6][4] + xor_out[96][6][4] + xor_out[97][6][4] + xor_out[98][6][4] + xor_out[99][6][4];

assign sum_out[0][6][5] = xor_out[0][6][5] + xor_out[1][6][5] + xor_out[2][6][5] + xor_out[3][6][5] + xor_out[4][6][5];
assign sum_out[1][6][5] = xor_out[5][6][5] + xor_out[6][6][5] + xor_out[7][6][5] + xor_out[8][6][5] + xor_out[9][6][5];
assign sum_out[2][6][5] = xor_out[10][6][5] + xor_out[11][6][5] + xor_out[12][6][5] + xor_out[13][6][5] + xor_out[14][6][5];
assign sum_out[3][6][5] = xor_out[15][6][5] + xor_out[16][6][5] + xor_out[17][6][5] + xor_out[18][6][5] + xor_out[19][6][5];
assign sum_out[4][6][5] = xor_out[20][6][5] + xor_out[21][6][5] + xor_out[22][6][5] + xor_out[23][6][5] + xor_out[24][6][5];
assign sum_out[5][6][5] = xor_out[25][6][5] + xor_out[26][6][5] + xor_out[27][6][5] + xor_out[28][6][5] + xor_out[29][6][5];
assign sum_out[6][6][5] = xor_out[30][6][5] + xor_out[31][6][5] + xor_out[32][6][5] + xor_out[33][6][5] + xor_out[34][6][5];
assign sum_out[7][6][5] = xor_out[35][6][5] + xor_out[36][6][5] + xor_out[37][6][5] + xor_out[38][6][5] + xor_out[39][6][5];
assign sum_out[8][6][5] = xor_out[40][6][5] + xor_out[41][6][5] + xor_out[42][6][5] + xor_out[43][6][5] + xor_out[44][6][5];
assign sum_out[9][6][5] = xor_out[45][6][5] + xor_out[46][6][5] + xor_out[47][6][5] + xor_out[48][6][5] + xor_out[49][6][5];
assign sum_out[10][6][5] = xor_out[50][6][5] + xor_out[51][6][5] + xor_out[52][6][5] + xor_out[53][6][5] + xor_out[54][6][5];
assign sum_out[11][6][5] = xor_out[55][6][5] + xor_out[56][6][5] + xor_out[57][6][5] + xor_out[58][6][5] + xor_out[59][6][5];
assign sum_out[12][6][5] = xor_out[60][6][5] + xor_out[61][6][5] + xor_out[62][6][5] + xor_out[63][6][5] + xor_out[64][6][5];
assign sum_out[13][6][5] = xor_out[65][6][5] + xor_out[66][6][5] + xor_out[67][6][5] + xor_out[68][6][5] + xor_out[69][6][5];
assign sum_out[14][6][5] = xor_out[70][6][5] + xor_out[71][6][5] + xor_out[72][6][5] + xor_out[73][6][5] + xor_out[74][6][5];
assign sum_out[15][6][5] = xor_out[75][6][5] + xor_out[76][6][5] + xor_out[77][6][5] + xor_out[78][6][5] + xor_out[79][6][5];
assign sum_out[16][6][5] = xor_out[80][6][5] + xor_out[81][6][5] + xor_out[82][6][5] + xor_out[83][6][5] + xor_out[84][6][5];
assign sum_out[17][6][5] = xor_out[85][6][5] + xor_out[86][6][5] + xor_out[87][6][5] + xor_out[88][6][5] + xor_out[89][6][5];
assign sum_out[18][6][5] = xor_out[90][6][5] + xor_out[91][6][5] + xor_out[92][6][5] + xor_out[93][6][5] + xor_out[94][6][5];
assign sum_out[19][6][5] = xor_out[95][6][5] + xor_out[96][6][5] + xor_out[97][6][5] + xor_out[98][6][5] + xor_out[99][6][5];

assign sum_out[0][6][6] = xor_out[0][6][6] + xor_out[1][6][6] + xor_out[2][6][6] + xor_out[3][6][6] + xor_out[4][6][6];
assign sum_out[1][6][6] = xor_out[5][6][6] + xor_out[6][6][6] + xor_out[7][6][6] + xor_out[8][6][6] + xor_out[9][6][6];
assign sum_out[2][6][6] = xor_out[10][6][6] + xor_out[11][6][6] + xor_out[12][6][6] + xor_out[13][6][6] + xor_out[14][6][6];
assign sum_out[3][6][6] = xor_out[15][6][6] + xor_out[16][6][6] + xor_out[17][6][6] + xor_out[18][6][6] + xor_out[19][6][6];
assign sum_out[4][6][6] = xor_out[20][6][6] + xor_out[21][6][6] + xor_out[22][6][6] + xor_out[23][6][6] + xor_out[24][6][6];
assign sum_out[5][6][6] = xor_out[25][6][6] + xor_out[26][6][6] + xor_out[27][6][6] + xor_out[28][6][6] + xor_out[29][6][6];
assign sum_out[6][6][6] = xor_out[30][6][6] + xor_out[31][6][6] + xor_out[32][6][6] + xor_out[33][6][6] + xor_out[34][6][6];
assign sum_out[7][6][6] = xor_out[35][6][6] + xor_out[36][6][6] + xor_out[37][6][6] + xor_out[38][6][6] + xor_out[39][6][6];
assign sum_out[8][6][6] = xor_out[40][6][6] + xor_out[41][6][6] + xor_out[42][6][6] + xor_out[43][6][6] + xor_out[44][6][6];
assign sum_out[9][6][6] = xor_out[45][6][6] + xor_out[46][6][6] + xor_out[47][6][6] + xor_out[48][6][6] + xor_out[49][6][6];
assign sum_out[10][6][6] = xor_out[50][6][6] + xor_out[51][6][6] + xor_out[52][6][6] + xor_out[53][6][6] + xor_out[54][6][6];
assign sum_out[11][6][6] = xor_out[55][6][6] + xor_out[56][6][6] + xor_out[57][6][6] + xor_out[58][6][6] + xor_out[59][6][6];
assign sum_out[12][6][6] = xor_out[60][6][6] + xor_out[61][6][6] + xor_out[62][6][6] + xor_out[63][6][6] + xor_out[64][6][6];
assign sum_out[13][6][6] = xor_out[65][6][6] + xor_out[66][6][6] + xor_out[67][6][6] + xor_out[68][6][6] + xor_out[69][6][6];
assign sum_out[14][6][6] = xor_out[70][6][6] + xor_out[71][6][6] + xor_out[72][6][6] + xor_out[73][6][6] + xor_out[74][6][6];
assign sum_out[15][6][6] = xor_out[75][6][6] + xor_out[76][6][6] + xor_out[77][6][6] + xor_out[78][6][6] + xor_out[79][6][6];
assign sum_out[16][6][6] = xor_out[80][6][6] + xor_out[81][6][6] + xor_out[82][6][6] + xor_out[83][6][6] + xor_out[84][6][6];
assign sum_out[17][6][6] = xor_out[85][6][6] + xor_out[86][6][6] + xor_out[87][6][6] + xor_out[88][6][6] + xor_out[89][6][6];
assign sum_out[18][6][6] = xor_out[90][6][6] + xor_out[91][6][6] + xor_out[92][6][6] + xor_out[93][6][6] + xor_out[94][6][6];
assign sum_out[19][6][6] = xor_out[95][6][6] + xor_out[96][6][6] + xor_out[97][6][6] + xor_out[98][6][6] + xor_out[99][6][6];

assign sum_out[0][6][7] = xor_out[0][6][7] + xor_out[1][6][7] + xor_out[2][6][7] + xor_out[3][6][7] + xor_out[4][6][7];
assign sum_out[1][6][7] = xor_out[5][6][7] + xor_out[6][6][7] + xor_out[7][6][7] + xor_out[8][6][7] + xor_out[9][6][7];
assign sum_out[2][6][7] = xor_out[10][6][7] + xor_out[11][6][7] + xor_out[12][6][7] + xor_out[13][6][7] + xor_out[14][6][7];
assign sum_out[3][6][7] = xor_out[15][6][7] + xor_out[16][6][7] + xor_out[17][6][7] + xor_out[18][6][7] + xor_out[19][6][7];
assign sum_out[4][6][7] = xor_out[20][6][7] + xor_out[21][6][7] + xor_out[22][6][7] + xor_out[23][6][7] + xor_out[24][6][7];
assign sum_out[5][6][7] = xor_out[25][6][7] + xor_out[26][6][7] + xor_out[27][6][7] + xor_out[28][6][7] + xor_out[29][6][7];
assign sum_out[6][6][7] = xor_out[30][6][7] + xor_out[31][6][7] + xor_out[32][6][7] + xor_out[33][6][7] + xor_out[34][6][7];
assign sum_out[7][6][7] = xor_out[35][6][7] + xor_out[36][6][7] + xor_out[37][6][7] + xor_out[38][6][7] + xor_out[39][6][7];
assign sum_out[8][6][7] = xor_out[40][6][7] + xor_out[41][6][7] + xor_out[42][6][7] + xor_out[43][6][7] + xor_out[44][6][7];
assign sum_out[9][6][7] = xor_out[45][6][7] + xor_out[46][6][7] + xor_out[47][6][7] + xor_out[48][6][7] + xor_out[49][6][7];
assign sum_out[10][6][7] = xor_out[50][6][7] + xor_out[51][6][7] + xor_out[52][6][7] + xor_out[53][6][7] + xor_out[54][6][7];
assign sum_out[11][6][7] = xor_out[55][6][7] + xor_out[56][6][7] + xor_out[57][6][7] + xor_out[58][6][7] + xor_out[59][6][7];
assign sum_out[12][6][7] = xor_out[60][6][7] + xor_out[61][6][7] + xor_out[62][6][7] + xor_out[63][6][7] + xor_out[64][6][7];
assign sum_out[13][6][7] = xor_out[65][6][7] + xor_out[66][6][7] + xor_out[67][6][7] + xor_out[68][6][7] + xor_out[69][6][7];
assign sum_out[14][6][7] = xor_out[70][6][7] + xor_out[71][6][7] + xor_out[72][6][7] + xor_out[73][6][7] + xor_out[74][6][7];
assign sum_out[15][6][7] = xor_out[75][6][7] + xor_out[76][6][7] + xor_out[77][6][7] + xor_out[78][6][7] + xor_out[79][6][7];
assign sum_out[16][6][7] = xor_out[80][6][7] + xor_out[81][6][7] + xor_out[82][6][7] + xor_out[83][6][7] + xor_out[84][6][7];
assign sum_out[17][6][7] = xor_out[85][6][7] + xor_out[86][6][7] + xor_out[87][6][7] + xor_out[88][6][7] + xor_out[89][6][7];
assign sum_out[18][6][7] = xor_out[90][6][7] + xor_out[91][6][7] + xor_out[92][6][7] + xor_out[93][6][7] + xor_out[94][6][7];
assign sum_out[19][6][7] = xor_out[95][6][7] + xor_out[96][6][7] + xor_out[97][6][7] + xor_out[98][6][7] + xor_out[99][6][7];

assign sum_out[0][6][8] = xor_out[0][6][8] + xor_out[1][6][8] + xor_out[2][6][8] + xor_out[3][6][8] + xor_out[4][6][8];
assign sum_out[1][6][8] = xor_out[5][6][8] + xor_out[6][6][8] + xor_out[7][6][8] + xor_out[8][6][8] + xor_out[9][6][8];
assign sum_out[2][6][8] = xor_out[10][6][8] + xor_out[11][6][8] + xor_out[12][6][8] + xor_out[13][6][8] + xor_out[14][6][8];
assign sum_out[3][6][8] = xor_out[15][6][8] + xor_out[16][6][8] + xor_out[17][6][8] + xor_out[18][6][8] + xor_out[19][6][8];
assign sum_out[4][6][8] = xor_out[20][6][8] + xor_out[21][6][8] + xor_out[22][6][8] + xor_out[23][6][8] + xor_out[24][6][8];
assign sum_out[5][6][8] = xor_out[25][6][8] + xor_out[26][6][8] + xor_out[27][6][8] + xor_out[28][6][8] + xor_out[29][6][8];
assign sum_out[6][6][8] = xor_out[30][6][8] + xor_out[31][6][8] + xor_out[32][6][8] + xor_out[33][6][8] + xor_out[34][6][8];
assign sum_out[7][6][8] = xor_out[35][6][8] + xor_out[36][6][8] + xor_out[37][6][8] + xor_out[38][6][8] + xor_out[39][6][8];
assign sum_out[8][6][8] = xor_out[40][6][8] + xor_out[41][6][8] + xor_out[42][6][8] + xor_out[43][6][8] + xor_out[44][6][8];
assign sum_out[9][6][8] = xor_out[45][6][8] + xor_out[46][6][8] + xor_out[47][6][8] + xor_out[48][6][8] + xor_out[49][6][8];
assign sum_out[10][6][8] = xor_out[50][6][8] + xor_out[51][6][8] + xor_out[52][6][8] + xor_out[53][6][8] + xor_out[54][6][8];
assign sum_out[11][6][8] = xor_out[55][6][8] + xor_out[56][6][8] + xor_out[57][6][8] + xor_out[58][6][8] + xor_out[59][6][8];
assign sum_out[12][6][8] = xor_out[60][6][8] + xor_out[61][6][8] + xor_out[62][6][8] + xor_out[63][6][8] + xor_out[64][6][8];
assign sum_out[13][6][8] = xor_out[65][6][8] + xor_out[66][6][8] + xor_out[67][6][8] + xor_out[68][6][8] + xor_out[69][6][8];
assign sum_out[14][6][8] = xor_out[70][6][8] + xor_out[71][6][8] + xor_out[72][6][8] + xor_out[73][6][8] + xor_out[74][6][8];
assign sum_out[15][6][8] = xor_out[75][6][8] + xor_out[76][6][8] + xor_out[77][6][8] + xor_out[78][6][8] + xor_out[79][6][8];
assign sum_out[16][6][8] = xor_out[80][6][8] + xor_out[81][6][8] + xor_out[82][6][8] + xor_out[83][6][8] + xor_out[84][6][8];
assign sum_out[17][6][8] = xor_out[85][6][8] + xor_out[86][6][8] + xor_out[87][6][8] + xor_out[88][6][8] + xor_out[89][6][8];
assign sum_out[18][6][8] = xor_out[90][6][8] + xor_out[91][6][8] + xor_out[92][6][8] + xor_out[93][6][8] + xor_out[94][6][8];
assign sum_out[19][6][8] = xor_out[95][6][8] + xor_out[96][6][8] + xor_out[97][6][8] + xor_out[98][6][8] + xor_out[99][6][8];

assign sum_out[0][6][9] = xor_out[0][6][9] + xor_out[1][6][9] + xor_out[2][6][9] + xor_out[3][6][9] + xor_out[4][6][9];
assign sum_out[1][6][9] = xor_out[5][6][9] + xor_out[6][6][9] + xor_out[7][6][9] + xor_out[8][6][9] + xor_out[9][6][9];
assign sum_out[2][6][9] = xor_out[10][6][9] + xor_out[11][6][9] + xor_out[12][6][9] + xor_out[13][6][9] + xor_out[14][6][9];
assign sum_out[3][6][9] = xor_out[15][6][9] + xor_out[16][6][9] + xor_out[17][6][9] + xor_out[18][6][9] + xor_out[19][6][9];
assign sum_out[4][6][9] = xor_out[20][6][9] + xor_out[21][6][9] + xor_out[22][6][9] + xor_out[23][6][9] + xor_out[24][6][9];
assign sum_out[5][6][9] = xor_out[25][6][9] + xor_out[26][6][9] + xor_out[27][6][9] + xor_out[28][6][9] + xor_out[29][6][9];
assign sum_out[6][6][9] = xor_out[30][6][9] + xor_out[31][6][9] + xor_out[32][6][9] + xor_out[33][6][9] + xor_out[34][6][9];
assign sum_out[7][6][9] = xor_out[35][6][9] + xor_out[36][6][9] + xor_out[37][6][9] + xor_out[38][6][9] + xor_out[39][6][9];
assign sum_out[8][6][9] = xor_out[40][6][9] + xor_out[41][6][9] + xor_out[42][6][9] + xor_out[43][6][9] + xor_out[44][6][9];
assign sum_out[9][6][9] = xor_out[45][6][9] + xor_out[46][6][9] + xor_out[47][6][9] + xor_out[48][6][9] + xor_out[49][6][9];
assign sum_out[10][6][9] = xor_out[50][6][9] + xor_out[51][6][9] + xor_out[52][6][9] + xor_out[53][6][9] + xor_out[54][6][9];
assign sum_out[11][6][9] = xor_out[55][6][9] + xor_out[56][6][9] + xor_out[57][6][9] + xor_out[58][6][9] + xor_out[59][6][9];
assign sum_out[12][6][9] = xor_out[60][6][9] + xor_out[61][6][9] + xor_out[62][6][9] + xor_out[63][6][9] + xor_out[64][6][9];
assign sum_out[13][6][9] = xor_out[65][6][9] + xor_out[66][6][9] + xor_out[67][6][9] + xor_out[68][6][9] + xor_out[69][6][9];
assign sum_out[14][6][9] = xor_out[70][6][9] + xor_out[71][6][9] + xor_out[72][6][9] + xor_out[73][6][9] + xor_out[74][6][9];
assign sum_out[15][6][9] = xor_out[75][6][9] + xor_out[76][6][9] + xor_out[77][6][9] + xor_out[78][6][9] + xor_out[79][6][9];
assign sum_out[16][6][9] = xor_out[80][6][9] + xor_out[81][6][9] + xor_out[82][6][9] + xor_out[83][6][9] + xor_out[84][6][9];
assign sum_out[17][6][9] = xor_out[85][6][9] + xor_out[86][6][9] + xor_out[87][6][9] + xor_out[88][6][9] + xor_out[89][6][9];
assign sum_out[18][6][9] = xor_out[90][6][9] + xor_out[91][6][9] + xor_out[92][6][9] + xor_out[93][6][9] + xor_out[94][6][9];
assign sum_out[19][6][9] = xor_out[95][6][9] + xor_out[96][6][9] + xor_out[97][6][9] + xor_out[98][6][9] + xor_out[99][6][9];

assign sum_out[0][6][10] = xor_out[0][6][10] + xor_out[1][6][10] + xor_out[2][6][10] + xor_out[3][6][10] + xor_out[4][6][10];
assign sum_out[1][6][10] = xor_out[5][6][10] + xor_out[6][6][10] + xor_out[7][6][10] + xor_out[8][6][10] + xor_out[9][6][10];
assign sum_out[2][6][10] = xor_out[10][6][10] + xor_out[11][6][10] + xor_out[12][6][10] + xor_out[13][6][10] + xor_out[14][6][10];
assign sum_out[3][6][10] = xor_out[15][6][10] + xor_out[16][6][10] + xor_out[17][6][10] + xor_out[18][6][10] + xor_out[19][6][10];
assign sum_out[4][6][10] = xor_out[20][6][10] + xor_out[21][6][10] + xor_out[22][6][10] + xor_out[23][6][10] + xor_out[24][6][10];
assign sum_out[5][6][10] = xor_out[25][6][10] + xor_out[26][6][10] + xor_out[27][6][10] + xor_out[28][6][10] + xor_out[29][6][10];
assign sum_out[6][6][10] = xor_out[30][6][10] + xor_out[31][6][10] + xor_out[32][6][10] + xor_out[33][6][10] + xor_out[34][6][10];
assign sum_out[7][6][10] = xor_out[35][6][10] + xor_out[36][6][10] + xor_out[37][6][10] + xor_out[38][6][10] + xor_out[39][6][10];
assign sum_out[8][6][10] = xor_out[40][6][10] + xor_out[41][6][10] + xor_out[42][6][10] + xor_out[43][6][10] + xor_out[44][6][10];
assign sum_out[9][6][10] = xor_out[45][6][10] + xor_out[46][6][10] + xor_out[47][6][10] + xor_out[48][6][10] + xor_out[49][6][10];
assign sum_out[10][6][10] = xor_out[50][6][10] + xor_out[51][6][10] + xor_out[52][6][10] + xor_out[53][6][10] + xor_out[54][6][10];
assign sum_out[11][6][10] = xor_out[55][6][10] + xor_out[56][6][10] + xor_out[57][6][10] + xor_out[58][6][10] + xor_out[59][6][10];
assign sum_out[12][6][10] = xor_out[60][6][10] + xor_out[61][6][10] + xor_out[62][6][10] + xor_out[63][6][10] + xor_out[64][6][10];
assign sum_out[13][6][10] = xor_out[65][6][10] + xor_out[66][6][10] + xor_out[67][6][10] + xor_out[68][6][10] + xor_out[69][6][10];
assign sum_out[14][6][10] = xor_out[70][6][10] + xor_out[71][6][10] + xor_out[72][6][10] + xor_out[73][6][10] + xor_out[74][6][10];
assign sum_out[15][6][10] = xor_out[75][6][10] + xor_out[76][6][10] + xor_out[77][6][10] + xor_out[78][6][10] + xor_out[79][6][10];
assign sum_out[16][6][10] = xor_out[80][6][10] + xor_out[81][6][10] + xor_out[82][6][10] + xor_out[83][6][10] + xor_out[84][6][10];
assign sum_out[17][6][10] = xor_out[85][6][10] + xor_out[86][6][10] + xor_out[87][6][10] + xor_out[88][6][10] + xor_out[89][6][10];
assign sum_out[18][6][10] = xor_out[90][6][10] + xor_out[91][6][10] + xor_out[92][6][10] + xor_out[93][6][10] + xor_out[94][6][10];
assign sum_out[19][6][10] = xor_out[95][6][10] + xor_out[96][6][10] + xor_out[97][6][10] + xor_out[98][6][10] + xor_out[99][6][10];

assign sum_out[0][6][11] = xor_out[0][6][11] + xor_out[1][6][11] + xor_out[2][6][11] + xor_out[3][6][11] + xor_out[4][6][11];
assign sum_out[1][6][11] = xor_out[5][6][11] + xor_out[6][6][11] + xor_out[7][6][11] + xor_out[8][6][11] + xor_out[9][6][11];
assign sum_out[2][6][11] = xor_out[10][6][11] + xor_out[11][6][11] + xor_out[12][6][11] + xor_out[13][6][11] + xor_out[14][6][11];
assign sum_out[3][6][11] = xor_out[15][6][11] + xor_out[16][6][11] + xor_out[17][6][11] + xor_out[18][6][11] + xor_out[19][6][11];
assign sum_out[4][6][11] = xor_out[20][6][11] + xor_out[21][6][11] + xor_out[22][6][11] + xor_out[23][6][11] + xor_out[24][6][11];
assign sum_out[5][6][11] = xor_out[25][6][11] + xor_out[26][6][11] + xor_out[27][6][11] + xor_out[28][6][11] + xor_out[29][6][11];
assign sum_out[6][6][11] = xor_out[30][6][11] + xor_out[31][6][11] + xor_out[32][6][11] + xor_out[33][6][11] + xor_out[34][6][11];
assign sum_out[7][6][11] = xor_out[35][6][11] + xor_out[36][6][11] + xor_out[37][6][11] + xor_out[38][6][11] + xor_out[39][6][11];
assign sum_out[8][6][11] = xor_out[40][6][11] + xor_out[41][6][11] + xor_out[42][6][11] + xor_out[43][6][11] + xor_out[44][6][11];
assign sum_out[9][6][11] = xor_out[45][6][11] + xor_out[46][6][11] + xor_out[47][6][11] + xor_out[48][6][11] + xor_out[49][6][11];
assign sum_out[10][6][11] = xor_out[50][6][11] + xor_out[51][6][11] + xor_out[52][6][11] + xor_out[53][6][11] + xor_out[54][6][11];
assign sum_out[11][6][11] = xor_out[55][6][11] + xor_out[56][6][11] + xor_out[57][6][11] + xor_out[58][6][11] + xor_out[59][6][11];
assign sum_out[12][6][11] = xor_out[60][6][11] + xor_out[61][6][11] + xor_out[62][6][11] + xor_out[63][6][11] + xor_out[64][6][11];
assign sum_out[13][6][11] = xor_out[65][6][11] + xor_out[66][6][11] + xor_out[67][6][11] + xor_out[68][6][11] + xor_out[69][6][11];
assign sum_out[14][6][11] = xor_out[70][6][11] + xor_out[71][6][11] + xor_out[72][6][11] + xor_out[73][6][11] + xor_out[74][6][11];
assign sum_out[15][6][11] = xor_out[75][6][11] + xor_out[76][6][11] + xor_out[77][6][11] + xor_out[78][6][11] + xor_out[79][6][11];
assign sum_out[16][6][11] = xor_out[80][6][11] + xor_out[81][6][11] + xor_out[82][6][11] + xor_out[83][6][11] + xor_out[84][6][11];
assign sum_out[17][6][11] = xor_out[85][6][11] + xor_out[86][6][11] + xor_out[87][6][11] + xor_out[88][6][11] + xor_out[89][6][11];
assign sum_out[18][6][11] = xor_out[90][6][11] + xor_out[91][6][11] + xor_out[92][6][11] + xor_out[93][6][11] + xor_out[94][6][11];
assign sum_out[19][6][11] = xor_out[95][6][11] + xor_out[96][6][11] + xor_out[97][6][11] + xor_out[98][6][11] + xor_out[99][6][11];

assign sum_out[0][6][12] = xor_out[0][6][12] + xor_out[1][6][12] + xor_out[2][6][12] + xor_out[3][6][12] + xor_out[4][6][12];
assign sum_out[1][6][12] = xor_out[5][6][12] + xor_out[6][6][12] + xor_out[7][6][12] + xor_out[8][6][12] + xor_out[9][6][12];
assign sum_out[2][6][12] = xor_out[10][6][12] + xor_out[11][6][12] + xor_out[12][6][12] + xor_out[13][6][12] + xor_out[14][6][12];
assign sum_out[3][6][12] = xor_out[15][6][12] + xor_out[16][6][12] + xor_out[17][6][12] + xor_out[18][6][12] + xor_out[19][6][12];
assign sum_out[4][6][12] = xor_out[20][6][12] + xor_out[21][6][12] + xor_out[22][6][12] + xor_out[23][6][12] + xor_out[24][6][12];
assign sum_out[5][6][12] = xor_out[25][6][12] + xor_out[26][6][12] + xor_out[27][6][12] + xor_out[28][6][12] + xor_out[29][6][12];
assign sum_out[6][6][12] = xor_out[30][6][12] + xor_out[31][6][12] + xor_out[32][6][12] + xor_out[33][6][12] + xor_out[34][6][12];
assign sum_out[7][6][12] = xor_out[35][6][12] + xor_out[36][6][12] + xor_out[37][6][12] + xor_out[38][6][12] + xor_out[39][6][12];
assign sum_out[8][6][12] = xor_out[40][6][12] + xor_out[41][6][12] + xor_out[42][6][12] + xor_out[43][6][12] + xor_out[44][6][12];
assign sum_out[9][6][12] = xor_out[45][6][12] + xor_out[46][6][12] + xor_out[47][6][12] + xor_out[48][6][12] + xor_out[49][6][12];
assign sum_out[10][6][12] = xor_out[50][6][12] + xor_out[51][6][12] + xor_out[52][6][12] + xor_out[53][6][12] + xor_out[54][6][12];
assign sum_out[11][6][12] = xor_out[55][6][12] + xor_out[56][6][12] + xor_out[57][6][12] + xor_out[58][6][12] + xor_out[59][6][12];
assign sum_out[12][6][12] = xor_out[60][6][12] + xor_out[61][6][12] + xor_out[62][6][12] + xor_out[63][6][12] + xor_out[64][6][12];
assign sum_out[13][6][12] = xor_out[65][6][12] + xor_out[66][6][12] + xor_out[67][6][12] + xor_out[68][6][12] + xor_out[69][6][12];
assign sum_out[14][6][12] = xor_out[70][6][12] + xor_out[71][6][12] + xor_out[72][6][12] + xor_out[73][6][12] + xor_out[74][6][12];
assign sum_out[15][6][12] = xor_out[75][6][12] + xor_out[76][6][12] + xor_out[77][6][12] + xor_out[78][6][12] + xor_out[79][6][12];
assign sum_out[16][6][12] = xor_out[80][6][12] + xor_out[81][6][12] + xor_out[82][6][12] + xor_out[83][6][12] + xor_out[84][6][12];
assign sum_out[17][6][12] = xor_out[85][6][12] + xor_out[86][6][12] + xor_out[87][6][12] + xor_out[88][6][12] + xor_out[89][6][12];
assign sum_out[18][6][12] = xor_out[90][6][12] + xor_out[91][6][12] + xor_out[92][6][12] + xor_out[93][6][12] + xor_out[94][6][12];
assign sum_out[19][6][12] = xor_out[95][6][12] + xor_out[96][6][12] + xor_out[97][6][12] + xor_out[98][6][12] + xor_out[99][6][12];

assign sum_out[0][6][13] = xor_out[0][6][13] + xor_out[1][6][13] + xor_out[2][6][13] + xor_out[3][6][13] + xor_out[4][6][13];
assign sum_out[1][6][13] = xor_out[5][6][13] + xor_out[6][6][13] + xor_out[7][6][13] + xor_out[8][6][13] + xor_out[9][6][13];
assign sum_out[2][6][13] = xor_out[10][6][13] + xor_out[11][6][13] + xor_out[12][6][13] + xor_out[13][6][13] + xor_out[14][6][13];
assign sum_out[3][6][13] = xor_out[15][6][13] + xor_out[16][6][13] + xor_out[17][6][13] + xor_out[18][6][13] + xor_out[19][6][13];
assign sum_out[4][6][13] = xor_out[20][6][13] + xor_out[21][6][13] + xor_out[22][6][13] + xor_out[23][6][13] + xor_out[24][6][13];
assign sum_out[5][6][13] = xor_out[25][6][13] + xor_out[26][6][13] + xor_out[27][6][13] + xor_out[28][6][13] + xor_out[29][6][13];
assign sum_out[6][6][13] = xor_out[30][6][13] + xor_out[31][6][13] + xor_out[32][6][13] + xor_out[33][6][13] + xor_out[34][6][13];
assign sum_out[7][6][13] = xor_out[35][6][13] + xor_out[36][6][13] + xor_out[37][6][13] + xor_out[38][6][13] + xor_out[39][6][13];
assign sum_out[8][6][13] = xor_out[40][6][13] + xor_out[41][6][13] + xor_out[42][6][13] + xor_out[43][6][13] + xor_out[44][6][13];
assign sum_out[9][6][13] = xor_out[45][6][13] + xor_out[46][6][13] + xor_out[47][6][13] + xor_out[48][6][13] + xor_out[49][6][13];
assign sum_out[10][6][13] = xor_out[50][6][13] + xor_out[51][6][13] + xor_out[52][6][13] + xor_out[53][6][13] + xor_out[54][6][13];
assign sum_out[11][6][13] = xor_out[55][6][13] + xor_out[56][6][13] + xor_out[57][6][13] + xor_out[58][6][13] + xor_out[59][6][13];
assign sum_out[12][6][13] = xor_out[60][6][13] + xor_out[61][6][13] + xor_out[62][6][13] + xor_out[63][6][13] + xor_out[64][6][13];
assign sum_out[13][6][13] = xor_out[65][6][13] + xor_out[66][6][13] + xor_out[67][6][13] + xor_out[68][6][13] + xor_out[69][6][13];
assign sum_out[14][6][13] = xor_out[70][6][13] + xor_out[71][6][13] + xor_out[72][6][13] + xor_out[73][6][13] + xor_out[74][6][13];
assign sum_out[15][6][13] = xor_out[75][6][13] + xor_out[76][6][13] + xor_out[77][6][13] + xor_out[78][6][13] + xor_out[79][6][13];
assign sum_out[16][6][13] = xor_out[80][6][13] + xor_out[81][6][13] + xor_out[82][6][13] + xor_out[83][6][13] + xor_out[84][6][13];
assign sum_out[17][6][13] = xor_out[85][6][13] + xor_out[86][6][13] + xor_out[87][6][13] + xor_out[88][6][13] + xor_out[89][6][13];
assign sum_out[18][6][13] = xor_out[90][6][13] + xor_out[91][6][13] + xor_out[92][6][13] + xor_out[93][6][13] + xor_out[94][6][13];
assign sum_out[19][6][13] = xor_out[95][6][13] + xor_out[96][6][13] + xor_out[97][6][13] + xor_out[98][6][13] + xor_out[99][6][13];

assign sum_out[0][6][14] = xor_out[0][6][14] + xor_out[1][6][14] + xor_out[2][6][14] + xor_out[3][6][14] + xor_out[4][6][14];
assign sum_out[1][6][14] = xor_out[5][6][14] + xor_out[6][6][14] + xor_out[7][6][14] + xor_out[8][6][14] + xor_out[9][6][14];
assign sum_out[2][6][14] = xor_out[10][6][14] + xor_out[11][6][14] + xor_out[12][6][14] + xor_out[13][6][14] + xor_out[14][6][14];
assign sum_out[3][6][14] = xor_out[15][6][14] + xor_out[16][6][14] + xor_out[17][6][14] + xor_out[18][6][14] + xor_out[19][6][14];
assign sum_out[4][6][14] = xor_out[20][6][14] + xor_out[21][6][14] + xor_out[22][6][14] + xor_out[23][6][14] + xor_out[24][6][14];
assign sum_out[5][6][14] = xor_out[25][6][14] + xor_out[26][6][14] + xor_out[27][6][14] + xor_out[28][6][14] + xor_out[29][6][14];
assign sum_out[6][6][14] = xor_out[30][6][14] + xor_out[31][6][14] + xor_out[32][6][14] + xor_out[33][6][14] + xor_out[34][6][14];
assign sum_out[7][6][14] = xor_out[35][6][14] + xor_out[36][6][14] + xor_out[37][6][14] + xor_out[38][6][14] + xor_out[39][6][14];
assign sum_out[8][6][14] = xor_out[40][6][14] + xor_out[41][6][14] + xor_out[42][6][14] + xor_out[43][6][14] + xor_out[44][6][14];
assign sum_out[9][6][14] = xor_out[45][6][14] + xor_out[46][6][14] + xor_out[47][6][14] + xor_out[48][6][14] + xor_out[49][6][14];
assign sum_out[10][6][14] = xor_out[50][6][14] + xor_out[51][6][14] + xor_out[52][6][14] + xor_out[53][6][14] + xor_out[54][6][14];
assign sum_out[11][6][14] = xor_out[55][6][14] + xor_out[56][6][14] + xor_out[57][6][14] + xor_out[58][6][14] + xor_out[59][6][14];
assign sum_out[12][6][14] = xor_out[60][6][14] + xor_out[61][6][14] + xor_out[62][6][14] + xor_out[63][6][14] + xor_out[64][6][14];
assign sum_out[13][6][14] = xor_out[65][6][14] + xor_out[66][6][14] + xor_out[67][6][14] + xor_out[68][6][14] + xor_out[69][6][14];
assign sum_out[14][6][14] = xor_out[70][6][14] + xor_out[71][6][14] + xor_out[72][6][14] + xor_out[73][6][14] + xor_out[74][6][14];
assign sum_out[15][6][14] = xor_out[75][6][14] + xor_out[76][6][14] + xor_out[77][6][14] + xor_out[78][6][14] + xor_out[79][6][14];
assign sum_out[16][6][14] = xor_out[80][6][14] + xor_out[81][6][14] + xor_out[82][6][14] + xor_out[83][6][14] + xor_out[84][6][14];
assign sum_out[17][6][14] = xor_out[85][6][14] + xor_out[86][6][14] + xor_out[87][6][14] + xor_out[88][6][14] + xor_out[89][6][14];
assign sum_out[18][6][14] = xor_out[90][6][14] + xor_out[91][6][14] + xor_out[92][6][14] + xor_out[93][6][14] + xor_out[94][6][14];
assign sum_out[19][6][14] = xor_out[95][6][14] + xor_out[96][6][14] + xor_out[97][6][14] + xor_out[98][6][14] + xor_out[99][6][14];

assign sum_out[0][6][15] = xor_out[0][6][15] + xor_out[1][6][15] + xor_out[2][6][15] + xor_out[3][6][15] + xor_out[4][6][15];
assign sum_out[1][6][15] = xor_out[5][6][15] + xor_out[6][6][15] + xor_out[7][6][15] + xor_out[8][6][15] + xor_out[9][6][15];
assign sum_out[2][6][15] = xor_out[10][6][15] + xor_out[11][6][15] + xor_out[12][6][15] + xor_out[13][6][15] + xor_out[14][6][15];
assign sum_out[3][6][15] = xor_out[15][6][15] + xor_out[16][6][15] + xor_out[17][6][15] + xor_out[18][6][15] + xor_out[19][6][15];
assign sum_out[4][6][15] = xor_out[20][6][15] + xor_out[21][6][15] + xor_out[22][6][15] + xor_out[23][6][15] + xor_out[24][6][15];
assign sum_out[5][6][15] = xor_out[25][6][15] + xor_out[26][6][15] + xor_out[27][6][15] + xor_out[28][6][15] + xor_out[29][6][15];
assign sum_out[6][6][15] = xor_out[30][6][15] + xor_out[31][6][15] + xor_out[32][6][15] + xor_out[33][6][15] + xor_out[34][6][15];
assign sum_out[7][6][15] = xor_out[35][6][15] + xor_out[36][6][15] + xor_out[37][6][15] + xor_out[38][6][15] + xor_out[39][6][15];
assign sum_out[8][6][15] = xor_out[40][6][15] + xor_out[41][6][15] + xor_out[42][6][15] + xor_out[43][6][15] + xor_out[44][6][15];
assign sum_out[9][6][15] = xor_out[45][6][15] + xor_out[46][6][15] + xor_out[47][6][15] + xor_out[48][6][15] + xor_out[49][6][15];
assign sum_out[10][6][15] = xor_out[50][6][15] + xor_out[51][6][15] + xor_out[52][6][15] + xor_out[53][6][15] + xor_out[54][6][15];
assign sum_out[11][6][15] = xor_out[55][6][15] + xor_out[56][6][15] + xor_out[57][6][15] + xor_out[58][6][15] + xor_out[59][6][15];
assign sum_out[12][6][15] = xor_out[60][6][15] + xor_out[61][6][15] + xor_out[62][6][15] + xor_out[63][6][15] + xor_out[64][6][15];
assign sum_out[13][6][15] = xor_out[65][6][15] + xor_out[66][6][15] + xor_out[67][6][15] + xor_out[68][6][15] + xor_out[69][6][15];
assign sum_out[14][6][15] = xor_out[70][6][15] + xor_out[71][6][15] + xor_out[72][6][15] + xor_out[73][6][15] + xor_out[74][6][15];
assign sum_out[15][6][15] = xor_out[75][6][15] + xor_out[76][6][15] + xor_out[77][6][15] + xor_out[78][6][15] + xor_out[79][6][15];
assign sum_out[16][6][15] = xor_out[80][6][15] + xor_out[81][6][15] + xor_out[82][6][15] + xor_out[83][6][15] + xor_out[84][6][15];
assign sum_out[17][6][15] = xor_out[85][6][15] + xor_out[86][6][15] + xor_out[87][6][15] + xor_out[88][6][15] + xor_out[89][6][15];
assign sum_out[18][6][15] = xor_out[90][6][15] + xor_out[91][6][15] + xor_out[92][6][15] + xor_out[93][6][15] + xor_out[94][6][15];
assign sum_out[19][6][15] = xor_out[95][6][15] + xor_out[96][6][15] + xor_out[97][6][15] + xor_out[98][6][15] + xor_out[99][6][15];

assign sum_out[0][6][16] = xor_out[0][6][16] + xor_out[1][6][16] + xor_out[2][6][16] + xor_out[3][6][16] + xor_out[4][6][16];
assign sum_out[1][6][16] = xor_out[5][6][16] + xor_out[6][6][16] + xor_out[7][6][16] + xor_out[8][6][16] + xor_out[9][6][16];
assign sum_out[2][6][16] = xor_out[10][6][16] + xor_out[11][6][16] + xor_out[12][6][16] + xor_out[13][6][16] + xor_out[14][6][16];
assign sum_out[3][6][16] = xor_out[15][6][16] + xor_out[16][6][16] + xor_out[17][6][16] + xor_out[18][6][16] + xor_out[19][6][16];
assign sum_out[4][6][16] = xor_out[20][6][16] + xor_out[21][6][16] + xor_out[22][6][16] + xor_out[23][6][16] + xor_out[24][6][16];
assign sum_out[5][6][16] = xor_out[25][6][16] + xor_out[26][6][16] + xor_out[27][6][16] + xor_out[28][6][16] + xor_out[29][6][16];
assign sum_out[6][6][16] = xor_out[30][6][16] + xor_out[31][6][16] + xor_out[32][6][16] + xor_out[33][6][16] + xor_out[34][6][16];
assign sum_out[7][6][16] = xor_out[35][6][16] + xor_out[36][6][16] + xor_out[37][6][16] + xor_out[38][6][16] + xor_out[39][6][16];
assign sum_out[8][6][16] = xor_out[40][6][16] + xor_out[41][6][16] + xor_out[42][6][16] + xor_out[43][6][16] + xor_out[44][6][16];
assign sum_out[9][6][16] = xor_out[45][6][16] + xor_out[46][6][16] + xor_out[47][6][16] + xor_out[48][6][16] + xor_out[49][6][16];
assign sum_out[10][6][16] = xor_out[50][6][16] + xor_out[51][6][16] + xor_out[52][6][16] + xor_out[53][6][16] + xor_out[54][6][16];
assign sum_out[11][6][16] = xor_out[55][6][16] + xor_out[56][6][16] + xor_out[57][6][16] + xor_out[58][6][16] + xor_out[59][6][16];
assign sum_out[12][6][16] = xor_out[60][6][16] + xor_out[61][6][16] + xor_out[62][6][16] + xor_out[63][6][16] + xor_out[64][6][16];
assign sum_out[13][6][16] = xor_out[65][6][16] + xor_out[66][6][16] + xor_out[67][6][16] + xor_out[68][6][16] + xor_out[69][6][16];
assign sum_out[14][6][16] = xor_out[70][6][16] + xor_out[71][6][16] + xor_out[72][6][16] + xor_out[73][6][16] + xor_out[74][6][16];
assign sum_out[15][6][16] = xor_out[75][6][16] + xor_out[76][6][16] + xor_out[77][6][16] + xor_out[78][6][16] + xor_out[79][6][16];
assign sum_out[16][6][16] = xor_out[80][6][16] + xor_out[81][6][16] + xor_out[82][6][16] + xor_out[83][6][16] + xor_out[84][6][16];
assign sum_out[17][6][16] = xor_out[85][6][16] + xor_out[86][6][16] + xor_out[87][6][16] + xor_out[88][6][16] + xor_out[89][6][16];
assign sum_out[18][6][16] = xor_out[90][6][16] + xor_out[91][6][16] + xor_out[92][6][16] + xor_out[93][6][16] + xor_out[94][6][16];
assign sum_out[19][6][16] = xor_out[95][6][16] + xor_out[96][6][16] + xor_out[97][6][16] + xor_out[98][6][16] + xor_out[99][6][16];

assign sum_out[0][6][17] = xor_out[0][6][17] + xor_out[1][6][17] + xor_out[2][6][17] + xor_out[3][6][17] + xor_out[4][6][17];
assign sum_out[1][6][17] = xor_out[5][6][17] + xor_out[6][6][17] + xor_out[7][6][17] + xor_out[8][6][17] + xor_out[9][6][17];
assign sum_out[2][6][17] = xor_out[10][6][17] + xor_out[11][6][17] + xor_out[12][6][17] + xor_out[13][6][17] + xor_out[14][6][17];
assign sum_out[3][6][17] = xor_out[15][6][17] + xor_out[16][6][17] + xor_out[17][6][17] + xor_out[18][6][17] + xor_out[19][6][17];
assign sum_out[4][6][17] = xor_out[20][6][17] + xor_out[21][6][17] + xor_out[22][6][17] + xor_out[23][6][17] + xor_out[24][6][17];
assign sum_out[5][6][17] = xor_out[25][6][17] + xor_out[26][6][17] + xor_out[27][6][17] + xor_out[28][6][17] + xor_out[29][6][17];
assign sum_out[6][6][17] = xor_out[30][6][17] + xor_out[31][6][17] + xor_out[32][6][17] + xor_out[33][6][17] + xor_out[34][6][17];
assign sum_out[7][6][17] = xor_out[35][6][17] + xor_out[36][6][17] + xor_out[37][6][17] + xor_out[38][6][17] + xor_out[39][6][17];
assign sum_out[8][6][17] = xor_out[40][6][17] + xor_out[41][6][17] + xor_out[42][6][17] + xor_out[43][6][17] + xor_out[44][6][17];
assign sum_out[9][6][17] = xor_out[45][6][17] + xor_out[46][6][17] + xor_out[47][6][17] + xor_out[48][6][17] + xor_out[49][6][17];
assign sum_out[10][6][17] = xor_out[50][6][17] + xor_out[51][6][17] + xor_out[52][6][17] + xor_out[53][6][17] + xor_out[54][6][17];
assign sum_out[11][6][17] = xor_out[55][6][17] + xor_out[56][6][17] + xor_out[57][6][17] + xor_out[58][6][17] + xor_out[59][6][17];
assign sum_out[12][6][17] = xor_out[60][6][17] + xor_out[61][6][17] + xor_out[62][6][17] + xor_out[63][6][17] + xor_out[64][6][17];
assign sum_out[13][6][17] = xor_out[65][6][17] + xor_out[66][6][17] + xor_out[67][6][17] + xor_out[68][6][17] + xor_out[69][6][17];
assign sum_out[14][6][17] = xor_out[70][6][17] + xor_out[71][6][17] + xor_out[72][6][17] + xor_out[73][6][17] + xor_out[74][6][17];
assign sum_out[15][6][17] = xor_out[75][6][17] + xor_out[76][6][17] + xor_out[77][6][17] + xor_out[78][6][17] + xor_out[79][6][17];
assign sum_out[16][6][17] = xor_out[80][6][17] + xor_out[81][6][17] + xor_out[82][6][17] + xor_out[83][6][17] + xor_out[84][6][17];
assign sum_out[17][6][17] = xor_out[85][6][17] + xor_out[86][6][17] + xor_out[87][6][17] + xor_out[88][6][17] + xor_out[89][6][17];
assign sum_out[18][6][17] = xor_out[90][6][17] + xor_out[91][6][17] + xor_out[92][6][17] + xor_out[93][6][17] + xor_out[94][6][17];
assign sum_out[19][6][17] = xor_out[95][6][17] + xor_out[96][6][17] + xor_out[97][6][17] + xor_out[98][6][17] + xor_out[99][6][17];

assign sum_out[0][6][18] = xor_out[0][6][18] + xor_out[1][6][18] + xor_out[2][6][18] + xor_out[3][6][18] + xor_out[4][6][18];
assign sum_out[1][6][18] = xor_out[5][6][18] + xor_out[6][6][18] + xor_out[7][6][18] + xor_out[8][6][18] + xor_out[9][6][18];
assign sum_out[2][6][18] = xor_out[10][6][18] + xor_out[11][6][18] + xor_out[12][6][18] + xor_out[13][6][18] + xor_out[14][6][18];
assign sum_out[3][6][18] = xor_out[15][6][18] + xor_out[16][6][18] + xor_out[17][6][18] + xor_out[18][6][18] + xor_out[19][6][18];
assign sum_out[4][6][18] = xor_out[20][6][18] + xor_out[21][6][18] + xor_out[22][6][18] + xor_out[23][6][18] + xor_out[24][6][18];
assign sum_out[5][6][18] = xor_out[25][6][18] + xor_out[26][6][18] + xor_out[27][6][18] + xor_out[28][6][18] + xor_out[29][6][18];
assign sum_out[6][6][18] = xor_out[30][6][18] + xor_out[31][6][18] + xor_out[32][6][18] + xor_out[33][6][18] + xor_out[34][6][18];
assign sum_out[7][6][18] = xor_out[35][6][18] + xor_out[36][6][18] + xor_out[37][6][18] + xor_out[38][6][18] + xor_out[39][6][18];
assign sum_out[8][6][18] = xor_out[40][6][18] + xor_out[41][6][18] + xor_out[42][6][18] + xor_out[43][6][18] + xor_out[44][6][18];
assign sum_out[9][6][18] = xor_out[45][6][18] + xor_out[46][6][18] + xor_out[47][6][18] + xor_out[48][6][18] + xor_out[49][6][18];
assign sum_out[10][6][18] = xor_out[50][6][18] + xor_out[51][6][18] + xor_out[52][6][18] + xor_out[53][6][18] + xor_out[54][6][18];
assign sum_out[11][6][18] = xor_out[55][6][18] + xor_out[56][6][18] + xor_out[57][6][18] + xor_out[58][6][18] + xor_out[59][6][18];
assign sum_out[12][6][18] = xor_out[60][6][18] + xor_out[61][6][18] + xor_out[62][6][18] + xor_out[63][6][18] + xor_out[64][6][18];
assign sum_out[13][6][18] = xor_out[65][6][18] + xor_out[66][6][18] + xor_out[67][6][18] + xor_out[68][6][18] + xor_out[69][6][18];
assign sum_out[14][6][18] = xor_out[70][6][18] + xor_out[71][6][18] + xor_out[72][6][18] + xor_out[73][6][18] + xor_out[74][6][18];
assign sum_out[15][6][18] = xor_out[75][6][18] + xor_out[76][6][18] + xor_out[77][6][18] + xor_out[78][6][18] + xor_out[79][6][18];
assign sum_out[16][6][18] = xor_out[80][6][18] + xor_out[81][6][18] + xor_out[82][6][18] + xor_out[83][6][18] + xor_out[84][6][18];
assign sum_out[17][6][18] = xor_out[85][6][18] + xor_out[86][6][18] + xor_out[87][6][18] + xor_out[88][6][18] + xor_out[89][6][18];
assign sum_out[18][6][18] = xor_out[90][6][18] + xor_out[91][6][18] + xor_out[92][6][18] + xor_out[93][6][18] + xor_out[94][6][18];
assign sum_out[19][6][18] = xor_out[95][6][18] + xor_out[96][6][18] + xor_out[97][6][18] + xor_out[98][6][18] + xor_out[99][6][18];

assign sum_out[0][6][19] = xor_out[0][6][19] + xor_out[1][6][19] + xor_out[2][6][19] + xor_out[3][6][19] + xor_out[4][6][19];
assign sum_out[1][6][19] = xor_out[5][6][19] + xor_out[6][6][19] + xor_out[7][6][19] + xor_out[8][6][19] + xor_out[9][6][19];
assign sum_out[2][6][19] = xor_out[10][6][19] + xor_out[11][6][19] + xor_out[12][6][19] + xor_out[13][6][19] + xor_out[14][6][19];
assign sum_out[3][6][19] = xor_out[15][6][19] + xor_out[16][6][19] + xor_out[17][6][19] + xor_out[18][6][19] + xor_out[19][6][19];
assign sum_out[4][6][19] = xor_out[20][6][19] + xor_out[21][6][19] + xor_out[22][6][19] + xor_out[23][6][19] + xor_out[24][6][19];
assign sum_out[5][6][19] = xor_out[25][6][19] + xor_out[26][6][19] + xor_out[27][6][19] + xor_out[28][6][19] + xor_out[29][6][19];
assign sum_out[6][6][19] = xor_out[30][6][19] + xor_out[31][6][19] + xor_out[32][6][19] + xor_out[33][6][19] + xor_out[34][6][19];
assign sum_out[7][6][19] = xor_out[35][6][19] + xor_out[36][6][19] + xor_out[37][6][19] + xor_out[38][6][19] + xor_out[39][6][19];
assign sum_out[8][6][19] = xor_out[40][6][19] + xor_out[41][6][19] + xor_out[42][6][19] + xor_out[43][6][19] + xor_out[44][6][19];
assign sum_out[9][6][19] = xor_out[45][6][19] + xor_out[46][6][19] + xor_out[47][6][19] + xor_out[48][6][19] + xor_out[49][6][19];
assign sum_out[10][6][19] = xor_out[50][6][19] + xor_out[51][6][19] + xor_out[52][6][19] + xor_out[53][6][19] + xor_out[54][6][19];
assign sum_out[11][6][19] = xor_out[55][6][19] + xor_out[56][6][19] + xor_out[57][6][19] + xor_out[58][6][19] + xor_out[59][6][19];
assign sum_out[12][6][19] = xor_out[60][6][19] + xor_out[61][6][19] + xor_out[62][6][19] + xor_out[63][6][19] + xor_out[64][6][19];
assign sum_out[13][6][19] = xor_out[65][6][19] + xor_out[66][6][19] + xor_out[67][6][19] + xor_out[68][6][19] + xor_out[69][6][19];
assign sum_out[14][6][19] = xor_out[70][6][19] + xor_out[71][6][19] + xor_out[72][6][19] + xor_out[73][6][19] + xor_out[74][6][19];
assign sum_out[15][6][19] = xor_out[75][6][19] + xor_out[76][6][19] + xor_out[77][6][19] + xor_out[78][6][19] + xor_out[79][6][19];
assign sum_out[16][6][19] = xor_out[80][6][19] + xor_out[81][6][19] + xor_out[82][6][19] + xor_out[83][6][19] + xor_out[84][6][19];
assign sum_out[17][6][19] = xor_out[85][6][19] + xor_out[86][6][19] + xor_out[87][6][19] + xor_out[88][6][19] + xor_out[89][6][19];
assign sum_out[18][6][19] = xor_out[90][6][19] + xor_out[91][6][19] + xor_out[92][6][19] + xor_out[93][6][19] + xor_out[94][6][19];
assign sum_out[19][6][19] = xor_out[95][6][19] + xor_out[96][6][19] + xor_out[97][6][19] + xor_out[98][6][19] + xor_out[99][6][19];

assign sum_out[0][6][20] = xor_out[0][6][20] + xor_out[1][6][20] + xor_out[2][6][20] + xor_out[3][6][20] + xor_out[4][6][20];
assign sum_out[1][6][20] = xor_out[5][6][20] + xor_out[6][6][20] + xor_out[7][6][20] + xor_out[8][6][20] + xor_out[9][6][20];
assign sum_out[2][6][20] = xor_out[10][6][20] + xor_out[11][6][20] + xor_out[12][6][20] + xor_out[13][6][20] + xor_out[14][6][20];
assign sum_out[3][6][20] = xor_out[15][6][20] + xor_out[16][6][20] + xor_out[17][6][20] + xor_out[18][6][20] + xor_out[19][6][20];
assign sum_out[4][6][20] = xor_out[20][6][20] + xor_out[21][6][20] + xor_out[22][6][20] + xor_out[23][6][20] + xor_out[24][6][20];
assign sum_out[5][6][20] = xor_out[25][6][20] + xor_out[26][6][20] + xor_out[27][6][20] + xor_out[28][6][20] + xor_out[29][6][20];
assign sum_out[6][6][20] = xor_out[30][6][20] + xor_out[31][6][20] + xor_out[32][6][20] + xor_out[33][6][20] + xor_out[34][6][20];
assign sum_out[7][6][20] = xor_out[35][6][20] + xor_out[36][6][20] + xor_out[37][6][20] + xor_out[38][6][20] + xor_out[39][6][20];
assign sum_out[8][6][20] = xor_out[40][6][20] + xor_out[41][6][20] + xor_out[42][6][20] + xor_out[43][6][20] + xor_out[44][6][20];
assign sum_out[9][6][20] = xor_out[45][6][20] + xor_out[46][6][20] + xor_out[47][6][20] + xor_out[48][6][20] + xor_out[49][6][20];
assign sum_out[10][6][20] = xor_out[50][6][20] + xor_out[51][6][20] + xor_out[52][6][20] + xor_out[53][6][20] + xor_out[54][6][20];
assign sum_out[11][6][20] = xor_out[55][6][20] + xor_out[56][6][20] + xor_out[57][6][20] + xor_out[58][6][20] + xor_out[59][6][20];
assign sum_out[12][6][20] = xor_out[60][6][20] + xor_out[61][6][20] + xor_out[62][6][20] + xor_out[63][6][20] + xor_out[64][6][20];
assign sum_out[13][6][20] = xor_out[65][6][20] + xor_out[66][6][20] + xor_out[67][6][20] + xor_out[68][6][20] + xor_out[69][6][20];
assign sum_out[14][6][20] = xor_out[70][6][20] + xor_out[71][6][20] + xor_out[72][6][20] + xor_out[73][6][20] + xor_out[74][6][20];
assign sum_out[15][6][20] = xor_out[75][6][20] + xor_out[76][6][20] + xor_out[77][6][20] + xor_out[78][6][20] + xor_out[79][6][20];
assign sum_out[16][6][20] = xor_out[80][6][20] + xor_out[81][6][20] + xor_out[82][6][20] + xor_out[83][6][20] + xor_out[84][6][20];
assign sum_out[17][6][20] = xor_out[85][6][20] + xor_out[86][6][20] + xor_out[87][6][20] + xor_out[88][6][20] + xor_out[89][6][20];
assign sum_out[18][6][20] = xor_out[90][6][20] + xor_out[91][6][20] + xor_out[92][6][20] + xor_out[93][6][20] + xor_out[94][6][20];
assign sum_out[19][6][20] = xor_out[95][6][20] + xor_out[96][6][20] + xor_out[97][6][20] + xor_out[98][6][20] + xor_out[99][6][20];

assign sum_out[0][6][21] = xor_out[0][6][21] + xor_out[1][6][21] + xor_out[2][6][21] + xor_out[3][6][21] + xor_out[4][6][21];
assign sum_out[1][6][21] = xor_out[5][6][21] + xor_out[6][6][21] + xor_out[7][6][21] + xor_out[8][6][21] + xor_out[9][6][21];
assign sum_out[2][6][21] = xor_out[10][6][21] + xor_out[11][6][21] + xor_out[12][6][21] + xor_out[13][6][21] + xor_out[14][6][21];
assign sum_out[3][6][21] = xor_out[15][6][21] + xor_out[16][6][21] + xor_out[17][6][21] + xor_out[18][6][21] + xor_out[19][6][21];
assign sum_out[4][6][21] = xor_out[20][6][21] + xor_out[21][6][21] + xor_out[22][6][21] + xor_out[23][6][21] + xor_out[24][6][21];
assign sum_out[5][6][21] = xor_out[25][6][21] + xor_out[26][6][21] + xor_out[27][6][21] + xor_out[28][6][21] + xor_out[29][6][21];
assign sum_out[6][6][21] = xor_out[30][6][21] + xor_out[31][6][21] + xor_out[32][6][21] + xor_out[33][6][21] + xor_out[34][6][21];
assign sum_out[7][6][21] = xor_out[35][6][21] + xor_out[36][6][21] + xor_out[37][6][21] + xor_out[38][6][21] + xor_out[39][6][21];
assign sum_out[8][6][21] = xor_out[40][6][21] + xor_out[41][6][21] + xor_out[42][6][21] + xor_out[43][6][21] + xor_out[44][6][21];
assign sum_out[9][6][21] = xor_out[45][6][21] + xor_out[46][6][21] + xor_out[47][6][21] + xor_out[48][6][21] + xor_out[49][6][21];
assign sum_out[10][6][21] = xor_out[50][6][21] + xor_out[51][6][21] + xor_out[52][6][21] + xor_out[53][6][21] + xor_out[54][6][21];
assign sum_out[11][6][21] = xor_out[55][6][21] + xor_out[56][6][21] + xor_out[57][6][21] + xor_out[58][6][21] + xor_out[59][6][21];
assign sum_out[12][6][21] = xor_out[60][6][21] + xor_out[61][6][21] + xor_out[62][6][21] + xor_out[63][6][21] + xor_out[64][6][21];
assign sum_out[13][6][21] = xor_out[65][6][21] + xor_out[66][6][21] + xor_out[67][6][21] + xor_out[68][6][21] + xor_out[69][6][21];
assign sum_out[14][6][21] = xor_out[70][6][21] + xor_out[71][6][21] + xor_out[72][6][21] + xor_out[73][6][21] + xor_out[74][6][21];
assign sum_out[15][6][21] = xor_out[75][6][21] + xor_out[76][6][21] + xor_out[77][6][21] + xor_out[78][6][21] + xor_out[79][6][21];
assign sum_out[16][6][21] = xor_out[80][6][21] + xor_out[81][6][21] + xor_out[82][6][21] + xor_out[83][6][21] + xor_out[84][6][21];
assign sum_out[17][6][21] = xor_out[85][6][21] + xor_out[86][6][21] + xor_out[87][6][21] + xor_out[88][6][21] + xor_out[89][6][21];
assign sum_out[18][6][21] = xor_out[90][6][21] + xor_out[91][6][21] + xor_out[92][6][21] + xor_out[93][6][21] + xor_out[94][6][21];
assign sum_out[19][6][21] = xor_out[95][6][21] + xor_out[96][6][21] + xor_out[97][6][21] + xor_out[98][6][21] + xor_out[99][6][21];

assign sum_out[0][6][22] = xor_out[0][6][22] + xor_out[1][6][22] + xor_out[2][6][22] + xor_out[3][6][22] + xor_out[4][6][22];
assign sum_out[1][6][22] = xor_out[5][6][22] + xor_out[6][6][22] + xor_out[7][6][22] + xor_out[8][6][22] + xor_out[9][6][22];
assign sum_out[2][6][22] = xor_out[10][6][22] + xor_out[11][6][22] + xor_out[12][6][22] + xor_out[13][6][22] + xor_out[14][6][22];
assign sum_out[3][6][22] = xor_out[15][6][22] + xor_out[16][6][22] + xor_out[17][6][22] + xor_out[18][6][22] + xor_out[19][6][22];
assign sum_out[4][6][22] = xor_out[20][6][22] + xor_out[21][6][22] + xor_out[22][6][22] + xor_out[23][6][22] + xor_out[24][6][22];
assign sum_out[5][6][22] = xor_out[25][6][22] + xor_out[26][6][22] + xor_out[27][6][22] + xor_out[28][6][22] + xor_out[29][6][22];
assign sum_out[6][6][22] = xor_out[30][6][22] + xor_out[31][6][22] + xor_out[32][6][22] + xor_out[33][6][22] + xor_out[34][6][22];
assign sum_out[7][6][22] = xor_out[35][6][22] + xor_out[36][6][22] + xor_out[37][6][22] + xor_out[38][6][22] + xor_out[39][6][22];
assign sum_out[8][6][22] = xor_out[40][6][22] + xor_out[41][6][22] + xor_out[42][6][22] + xor_out[43][6][22] + xor_out[44][6][22];
assign sum_out[9][6][22] = xor_out[45][6][22] + xor_out[46][6][22] + xor_out[47][6][22] + xor_out[48][6][22] + xor_out[49][6][22];
assign sum_out[10][6][22] = xor_out[50][6][22] + xor_out[51][6][22] + xor_out[52][6][22] + xor_out[53][6][22] + xor_out[54][6][22];
assign sum_out[11][6][22] = xor_out[55][6][22] + xor_out[56][6][22] + xor_out[57][6][22] + xor_out[58][6][22] + xor_out[59][6][22];
assign sum_out[12][6][22] = xor_out[60][6][22] + xor_out[61][6][22] + xor_out[62][6][22] + xor_out[63][6][22] + xor_out[64][6][22];
assign sum_out[13][6][22] = xor_out[65][6][22] + xor_out[66][6][22] + xor_out[67][6][22] + xor_out[68][6][22] + xor_out[69][6][22];
assign sum_out[14][6][22] = xor_out[70][6][22] + xor_out[71][6][22] + xor_out[72][6][22] + xor_out[73][6][22] + xor_out[74][6][22];
assign sum_out[15][6][22] = xor_out[75][6][22] + xor_out[76][6][22] + xor_out[77][6][22] + xor_out[78][6][22] + xor_out[79][6][22];
assign sum_out[16][6][22] = xor_out[80][6][22] + xor_out[81][6][22] + xor_out[82][6][22] + xor_out[83][6][22] + xor_out[84][6][22];
assign sum_out[17][6][22] = xor_out[85][6][22] + xor_out[86][6][22] + xor_out[87][6][22] + xor_out[88][6][22] + xor_out[89][6][22];
assign sum_out[18][6][22] = xor_out[90][6][22] + xor_out[91][6][22] + xor_out[92][6][22] + xor_out[93][6][22] + xor_out[94][6][22];
assign sum_out[19][6][22] = xor_out[95][6][22] + xor_out[96][6][22] + xor_out[97][6][22] + xor_out[98][6][22] + xor_out[99][6][22];

assign sum_out[0][6][23] = xor_out[0][6][23] + xor_out[1][6][23] + xor_out[2][6][23] + xor_out[3][6][23] + xor_out[4][6][23];
assign sum_out[1][6][23] = xor_out[5][6][23] + xor_out[6][6][23] + xor_out[7][6][23] + xor_out[8][6][23] + xor_out[9][6][23];
assign sum_out[2][6][23] = xor_out[10][6][23] + xor_out[11][6][23] + xor_out[12][6][23] + xor_out[13][6][23] + xor_out[14][6][23];
assign sum_out[3][6][23] = xor_out[15][6][23] + xor_out[16][6][23] + xor_out[17][6][23] + xor_out[18][6][23] + xor_out[19][6][23];
assign sum_out[4][6][23] = xor_out[20][6][23] + xor_out[21][6][23] + xor_out[22][6][23] + xor_out[23][6][23] + xor_out[24][6][23];
assign sum_out[5][6][23] = xor_out[25][6][23] + xor_out[26][6][23] + xor_out[27][6][23] + xor_out[28][6][23] + xor_out[29][6][23];
assign sum_out[6][6][23] = xor_out[30][6][23] + xor_out[31][6][23] + xor_out[32][6][23] + xor_out[33][6][23] + xor_out[34][6][23];
assign sum_out[7][6][23] = xor_out[35][6][23] + xor_out[36][6][23] + xor_out[37][6][23] + xor_out[38][6][23] + xor_out[39][6][23];
assign sum_out[8][6][23] = xor_out[40][6][23] + xor_out[41][6][23] + xor_out[42][6][23] + xor_out[43][6][23] + xor_out[44][6][23];
assign sum_out[9][6][23] = xor_out[45][6][23] + xor_out[46][6][23] + xor_out[47][6][23] + xor_out[48][6][23] + xor_out[49][6][23];
assign sum_out[10][6][23] = xor_out[50][6][23] + xor_out[51][6][23] + xor_out[52][6][23] + xor_out[53][6][23] + xor_out[54][6][23];
assign sum_out[11][6][23] = xor_out[55][6][23] + xor_out[56][6][23] + xor_out[57][6][23] + xor_out[58][6][23] + xor_out[59][6][23];
assign sum_out[12][6][23] = xor_out[60][6][23] + xor_out[61][6][23] + xor_out[62][6][23] + xor_out[63][6][23] + xor_out[64][6][23];
assign sum_out[13][6][23] = xor_out[65][6][23] + xor_out[66][6][23] + xor_out[67][6][23] + xor_out[68][6][23] + xor_out[69][6][23];
assign sum_out[14][6][23] = xor_out[70][6][23] + xor_out[71][6][23] + xor_out[72][6][23] + xor_out[73][6][23] + xor_out[74][6][23];
assign sum_out[15][6][23] = xor_out[75][6][23] + xor_out[76][6][23] + xor_out[77][6][23] + xor_out[78][6][23] + xor_out[79][6][23];
assign sum_out[16][6][23] = xor_out[80][6][23] + xor_out[81][6][23] + xor_out[82][6][23] + xor_out[83][6][23] + xor_out[84][6][23];
assign sum_out[17][6][23] = xor_out[85][6][23] + xor_out[86][6][23] + xor_out[87][6][23] + xor_out[88][6][23] + xor_out[89][6][23];
assign sum_out[18][6][23] = xor_out[90][6][23] + xor_out[91][6][23] + xor_out[92][6][23] + xor_out[93][6][23] + xor_out[94][6][23];
assign sum_out[19][6][23] = xor_out[95][6][23] + xor_out[96][6][23] + xor_out[97][6][23] + xor_out[98][6][23] + xor_out[99][6][23];

assign sum_out[0][7][0] = xor_out[0][7][0] + xor_out[1][7][0] + xor_out[2][7][0] + xor_out[3][7][0] + xor_out[4][7][0];
assign sum_out[1][7][0] = xor_out[5][7][0] + xor_out[6][7][0] + xor_out[7][7][0] + xor_out[8][7][0] + xor_out[9][7][0];
assign sum_out[2][7][0] = xor_out[10][7][0] + xor_out[11][7][0] + xor_out[12][7][0] + xor_out[13][7][0] + xor_out[14][7][0];
assign sum_out[3][7][0] = xor_out[15][7][0] + xor_out[16][7][0] + xor_out[17][7][0] + xor_out[18][7][0] + xor_out[19][7][0];
assign sum_out[4][7][0] = xor_out[20][7][0] + xor_out[21][7][0] + xor_out[22][7][0] + xor_out[23][7][0] + xor_out[24][7][0];
assign sum_out[5][7][0] = xor_out[25][7][0] + xor_out[26][7][0] + xor_out[27][7][0] + xor_out[28][7][0] + xor_out[29][7][0];
assign sum_out[6][7][0] = xor_out[30][7][0] + xor_out[31][7][0] + xor_out[32][7][0] + xor_out[33][7][0] + xor_out[34][7][0];
assign sum_out[7][7][0] = xor_out[35][7][0] + xor_out[36][7][0] + xor_out[37][7][0] + xor_out[38][7][0] + xor_out[39][7][0];
assign sum_out[8][7][0] = xor_out[40][7][0] + xor_out[41][7][0] + xor_out[42][7][0] + xor_out[43][7][0] + xor_out[44][7][0];
assign sum_out[9][7][0] = xor_out[45][7][0] + xor_out[46][7][0] + xor_out[47][7][0] + xor_out[48][7][0] + xor_out[49][7][0];
assign sum_out[10][7][0] = xor_out[50][7][0] + xor_out[51][7][0] + xor_out[52][7][0] + xor_out[53][7][0] + xor_out[54][7][0];
assign sum_out[11][7][0] = xor_out[55][7][0] + xor_out[56][7][0] + xor_out[57][7][0] + xor_out[58][7][0] + xor_out[59][7][0];
assign sum_out[12][7][0] = xor_out[60][7][0] + xor_out[61][7][0] + xor_out[62][7][0] + xor_out[63][7][0] + xor_out[64][7][0];
assign sum_out[13][7][0] = xor_out[65][7][0] + xor_out[66][7][0] + xor_out[67][7][0] + xor_out[68][7][0] + xor_out[69][7][0];
assign sum_out[14][7][0] = xor_out[70][7][0] + xor_out[71][7][0] + xor_out[72][7][0] + xor_out[73][7][0] + xor_out[74][7][0];
assign sum_out[15][7][0] = xor_out[75][7][0] + xor_out[76][7][0] + xor_out[77][7][0] + xor_out[78][7][0] + xor_out[79][7][0];
assign sum_out[16][7][0] = xor_out[80][7][0] + xor_out[81][7][0] + xor_out[82][7][0] + xor_out[83][7][0] + xor_out[84][7][0];
assign sum_out[17][7][0] = xor_out[85][7][0] + xor_out[86][7][0] + xor_out[87][7][0] + xor_out[88][7][0] + xor_out[89][7][0];
assign sum_out[18][7][0] = xor_out[90][7][0] + xor_out[91][7][0] + xor_out[92][7][0] + xor_out[93][7][0] + xor_out[94][7][0];
assign sum_out[19][7][0] = xor_out[95][7][0] + xor_out[96][7][0] + xor_out[97][7][0] + xor_out[98][7][0] + xor_out[99][7][0];

assign sum_out[0][7][1] = xor_out[0][7][1] + xor_out[1][7][1] + xor_out[2][7][1] + xor_out[3][7][1] + xor_out[4][7][1];
assign sum_out[1][7][1] = xor_out[5][7][1] + xor_out[6][7][1] + xor_out[7][7][1] + xor_out[8][7][1] + xor_out[9][7][1];
assign sum_out[2][7][1] = xor_out[10][7][1] + xor_out[11][7][1] + xor_out[12][7][1] + xor_out[13][7][1] + xor_out[14][7][1];
assign sum_out[3][7][1] = xor_out[15][7][1] + xor_out[16][7][1] + xor_out[17][7][1] + xor_out[18][7][1] + xor_out[19][7][1];
assign sum_out[4][7][1] = xor_out[20][7][1] + xor_out[21][7][1] + xor_out[22][7][1] + xor_out[23][7][1] + xor_out[24][7][1];
assign sum_out[5][7][1] = xor_out[25][7][1] + xor_out[26][7][1] + xor_out[27][7][1] + xor_out[28][7][1] + xor_out[29][7][1];
assign sum_out[6][7][1] = xor_out[30][7][1] + xor_out[31][7][1] + xor_out[32][7][1] + xor_out[33][7][1] + xor_out[34][7][1];
assign sum_out[7][7][1] = xor_out[35][7][1] + xor_out[36][7][1] + xor_out[37][7][1] + xor_out[38][7][1] + xor_out[39][7][1];
assign sum_out[8][7][1] = xor_out[40][7][1] + xor_out[41][7][1] + xor_out[42][7][1] + xor_out[43][7][1] + xor_out[44][7][1];
assign sum_out[9][7][1] = xor_out[45][7][1] + xor_out[46][7][1] + xor_out[47][7][1] + xor_out[48][7][1] + xor_out[49][7][1];
assign sum_out[10][7][1] = xor_out[50][7][1] + xor_out[51][7][1] + xor_out[52][7][1] + xor_out[53][7][1] + xor_out[54][7][1];
assign sum_out[11][7][1] = xor_out[55][7][1] + xor_out[56][7][1] + xor_out[57][7][1] + xor_out[58][7][1] + xor_out[59][7][1];
assign sum_out[12][7][1] = xor_out[60][7][1] + xor_out[61][7][1] + xor_out[62][7][1] + xor_out[63][7][1] + xor_out[64][7][1];
assign sum_out[13][7][1] = xor_out[65][7][1] + xor_out[66][7][1] + xor_out[67][7][1] + xor_out[68][7][1] + xor_out[69][7][1];
assign sum_out[14][7][1] = xor_out[70][7][1] + xor_out[71][7][1] + xor_out[72][7][1] + xor_out[73][7][1] + xor_out[74][7][1];
assign sum_out[15][7][1] = xor_out[75][7][1] + xor_out[76][7][1] + xor_out[77][7][1] + xor_out[78][7][1] + xor_out[79][7][1];
assign sum_out[16][7][1] = xor_out[80][7][1] + xor_out[81][7][1] + xor_out[82][7][1] + xor_out[83][7][1] + xor_out[84][7][1];
assign sum_out[17][7][1] = xor_out[85][7][1] + xor_out[86][7][1] + xor_out[87][7][1] + xor_out[88][7][1] + xor_out[89][7][1];
assign sum_out[18][7][1] = xor_out[90][7][1] + xor_out[91][7][1] + xor_out[92][7][1] + xor_out[93][7][1] + xor_out[94][7][1];
assign sum_out[19][7][1] = xor_out[95][7][1] + xor_out[96][7][1] + xor_out[97][7][1] + xor_out[98][7][1] + xor_out[99][7][1];

assign sum_out[0][7][2] = xor_out[0][7][2] + xor_out[1][7][2] + xor_out[2][7][2] + xor_out[3][7][2] + xor_out[4][7][2];
assign sum_out[1][7][2] = xor_out[5][7][2] + xor_out[6][7][2] + xor_out[7][7][2] + xor_out[8][7][2] + xor_out[9][7][2];
assign sum_out[2][7][2] = xor_out[10][7][2] + xor_out[11][7][2] + xor_out[12][7][2] + xor_out[13][7][2] + xor_out[14][7][2];
assign sum_out[3][7][2] = xor_out[15][7][2] + xor_out[16][7][2] + xor_out[17][7][2] + xor_out[18][7][2] + xor_out[19][7][2];
assign sum_out[4][7][2] = xor_out[20][7][2] + xor_out[21][7][2] + xor_out[22][7][2] + xor_out[23][7][2] + xor_out[24][7][2];
assign sum_out[5][7][2] = xor_out[25][7][2] + xor_out[26][7][2] + xor_out[27][7][2] + xor_out[28][7][2] + xor_out[29][7][2];
assign sum_out[6][7][2] = xor_out[30][7][2] + xor_out[31][7][2] + xor_out[32][7][2] + xor_out[33][7][2] + xor_out[34][7][2];
assign sum_out[7][7][2] = xor_out[35][7][2] + xor_out[36][7][2] + xor_out[37][7][2] + xor_out[38][7][2] + xor_out[39][7][2];
assign sum_out[8][7][2] = xor_out[40][7][2] + xor_out[41][7][2] + xor_out[42][7][2] + xor_out[43][7][2] + xor_out[44][7][2];
assign sum_out[9][7][2] = xor_out[45][7][2] + xor_out[46][7][2] + xor_out[47][7][2] + xor_out[48][7][2] + xor_out[49][7][2];
assign sum_out[10][7][2] = xor_out[50][7][2] + xor_out[51][7][2] + xor_out[52][7][2] + xor_out[53][7][2] + xor_out[54][7][2];
assign sum_out[11][7][2] = xor_out[55][7][2] + xor_out[56][7][2] + xor_out[57][7][2] + xor_out[58][7][2] + xor_out[59][7][2];
assign sum_out[12][7][2] = xor_out[60][7][2] + xor_out[61][7][2] + xor_out[62][7][2] + xor_out[63][7][2] + xor_out[64][7][2];
assign sum_out[13][7][2] = xor_out[65][7][2] + xor_out[66][7][2] + xor_out[67][7][2] + xor_out[68][7][2] + xor_out[69][7][2];
assign sum_out[14][7][2] = xor_out[70][7][2] + xor_out[71][7][2] + xor_out[72][7][2] + xor_out[73][7][2] + xor_out[74][7][2];
assign sum_out[15][7][2] = xor_out[75][7][2] + xor_out[76][7][2] + xor_out[77][7][2] + xor_out[78][7][2] + xor_out[79][7][2];
assign sum_out[16][7][2] = xor_out[80][7][2] + xor_out[81][7][2] + xor_out[82][7][2] + xor_out[83][7][2] + xor_out[84][7][2];
assign sum_out[17][7][2] = xor_out[85][7][2] + xor_out[86][7][2] + xor_out[87][7][2] + xor_out[88][7][2] + xor_out[89][7][2];
assign sum_out[18][7][2] = xor_out[90][7][2] + xor_out[91][7][2] + xor_out[92][7][2] + xor_out[93][7][2] + xor_out[94][7][2];
assign sum_out[19][7][2] = xor_out[95][7][2] + xor_out[96][7][2] + xor_out[97][7][2] + xor_out[98][7][2] + xor_out[99][7][2];

assign sum_out[0][7][3] = xor_out[0][7][3] + xor_out[1][7][3] + xor_out[2][7][3] + xor_out[3][7][3] + xor_out[4][7][3];
assign sum_out[1][7][3] = xor_out[5][7][3] + xor_out[6][7][3] + xor_out[7][7][3] + xor_out[8][7][3] + xor_out[9][7][3];
assign sum_out[2][7][3] = xor_out[10][7][3] + xor_out[11][7][3] + xor_out[12][7][3] + xor_out[13][7][3] + xor_out[14][7][3];
assign sum_out[3][7][3] = xor_out[15][7][3] + xor_out[16][7][3] + xor_out[17][7][3] + xor_out[18][7][3] + xor_out[19][7][3];
assign sum_out[4][7][3] = xor_out[20][7][3] + xor_out[21][7][3] + xor_out[22][7][3] + xor_out[23][7][3] + xor_out[24][7][3];
assign sum_out[5][7][3] = xor_out[25][7][3] + xor_out[26][7][3] + xor_out[27][7][3] + xor_out[28][7][3] + xor_out[29][7][3];
assign sum_out[6][7][3] = xor_out[30][7][3] + xor_out[31][7][3] + xor_out[32][7][3] + xor_out[33][7][3] + xor_out[34][7][3];
assign sum_out[7][7][3] = xor_out[35][7][3] + xor_out[36][7][3] + xor_out[37][7][3] + xor_out[38][7][3] + xor_out[39][7][3];
assign sum_out[8][7][3] = xor_out[40][7][3] + xor_out[41][7][3] + xor_out[42][7][3] + xor_out[43][7][3] + xor_out[44][7][3];
assign sum_out[9][7][3] = xor_out[45][7][3] + xor_out[46][7][3] + xor_out[47][7][3] + xor_out[48][7][3] + xor_out[49][7][3];
assign sum_out[10][7][3] = xor_out[50][7][3] + xor_out[51][7][3] + xor_out[52][7][3] + xor_out[53][7][3] + xor_out[54][7][3];
assign sum_out[11][7][3] = xor_out[55][7][3] + xor_out[56][7][3] + xor_out[57][7][3] + xor_out[58][7][3] + xor_out[59][7][3];
assign sum_out[12][7][3] = xor_out[60][7][3] + xor_out[61][7][3] + xor_out[62][7][3] + xor_out[63][7][3] + xor_out[64][7][3];
assign sum_out[13][7][3] = xor_out[65][7][3] + xor_out[66][7][3] + xor_out[67][7][3] + xor_out[68][7][3] + xor_out[69][7][3];
assign sum_out[14][7][3] = xor_out[70][7][3] + xor_out[71][7][3] + xor_out[72][7][3] + xor_out[73][7][3] + xor_out[74][7][3];
assign sum_out[15][7][3] = xor_out[75][7][3] + xor_out[76][7][3] + xor_out[77][7][3] + xor_out[78][7][3] + xor_out[79][7][3];
assign sum_out[16][7][3] = xor_out[80][7][3] + xor_out[81][7][3] + xor_out[82][7][3] + xor_out[83][7][3] + xor_out[84][7][3];
assign sum_out[17][7][3] = xor_out[85][7][3] + xor_out[86][7][3] + xor_out[87][7][3] + xor_out[88][7][3] + xor_out[89][7][3];
assign sum_out[18][7][3] = xor_out[90][7][3] + xor_out[91][7][3] + xor_out[92][7][3] + xor_out[93][7][3] + xor_out[94][7][3];
assign sum_out[19][7][3] = xor_out[95][7][3] + xor_out[96][7][3] + xor_out[97][7][3] + xor_out[98][7][3] + xor_out[99][7][3];

assign sum_out[0][7][4] = xor_out[0][7][4] + xor_out[1][7][4] + xor_out[2][7][4] + xor_out[3][7][4] + xor_out[4][7][4];
assign sum_out[1][7][4] = xor_out[5][7][4] + xor_out[6][7][4] + xor_out[7][7][4] + xor_out[8][7][4] + xor_out[9][7][4];
assign sum_out[2][7][4] = xor_out[10][7][4] + xor_out[11][7][4] + xor_out[12][7][4] + xor_out[13][7][4] + xor_out[14][7][4];
assign sum_out[3][7][4] = xor_out[15][7][4] + xor_out[16][7][4] + xor_out[17][7][4] + xor_out[18][7][4] + xor_out[19][7][4];
assign sum_out[4][7][4] = xor_out[20][7][4] + xor_out[21][7][4] + xor_out[22][7][4] + xor_out[23][7][4] + xor_out[24][7][4];
assign sum_out[5][7][4] = xor_out[25][7][4] + xor_out[26][7][4] + xor_out[27][7][4] + xor_out[28][7][4] + xor_out[29][7][4];
assign sum_out[6][7][4] = xor_out[30][7][4] + xor_out[31][7][4] + xor_out[32][7][4] + xor_out[33][7][4] + xor_out[34][7][4];
assign sum_out[7][7][4] = xor_out[35][7][4] + xor_out[36][7][4] + xor_out[37][7][4] + xor_out[38][7][4] + xor_out[39][7][4];
assign sum_out[8][7][4] = xor_out[40][7][4] + xor_out[41][7][4] + xor_out[42][7][4] + xor_out[43][7][4] + xor_out[44][7][4];
assign sum_out[9][7][4] = xor_out[45][7][4] + xor_out[46][7][4] + xor_out[47][7][4] + xor_out[48][7][4] + xor_out[49][7][4];
assign sum_out[10][7][4] = xor_out[50][7][4] + xor_out[51][7][4] + xor_out[52][7][4] + xor_out[53][7][4] + xor_out[54][7][4];
assign sum_out[11][7][4] = xor_out[55][7][4] + xor_out[56][7][4] + xor_out[57][7][4] + xor_out[58][7][4] + xor_out[59][7][4];
assign sum_out[12][7][4] = xor_out[60][7][4] + xor_out[61][7][4] + xor_out[62][7][4] + xor_out[63][7][4] + xor_out[64][7][4];
assign sum_out[13][7][4] = xor_out[65][7][4] + xor_out[66][7][4] + xor_out[67][7][4] + xor_out[68][7][4] + xor_out[69][7][4];
assign sum_out[14][7][4] = xor_out[70][7][4] + xor_out[71][7][4] + xor_out[72][7][4] + xor_out[73][7][4] + xor_out[74][7][4];
assign sum_out[15][7][4] = xor_out[75][7][4] + xor_out[76][7][4] + xor_out[77][7][4] + xor_out[78][7][4] + xor_out[79][7][4];
assign sum_out[16][7][4] = xor_out[80][7][4] + xor_out[81][7][4] + xor_out[82][7][4] + xor_out[83][7][4] + xor_out[84][7][4];
assign sum_out[17][7][4] = xor_out[85][7][4] + xor_out[86][7][4] + xor_out[87][7][4] + xor_out[88][7][4] + xor_out[89][7][4];
assign sum_out[18][7][4] = xor_out[90][7][4] + xor_out[91][7][4] + xor_out[92][7][4] + xor_out[93][7][4] + xor_out[94][7][4];
assign sum_out[19][7][4] = xor_out[95][7][4] + xor_out[96][7][4] + xor_out[97][7][4] + xor_out[98][7][4] + xor_out[99][7][4];

assign sum_out[0][7][5] = xor_out[0][7][5] + xor_out[1][7][5] + xor_out[2][7][5] + xor_out[3][7][5] + xor_out[4][7][5];
assign sum_out[1][7][5] = xor_out[5][7][5] + xor_out[6][7][5] + xor_out[7][7][5] + xor_out[8][7][5] + xor_out[9][7][5];
assign sum_out[2][7][5] = xor_out[10][7][5] + xor_out[11][7][5] + xor_out[12][7][5] + xor_out[13][7][5] + xor_out[14][7][5];
assign sum_out[3][7][5] = xor_out[15][7][5] + xor_out[16][7][5] + xor_out[17][7][5] + xor_out[18][7][5] + xor_out[19][7][5];
assign sum_out[4][7][5] = xor_out[20][7][5] + xor_out[21][7][5] + xor_out[22][7][5] + xor_out[23][7][5] + xor_out[24][7][5];
assign sum_out[5][7][5] = xor_out[25][7][5] + xor_out[26][7][5] + xor_out[27][7][5] + xor_out[28][7][5] + xor_out[29][7][5];
assign sum_out[6][7][5] = xor_out[30][7][5] + xor_out[31][7][5] + xor_out[32][7][5] + xor_out[33][7][5] + xor_out[34][7][5];
assign sum_out[7][7][5] = xor_out[35][7][5] + xor_out[36][7][5] + xor_out[37][7][5] + xor_out[38][7][5] + xor_out[39][7][5];
assign sum_out[8][7][5] = xor_out[40][7][5] + xor_out[41][7][5] + xor_out[42][7][5] + xor_out[43][7][5] + xor_out[44][7][5];
assign sum_out[9][7][5] = xor_out[45][7][5] + xor_out[46][7][5] + xor_out[47][7][5] + xor_out[48][7][5] + xor_out[49][7][5];
assign sum_out[10][7][5] = xor_out[50][7][5] + xor_out[51][7][5] + xor_out[52][7][5] + xor_out[53][7][5] + xor_out[54][7][5];
assign sum_out[11][7][5] = xor_out[55][7][5] + xor_out[56][7][5] + xor_out[57][7][5] + xor_out[58][7][5] + xor_out[59][7][5];
assign sum_out[12][7][5] = xor_out[60][7][5] + xor_out[61][7][5] + xor_out[62][7][5] + xor_out[63][7][5] + xor_out[64][7][5];
assign sum_out[13][7][5] = xor_out[65][7][5] + xor_out[66][7][5] + xor_out[67][7][5] + xor_out[68][7][5] + xor_out[69][7][5];
assign sum_out[14][7][5] = xor_out[70][7][5] + xor_out[71][7][5] + xor_out[72][7][5] + xor_out[73][7][5] + xor_out[74][7][5];
assign sum_out[15][7][5] = xor_out[75][7][5] + xor_out[76][7][5] + xor_out[77][7][5] + xor_out[78][7][5] + xor_out[79][7][5];
assign sum_out[16][7][5] = xor_out[80][7][5] + xor_out[81][7][5] + xor_out[82][7][5] + xor_out[83][7][5] + xor_out[84][7][5];
assign sum_out[17][7][5] = xor_out[85][7][5] + xor_out[86][7][5] + xor_out[87][7][5] + xor_out[88][7][5] + xor_out[89][7][5];
assign sum_out[18][7][5] = xor_out[90][7][5] + xor_out[91][7][5] + xor_out[92][7][5] + xor_out[93][7][5] + xor_out[94][7][5];
assign sum_out[19][7][5] = xor_out[95][7][5] + xor_out[96][7][5] + xor_out[97][7][5] + xor_out[98][7][5] + xor_out[99][7][5];

assign sum_out[0][7][6] = xor_out[0][7][6] + xor_out[1][7][6] + xor_out[2][7][6] + xor_out[3][7][6] + xor_out[4][7][6];
assign sum_out[1][7][6] = xor_out[5][7][6] + xor_out[6][7][6] + xor_out[7][7][6] + xor_out[8][7][6] + xor_out[9][7][6];
assign sum_out[2][7][6] = xor_out[10][7][6] + xor_out[11][7][6] + xor_out[12][7][6] + xor_out[13][7][6] + xor_out[14][7][6];
assign sum_out[3][7][6] = xor_out[15][7][6] + xor_out[16][7][6] + xor_out[17][7][6] + xor_out[18][7][6] + xor_out[19][7][6];
assign sum_out[4][7][6] = xor_out[20][7][6] + xor_out[21][7][6] + xor_out[22][7][6] + xor_out[23][7][6] + xor_out[24][7][6];
assign sum_out[5][7][6] = xor_out[25][7][6] + xor_out[26][7][6] + xor_out[27][7][6] + xor_out[28][7][6] + xor_out[29][7][6];
assign sum_out[6][7][6] = xor_out[30][7][6] + xor_out[31][7][6] + xor_out[32][7][6] + xor_out[33][7][6] + xor_out[34][7][6];
assign sum_out[7][7][6] = xor_out[35][7][6] + xor_out[36][7][6] + xor_out[37][7][6] + xor_out[38][7][6] + xor_out[39][7][6];
assign sum_out[8][7][6] = xor_out[40][7][6] + xor_out[41][7][6] + xor_out[42][7][6] + xor_out[43][7][6] + xor_out[44][7][6];
assign sum_out[9][7][6] = xor_out[45][7][6] + xor_out[46][7][6] + xor_out[47][7][6] + xor_out[48][7][6] + xor_out[49][7][6];
assign sum_out[10][7][6] = xor_out[50][7][6] + xor_out[51][7][6] + xor_out[52][7][6] + xor_out[53][7][6] + xor_out[54][7][6];
assign sum_out[11][7][6] = xor_out[55][7][6] + xor_out[56][7][6] + xor_out[57][7][6] + xor_out[58][7][6] + xor_out[59][7][6];
assign sum_out[12][7][6] = xor_out[60][7][6] + xor_out[61][7][6] + xor_out[62][7][6] + xor_out[63][7][6] + xor_out[64][7][6];
assign sum_out[13][7][6] = xor_out[65][7][6] + xor_out[66][7][6] + xor_out[67][7][6] + xor_out[68][7][6] + xor_out[69][7][6];
assign sum_out[14][7][6] = xor_out[70][7][6] + xor_out[71][7][6] + xor_out[72][7][6] + xor_out[73][7][6] + xor_out[74][7][6];
assign sum_out[15][7][6] = xor_out[75][7][6] + xor_out[76][7][6] + xor_out[77][7][6] + xor_out[78][7][6] + xor_out[79][7][6];
assign sum_out[16][7][6] = xor_out[80][7][6] + xor_out[81][7][6] + xor_out[82][7][6] + xor_out[83][7][6] + xor_out[84][7][6];
assign sum_out[17][7][6] = xor_out[85][7][6] + xor_out[86][7][6] + xor_out[87][7][6] + xor_out[88][7][6] + xor_out[89][7][6];
assign sum_out[18][7][6] = xor_out[90][7][6] + xor_out[91][7][6] + xor_out[92][7][6] + xor_out[93][7][6] + xor_out[94][7][6];
assign sum_out[19][7][6] = xor_out[95][7][6] + xor_out[96][7][6] + xor_out[97][7][6] + xor_out[98][7][6] + xor_out[99][7][6];

assign sum_out[0][7][7] = xor_out[0][7][7] + xor_out[1][7][7] + xor_out[2][7][7] + xor_out[3][7][7] + xor_out[4][7][7];
assign sum_out[1][7][7] = xor_out[5][7][7] + xor_out[6][7][7] + xor_out[7][7][7] + xor_out[8][7][7] + xor_out[9][7][7];
assign sum_out[2][7][7] = xor_out[10][7][7] + xor_out[11][7][7] + xor_out[12][7][7] + xor_out[13][7][7] + xor_out[14][7][7];
assign sum_out[3][7][7] = xor_out[15][7][7] + xor_out[16][7][7] + xor_out[17][7][7] + xor_out[18][7][7] + xor_out[19][7][7];
assign sum_out[4][7][7] = xor_out[20][7][7] + xor_out[21][7][7] + xor_out[22][7][7] + xor_out[23][7][7] + xor_out[24][7][7];
assign sum_out[5][7][7] = xor_out[25][7][7] + xor_out[26][7][7] + xor_out[27][7][7] + xor_out[28][7][7] + xor_out[29][7][7];
assign sum_out[6][7][7] = xor_out[30][7][7] + xor_out[31][7][7] + xor_out[32][7][7] + xor_out[33][7][7] + xor_out[34][7][7];
assign sum_out[7][7][7] = xor_out[35][7][7] + xor_out[36][7][7] + xor_out[37][7][7] + xor_out[38][7][7] + xor_out[39][7][7];
assign sum_out[8][7][7] = xor_out[40][7][7] + xor_out[41][7][7] + xor_out[42][7][7] + xor_out[43][7][7] + xor_out[44][7][7];
assign sum_out[9][7][7] = xor_out[45][7][7] + xor_out[46][7][7] + xor_out[47][7][7] + xor_out[48][7][7] + xor_out[49][7][7];
assign sum_out[10][7][7] = xor_out[50][7][7] + xor_out[51][7][7] + xor_out[52][7][7] + xor_out[53][7][7] + xor_out[54][7][7];
assign sum_out[11][7][7] = xor_out[55][7][7] + xor_out[56][7][7] + xor_out[57][7][7] + xor_out[58][7][7] + xor_out[59][7][7];
assign sum_out[12][7][7] = xor_out[60][7][7] + xor_out[61][7][7] + xor_out[62][7][7] + xor_out[63][7][7] + xor_out[64][7][7];
assign sum_out[13][7][7] = xor_out[65][7][7] + xor_out[66][7][7] + xor_out[67][7][7] + xor_out[68][7][7] + xor_out[69][7][7];
assign sum_out[14][7][7] = xor_out[70][7][7] + xor_out[71][7][7] + xor_out[72][7][7] + xor_out[73][7][7] + xor_out[74][7][7];
assign sum_out[15][7][7] = xor_out[75][7][7] + xor_out[76][7][7] + xor_out[77][7][7] + xor_out[78][7][7] + xor_out[79][7][7];
assign sum_out[16][7][7] = xor_out[80][7][7] + xor_out[81][7][7] + xor_out[82][7][7] + xor_out[83][7][7] + xor_out[84][7][7];
assign sum_out[17][7][7] = xor_out[85][7][7] + xor_out[86][7][7] + xor_out[87][7][7] + xor_out[88][7][7] + xor_out[89][7][7];
assign sum_out[18][7][7] = xor_out[90][7][7] + xor_out[91][7][7] + xor_out[92][7][7] + xor_out[93][7][7] + xor_out[94][7][7];
assign sum_out[19][7][7] = xor_out[95][7][7] + xor_out[96][7][7] + xor_out[97][7][7] + xor_out[98][7][7] + xor_out[99][7][7];

assign sum_out[0][7][8] = xor_out[0][7][8] + xor_out[1][7][8] + xor_out[2][7][8] + xor_out[3][7][8] + xor_out[4][7][8];
assign sum_out[1][7][8] = xor_out[5][7][8] + xor_out[6][7][8] + xor_out[7][7][8] + xor_out[8][7][8] + xor_out[9][7][8];
assign sum_out[2][7][8] = xor_out[10][7][8] + xor_out[11][7][8] + xor_out[12][7][8] + xor_out[13][7][8] + xor_out[14][7][8];
assign sum_out[3][7][8] = xor_out[15][7][8] + xor_out[16][7][8] + xor_out[17][7][8] + xor_out[18][7][8] + xor_out[19][7][8];
assign sum_out[4][7][8] = xor_out[20][7][8] + xor_out[21][7][8] + xor_out[22][7][8] + xor_out[23][7][8] + xor_out[24][7][8];
assign sum_out[5][7][8] = xor_out[25][7][8] + xor_out[26][7][8] + xor_out[27][7][8] + xor_out[28][7][8] + xor_out[29][7][8];
assign sum_out[6][7][8] = xor_out[30][7][8] + xor_out[31][7][8] + xor_out[32][7][8] + xor_out[33][7][8] + xor_out[34][7][8];
assign sum_out[7][7][8] = xor_out[35][7][8] + xor_out[36][7][8] + xor_out[37][7][8] + xor_out[38][7][8] + xor_out[39][7][8];
assign sum_out[8][7][8] = xor_out[40][7][8] + xor_out[41][7][8] + xor_out[42][7][8] + xor_out[43][7][8] + xor_out[44][7][8];
assign sum_out[9][7][8] = xor_out[45][7][8] + xor_out[46][7][8] + xor_out[47][7][8] + xor_out[48][7][8] + xor_out[49][7][8];
assign sum_out[10][7][8] = xor_out[50][7][8] + xor_out[51][7][8] + xor_out[52][7][8] + xor_out[53][7][8] + xor_out[54][7][8];
assign sum_out[11][7][8] = xor_out[55][7][8] + xor_out[56][7][8] + xor_out[57][7][8] + xor_out[58][7][8] + xor_out[59][7][8];
assign sum_out[12][7][8] = xor_out[60][7][8] + xor_out[61][7][8] + xor_out[62][7][8] + xor_out[63][7][8] + xor_out[64][7][8];
assign sum_out[13][7][8] = xor_out[65][7][8] + xor_out[66][7][8] + xor_out[67][7][8] + xor_out[68][7][8] + xor_out[69][7][8];
assign sum_out[14][7][8] = xor_out[70][7][8] + xor_out[71][7][8] + xor_out[72][7][8] + xor_out[73][7][8] + xor_out[74][7][8];
assign sum_out[15][7][8] = xor_out[75][7][8] + xor_out[76][7][8] + xor_out[77][7][8] + xor_out[78][7][8] + xor_out[79][7][8];
assign sum_out[16][7][8] = xor_out[80][7][8] + xor_out[81][7][8] + xor_out[82][7][8] + xor_out[83][7][8] + xor_out[84][7][8];
assign sum_out[17][7][8] = xor_out[85][7][8] + xor_out[86][7][8] + xor_out[87][7][8] + xor_out[88][7][8] + xor_out[89][7][8];
assign sum_out[18][7][8] = xor_out[90][7][8] + xor_out[91][7][8] + xor_out[92][7][8] + xor_out[93][7][8] + xor_out[94][7][8];
assign sum_out[19][7][8] = xor_out[95][7][8] + xor_out[96][7][8] + xor_out[97][7][8] + xor_out[98][7][8] + xor_out[99][7][8];

assign sum_out[0][7][9] = xor_out[0][7][9] + xor_out[1][7][9] + xor_out[2][7][9] + xor_out[3][7][9] + xor_out[4][7][9];
assign sum_out[1][7][9] = xor_out[5][7][9] + xor_out[6][7][9] + xor_out[7][7][9] + xor_out[8][7][9] + xor_out[9][7][9];
assign sum_out[2][7][9] = xor_out[10][7][9] + xor_out[11][7][9] + xor_out[12][7][9] + xor_out[13][7][9] + xor_out[14][7][9];
assign sum_out[3][7][9] = xor_out[15][7][9] + xor_out[16][7][9] + xor_out[17][7][9] + xor_out[18][7][9] + xor_out[19][7][9];
assign sum_out[4][7][9] = xor_out[20][7][9] + xor_out[21][7][9] + xor_out[22][7][9] + xor_out[23][7][9] + xor_out[24][7][9];
assign sum_out[5][7][9] = xor_out[25][7][9] + xor_out[26][7][9] + xor_out[27][7][9] + xor_out[28][7][9] + xor_out[29][7][9];
assign sum_out[6][7][9] = xor_out[30][7][9] + xor_out[31][7][9] + xor_out[32][7][9] + xor_out[33][7][9] + xor_out[34][7][9];
assign sum_out[7][7][9] = xor_out[35][7][9] + xor_out[36][7][9] + xor_out[37][7][9] + xor_out[38][7][9] + xor_out[39][7][9];
assign sum_out[8][7][9] = xor_out[40][7][9] + xor_out[41][7][9] + xor_out[42][7][9] + xor_out[43][7][9] + xor_out[44][7][9];
assign sum_out[9][7][9] = xor_out[45][7][9] + xor_out[46][7][9] + xor_out[47][7][9] + xor_out[48][7][9] + xor_out[49][7][9];
assign sum_out[10][7][9] = xor_out[50][7][9] + xor_out[51][7][9] + xor_out[52][7][9] + xor_out[53][7][9] + xor_out[54][7][9];
assign sum_out[11][7][9] = xor_out[55][7][9] + xor_out[56][7][9] + xor_out[57][7][9] + xor_out[58][7][9] + xor_out[59][7][9];
assign sum_out[12][7][9] = xor_out[60][7][9] + xor_out[61][7][9] + xor_out[62][7][9] + xor_out[63][7][9] + xor_out[64][7][9];
assign sum_out[13][7][9] = xor_out[65][7][9] + xor_out[66][7][9] + xor_out[67][7][9] + xor_out[68][7][9] + xor_out[69][7][9];
assign sum_out[14][7][9] = xor_out[70][7][9] + xor_out[71][7][9] + xor_out[72][7][9] + xor_out[73][7][9] + xor_out[74][7][9];
assign sum_out[15][7][9] = xor_out[75][7][9] + xor_out[76][7][9] + xor_out[77][7][9] + xor_out[78][7][9] + xor_out[79][7][9];
assign sum_out[16][7][9] = xor_out[80][7][9] + xor_out[81][7][9] + xor_out[82][7][9] + xor_out[83][7][9] + xor_out[84][7][9];
assign sum_out[17][7][9] = xor_out[85][7][9] + xor_out[86][7][9] + xor_out[87][7][9] + xor_out[88][7][9] + xor_out[89][7][9];
assign sum_out[18][7][9] = xor_out[90][7][9] + xor_out[91][7][9] + xor_out[92][7][9] + xor_out[93][7][9] + xor_out[94][7][9];
assign sum_out[19][7][9] = xor_out[95][7][9] + xor_out[96][7][9] + xor_out[97][7][9] + xor_out[98][7][9] + xor_out[99][7][9];

assign sum_out[0][7][10] = xor_out[0][7][10] + xor_out[1][7][10] + xor_out[2][7][10] + xor_out[3][7][10] + xor_out[4][7][10];
assign sum_out[1][7][10] = xor_out[5][7][10] + xor_out[6][7][10] + xor_out[7][7][10] + xor_out[8][7][10] + xor_out[9][7][10];
assign sum_out[2][7][10] = xor_out[10][7][10] + xor_out[11][7][10] + xor_out[12][7][10] + xor_out[13][7][10] + xor_out[14][7][10];
assign sum_out[3][7][10] = xor_out[15][7][10] + xor_out[16][7][10] + xor_out[17][7][10] + xor_out[18][7][10] + xor_out[19][7][10];
assign sum_out[4][7][10] = xor_out[20][7][10] + xor_out[21][7][10] + xor_out[22][7][10] + xor_out[23][7][10] + xor_out[24][7][10];
assign sum_out[5][7][10] = xor_out[25][7][10] + xor_out[26][7][10] + xor_out[27][7][10] + xor_out[28][7][10] + xor_out[29][7][10];
assign sum_out[6][7][10] = xor_out[30][7][10] + xor_out[31][7][10] + xor_out[32][7][10] + xor_out[33][7][10] + xor_out[34][7][10];
assign sum_out[7][7][10] = xor_out[35][7][10] + xor_out[36][7][10] + xor_out[37][7][10] + xor_out[38][7][10] + xor_out[39][7][10];
assign sum_out[8][7][10] = xor_out[40][7][10] + xor_out[41][7][10] + xor_out[42][7][10] + xor_out[43][7][10] + xor_out[44][7][10];
assign sum_out[9][7][10] = xor_out[45][7][10] + xor_out[46][7][10] + xor_out[47][7][10] + xor_out[48][7][10] + xor_out[49][7][10];
assign sum_out[10][7][10] = xor_out[50][7][10] + xor_out[51][7][10] + xor_out[52][7][10] + xor_out[53][7][10] + xor_out[54][7][10];
assign sum_out[11][7][10] = xor_out[55][7][10] + xor_out[56][7][10] + xor_out[57][7][10] + xor_out[58][7][10] + xor_out[59][7][10];
assign sum_out[12][7][10] = xor_out[60][7][10] + xor_out[61][7][10] + xor_out[62][7][10] + xor_out[63][7][10] + xor_out[64][7][10];
assign sum_out[13][7][10] = xor_out[65][7][10] + xor_out[66][7][10] + xor_out[67][7][10] + xor_out[68][7][10] + xor_out[69][7][10];
assign sum_out[14][7][10] = xor_out[70][7][10] + xor_out[71][7][10] + xor_out[72][7][10] + xor_out[73][7][10] + xor_out[74][7][10];
assign sum_out[15][7][10] = xor_out[75][7][10] + xor_out[76][7][10] + xor_out[77][7][10] + xor_out[78][7][10] + xor_out[79][7][10];
assign sum_out[16][7][10] = xor_out[80][7][10] + xor_out[81][7][10] + xor_out[82][7][10] + xor_out[83][7][10] + xor_out[84][7][10];
assign sum_out[17][7][10] = xor_out[85][7][10] + xor_out[86][7][10] + xor_out[87][7][10] + xor_out[88][7][10] + xor_out[89][7][10];
assign sum_out[18][7][10] = xor_out[90][7][10] + xor_out[91][7][10] + xor_out[92][7][10] + xor_out[93][7][10] + xor_out[94][7][10];
assign sum_out[19][7][10] = xor_out[95][7][10] + xor_out[96][7][10] + xor_out[97][7][10] + xor_out[98][7][10] + xor_out[99][7][10];

assign sum_out[0][7][11] = xor_out[0][7][11] + xor_out[1][7][11] + xor_out[2][7][11] + xor_out[3][7][11] + xor_out[4][7][11];
assign sum_out[1][7][11] = xor_out[5][7][11] + xor_out[6][7][11] + xor_out[7][7][11] + xor_out[8][7][11] + xor_out[9][7][11];
assign sum_out[2][7][11] = xor_out[10][7][11] + xor_out[11][7][11] + xor_out[12][7][11] + xor_out[13][7][11] + xor_out[14][7][11];
assign sum_out[3][7][11] = xor_out[15][7][11] + xor_out[16][7][11] + xor_out[17][7][11] + xor_out[18][7][11] + xor_out[19][7][11];
assign sum_out[4][7][11] = xor_out[20][7][11] + xor_out[21][7][11] + xor_out[22][7][11] + xor_out[23][7][11] + xor_out[24][7][11];
assign sum_out[5][7][11] = xor_out[25][7][11] + xor_out[26][7][11] + xor_out[27][7][11] + xor_out[28][7][11] + xor_out[29][7][11];
assign sum_out[6][7][11] = xor_out[30][7][11] + xor_out[31][7][11] + xor_out[32][7][11] + xor_out[33][7][11] + xor_out[34][7][11];
assign sum_out[7][7][11] = xor_out[35][7][11] + xor_out[36][7][11] + xor_out[37][7][11] + xor_out[38][7][11] + xor_out[39][7][11];
assign sum_out[8][7][11] = xor_out[40][7][11] + xor_out[41][7][11] + xor_out[42][7][11] + xor_out[43][7][11] + xor_out[44][7][11];
assign sum_out[9][7][11] = xor_out[45][7][11] + xor_out[46][7][11] + xor_out[47][7][11] + xor_out[48][7][11] + xor_out[49][7][11];
assign sum_out[10][7][11] = xor_out[50][7][11] + xor_out[51][7][11] + xor_out[52][7][11] + xor_out[53][7][11] + xor_out[54][7][11];
assign sum_out[11][7][11] = xor_out[55][7][11] + xor_out[56][7][11] + xor_out[57][7][11] + xor_out[58][7][11] + xor_out[59][7][11];
assign sum_out[12][7][11] = xor_out[60][7][11] + xor_out[61][7][11] + xor_out[62][7][11] + xor_out[63][7][11] + xor_out[64][7][11];
assign sum_out[13][7][11] = xor_out[65][7][11] + xor_out[66][7][11] + xor_out[67][7][11] + xor_out[68][7][11] + xor_out[69][7][11];
assign sum_out[14][7][11] = xor_out[70][7][11] + xor_out[71][7][11] + xor_out[72][7][11] + xor_out[73][7][11] + xor_out[74][7][11];
assign sum_out[15][7][11] = xor_out[75][7][11] + xor_out[76][7][11] + xor_out[77][7][11] + xor_out[78][7][11] + xor_out[79][7][11];
assign sum_out[16][7][11] = xor_out[80][7][11] + xor_out[81][7][11] + xor_out[82][7][11] + xor_out[83][7][11] + xor_out[84][7][11];
assign sum_out[17][7][11] = xor_out[85][7][11] + xor_out[86][7][11] + xor_out[87][7][11] + xor_out[88][7][11] + xor_out[89][7][11];
assign sum_out[18][7][11] = xor_out[90][7][11] + xor_out[91][7][11] + xor_out[92][7][11] + xor_out[93][7][11] + xor_out[94][7][11];
assign sum_out[19][7][11] = xor_out[95][7][11] + xor_out[96][7][11] + xor_out[97][7][11] + xor_out[98][7][11] + xor_out[99][7][11];

assign sum_out[0][7][12] = xor_out[0][7][12] + xor_out[1][7][12] + xor_out[2][7][12] + xor_out[3][7][12] + xor_out[4][7][12];
assign sum_out[1][7][12] = xor_out[5][7][12] + xor_out[6][7][12] + xor_out[7][7][12] + xor_out[8][7][12] + xor_out[9][7][12];
assign sum_out[2][7][12] = xor_out[10][7][12] + xor_out[11][7][12] + xor_out[12][7][12] + xor_out[13][7][12] + xor_out[14][7][12];
assign sum_out[3][7][12] = xor_out[15][7][12] + xor_out[16][7][12] + xor_out[17][7][12] + xor_out[18][7][12] + xor_out[19][7][12];
assign sum_out[4][7][12] = xor_out[20][7][12] + xor_out[21][7][12] + xor_out[22][7][12] + xor_out[23][7][12] + xor_out[24][7][12];
assign sum_out[5][7][12] = xor_out[25][7][12] + xor_out[26][7][12] + xor_out[27][7][12] + xor_out[28][7][12] + xor_out[29][7][12];
assign sum_out[6][7][12] = xor_out[30][7][12] + xor_out[31][7][12] + xor_out[32][7][12] + xor_out[33][7][12] + xor_out[34][7][12];
assign sum_out[7][7][12] = xor_out[35][7][12] + xor_out[36][7][12] + xor_out[37][7][12] + xor_out[38][7][12] + xor_out[39][7][12];
assign sum_out[8][7][12] = xor_out[40][7][12] + xor_out[41][7][12] + xor_out[42][7][12] + xor_out[43][7][12] + xor_out[44][7][12];
assign sum_out[9][7][12] = xor_out[45][7][12] + xor_out[46][7][12] + xor_out[47][7][12] + xor_out[48][7][12] + xor_out[49][7][12];
assign sum_out[10][7][12] = xor_out[50][7][12] + xor_out[51][7][12] + xor_out[52][7][12] + xor_out[53][7][12] + xor_out[54][7][12];
assign sum_out[11][7][12] = xor_out[55][7][12] + xor_out[56][7][12] + xor_out[57][7][12] + xor_out[58][7][12] + xor_out[59][7][12];
assign sum_out[12][7][12] = xor_out[60][7][12] + xor_out[61][7][12] + xor_out[62][7][12] + xor_out[63][7][12] + xor_out[64][7][12];
assign sum_out[13][7][12] = xor_out[65][7][12] + xor_out[66][7][12] + xor_out[67][7][12] + xor_out[68][7][12] + xor_out[69][7][12];
assign sum_out[14][7][12] = xor_out[70][7][12] + xor_out[71][7][12] + xor_out[72][7][12] + xor_out[73][7][12] + xor_out[74][7][12];
assign sum_out[15][7][12] = xor_out[75][7][12] + xor_out[76][7][12] + xor_out[77][7][12] + xor_out[78][7][12] + xor_out[79][7][12];
assign sum_out[16][7][12] = xor_out[80][7][12] + xor_out[81][7][12] + xor_out[82][7][12] + xor_out[83][7][12] + xor_out[84][7][12];
assign sum_out[17][7][12] = xor_out[85][7][12] + xor_out[86][7][12] + xor_out[87][7][12] + xor_out[88][7][12] + xor_out[89][7][12];
assign sum_out[18][7][12] = xor_out[90][7][12] + xor_out[91][7][12] + xor_out[92][7][12] + xor_out[93][7][12] + xor_out[94][7][12];
assign sum_out[19][7][12] = xor_out[95][7][12] + xor_out[96][7][12] + xor_out[97][7][12] + xor_out[98][7][12] + xor_out[99][7][12];

assign sum_out[0][7][13] = xor_out[0][7][13] + xor_out[1][7][13] + xor_out[2][7][13] + xor_out[3][7][13] + xor_out[4][7][13];
assign sum_out[1][7][13] = xor_out[5][7][13] + xor_out[6][7][13] + xor_out[7][7][13] + xor_out[8][7][13] + xor_out[9][7][13];
assign sum_out[2][7][13] = xor_out[10][7][13] + xor_out[11][7][13] + xor_out[12][7][13] + xor_out[13][7][13] + xor_out[14][7][13];
assign sum_out[3][7][13] = xor_out[15][7][13] + xor_out[16][7][13] + xor_out[17][7][13] + xor_out[18][7][13] + xor_out[19][7][13];
assign sum_out[4][7][13] = xor_out[20][7][13] + xor_out[21][7][13] + xor_out[22][7][13] + xor_out[23][7][13] + xor_out[24][7][13];
assign sum_out[5][7][13] = xor_out[25][7][13] + xor_out[26][7][13] + xor_out[27][7][13] + xor_out[28][7][13] + xor_out[29][7][13];
assign sum_out[6][7][13] = xor_out[30][7][13] + xor_out[31][7][13] + xor_out[32][7][13] + xor_out[33][7][13] + xor_out[34][7][13];
assign sum_out[7][7][13] = xor_out[35][7][13] + xor_out[36][7][13] + xor_out[37][7][13] + xor_out[38][7][13] + xor_out[39][7][13];
assign sum_out[8][7][13] = xor_out[40][7][13] + xor_out[41][7][13] + xor_out[42][7][13] + xor_out[43][7][13] + xor_out[44][7][13];
assign sum_out[9][7][13] = xor_out[45][7][13] + xor_out[46][7][13] + xor_out[47][7][13] + xor_out[48][7][13] + xor_out[49][7][13];
assign sum_out[10][7][13] = xor_out[50][7][13] + xor_out[51][7][13] + xor_out[52][7][13] + xor_out[53][7][13] + xor_out[54][7][13];
assign sum_out[11][7][13] = xor_out[55][7][13] + xor_out[56][7][13] + xor_out[57][7][13] + xor_out[58][7][13] + xor_out[59][7][13];
assign sum_out[12][7][13] = xor_out[60][7][13] + xor_out[61][7][13] + xor_out[62][7][13] + xor_out[63][7][13] + xor_out[64][7][13];
assign sum_out[13][7][13] = xor_out[65][7][13] + xor_out[66][7][13] + xor_out[67][7][13] + xor_out[68][7][13] + xor_out[69][7][13];
assign sum_out[14][7][13] = xor_out[70][7][13] + xor_out[71][7][13] + xor_out[72][7][13] + xor_out[73][7][13] + xor_out[74][7][13];
assign sum_out[15][7][13] = xor_out[75][7][13] + xor_out[76][7][13] + xor_out[77][7][13] + xor_out[78][7][13] + xor_out[79][7][13];
assign sum_out[16][7][13] = xor_out[80][7][13] + xor_out[81][7][13] + xor_out[82][7][13] + xor_out[83][7][13] + xor_out[84][7][13];
assign sum_out[17][7][13] = xor_out[85][7][13] + xor_out[86][7][13] + xor_out[87][7][13] + xor_out[88][7][13] + xor_out[89][7][13];
assign sum_out[18][7][13] = xor_out[90][7][13] + xor_out[91][7][13] + xor_out[92][7][13] + xor_out[93][7][13] + xor_out[94][7][13];
assign sum_out[19][7][13] = xor_out[95][7][13] + xor_out[96][7][13] + xor_out[97][7][13] + xor_out[98][7][13] + xor_out[99][7][13];

assign sum_out[0][7][14] = xor_out[0][7][14] + xor_out[1][7][14] + xor_out[2][7][14] + xor_out[3][7][14] + xor_out[4][7][14];
assign sum_out[1][7][14] = xor_out[5][7][14] + xor_out[6][7][14] + xor_out[7][7][14] + xor_out[8][7][14] + xor_out[9][7][14];
assign sum_out[2][7][14] = xor_out[10][7][14] + xor_out[11][7][14] + xor_out[12][7][14] + xor_out[13][7][14] + xor_out[14][7][14];
assign sum_out[3][7][14] = xor_out[15][7][14] + xor_out[16][7][14] + xor_out[17][7][14] + xor_out[18][7][14] + xor_out[19][7][14];
assign sum_out[4][7][14] = xor_out[20][7][14] + xor_out[21][7][14] + xor_out[22][7][14] + xor_out[23][7][14] + xor_out[24][7][14];
assign sum_out[5][7][14] = xor_out[25][7][14] + xor_out[26][7][14] + xor_out[27][7][14] + xor_out[28][7][14] + xor_out[29][7][14];
assign sum_out[6][7][14] = xor_out[30][7][14] + xor_out[31][7][14] + xor_out[32][7][14] + xor_out[33][7][14] + xor_out[34][7][14];
assign sum_out[7][7][14] = xor_out[35][7][14] + xor_out[36][7][14] + xor_out[37][7][14] + xor_out[38][7][14] + xor_out[39][7][14];
assign sum_out[8][7][14] = xor_out[40][7][14] + xor_out[41][7][14] + xor_out[42][7][14] + xor_out[43][7][14] + xor_out[44][7][14];
assign sum_out[9][7][14] = xor_out[45][7][14] + xor_out[46][7][14] + xor_out[47][7][14] + xor_out[48][7][14] + xor_out[49][7][14];
assign sum_out[10][7][14] = xor_out[50][7][14] + xor_out[51][7][14] + xor_out[52][7][14] + xor_out[53][7][14] + xor_out[54][7][14];
assign sum_out[11][7][14] = xor_out[55][7][14] + xor_out[56][7][14] + xor_out[57][7][14] + xor_out[58][7][14] + xor_out[59][7][14];
assign sum_out[12][7][14] = xor_out[60][7][14] + xor_out[61][7][14] + xor_out[62][7][14] + xor_out[63][7][14] + xor_out[64][7][14];
assign sum_out[13][7][14] = xor_out[65][7][14] + xor_out[66][7][14] + xor_out[67][7][14] + xor_out[68][7][14] + xor_out[69][7][14];
assign sum_out[14][7][14] = xor_out[70][7][14] + xor_out[71][7][14] + xor_out[72][7][14] + xor_out[73][7][14] + xor_out[74][7][14];
assign sum_out[15][7][14] = xor_out[75][7][14] + xor_out[76][7][14] + xor_out[77][7][14] + xor_out[78][7][14] + xor_out[79][7][14];
assign sum_out[16][7][14] = xor_out[80][7][14] + xor_out[81][7][14] + xor_out[82][7][14] + xor_out[83][7][14] + xor_out[84][7][14];
assign sum_out[17][7][14] = xor_out[85][7][14] + xor_out[86][7][14] + xor_out[87][7][14] + xor_out[88][7][14] + xor_out[89][7][14];
assign sum_out[18][7][14] = xor_out[90][7][14] + xor_out[91][7][14] + xor_out[92][7][14] + xor_out[93][7][14] + xor_out[94][7][14];
assign sum_out[19][7][14] = xor_out[95][7][14] + xor_out[96][7][14] + xor_out[97][7][14] + xor_out[98][7][14] + xor_out[99][7][14];

assign sum_out[0][7][15] = xor_out[0][7][15] + xor_out[1][7][15] + xor_out[2][7][15] + xor_out[3][7][15] + xor_out[4][7][15];
assign sum_out[1][7][15] = xor_out[5][7][15] + xor_out[6][7][15] + xor_out[7][7][15] + xor_out[8][7][15] + xor_out[9][7][15];
assign sum_out[2][7][15] = xor_out[10][7][15] + xor_out[11][7][15] + xor_out[12][7][15] + xor_out[13][7][15] + xor_out[14][7][15];
assign sum_out[3][7][15] = xor_out[15][7][15] + xor_out[16][7][15] + xor_out[17][7][15] + xor_out[18][7][15] + xor_out[19][7][15];
assign sum_out[4][7][15] = xor_out[20][7][15] + xor_out[21][7][15] + xor_out[22][7][15] + xor_out[23][7][15] + xor_out[24][7][15];
assign sum_out[5][7][15] = xor_out[25][7][15] + xor_out[26][7][15] + xor_out[27][7][15] + xor_out[28][7][15] + xor_out[29][7][15];
assign sum_out[6][7][15] = xor_out[30][7][15] + xor_out[31][7][15] + xor_out[32][7][15] + xor_out[33][7][15] + xor_out[34][7][15];
assign sum_out[7][7][15] = xor_out[35][7][15] + xor_out[36][7][15] + xor_out[37][7][15] + xor_out[38][7][15] + xor_out[39][7][15];
assign sum_out[8][7][15] = xor_out[40][7][15] + xor_out[41][7][15] + xor_out[42][7][15] + xor_out[43][7][15] + xor_out[44][7][15];
assign sum_out[9][7][15] = xor_out[45][7][15] + xor_out[46][7][15] + xor_out[47][7][15] + xor_out[48][7][15] + xor_out[49][7][15];
assign sum_out[10][7][15] = xor_out[50][7][15] + xor_out[51][7][15] + xor_out[52][7][15] + xor_out[53][7][15] + xor_out[54][7][15];
assign sum_out[11][7][15] = xor_out[55][7][15] + xor_out[56][7][15] + xor_out[57][7][15] + xor_out[58][7][15] + xor_out[59][7][15];
assign sum_out[12][7][15] = xor_out[60][7][15] + xor_out[61][7][15] + xor_out[62][7][15] + xor_out[63][7][15] + xor_out[64][7][15];
assign sum_out[13][7][15] = xor_out[65][7][15] + xor_out[66][7][15] + xor_out[67][7][15] + xor_out[68][7][15] + xor_out[69][7][15];
assign sum_out[14][7][15] = xor_out[70][7][15] + xor_out[71][7][15] + xor_out[72][7][15] + xor_out[73][7][15] + xor_out[74][7][15];
assign sum_out[15][7][15] = xor_out[75][7][15] + xor_out[76][7][15] + xor_out[77][7][15] + xor_out[78][7][15] + xor_out[79][7][15];
assign sum_out[16][7][15] = xor_out[80][7][15] + xor_out[81][7][15] + xor_out[82][7][15] + xor_out[83][7][15] + xor_out[84][7][15];
assign sum_out[17][7][15] = xor_out[85][7][15] + xor_out[86][7][15] + xor_out[87][7][15] + xor_out[88][7][15] + xor_out[89][7][15];
assign sum_out[18][7][15] = xor_out[90][7][15] + xor_out[91][7][15] + xor_out[92][7][15] + xor_out[93][7][15] + xor_out[94][7][15];
assign sum_out[19][7][15] = xor_out[95][7][15] + xor_out[96][7][15] + xor_out[97][7][15] + xor_out[98][7][15] + xor_out[99][7][15];

assign sum_out[0][7][16] = xor_out[0][7][16] + xor_out[1][7][16] + xor_out[2][7][16] + xor_out[3][7][16] + xor_out[4][7][16];
assign sum_out[1][7][16] = xor_out[5][7][16] + xor_out[6][7][16] + xor_out[7][7][16] + xor_out[8][7][16] + xor_out[9][7][16];
assign sum_out[2][7][16] = xor_out[10][7][16] + xor_out[11][7][16] + xor_out[12][7][16] + xor_out[13][7][16] + xor_out[14][7][16];
assign sum_out[3][7][16] = xor_out[15][7][16] + xor_out[16][7][16] + xor_out[17][7][16] + xor_out[18][7][16] + xor_out[19][7][16];
assign sum_out[4][7][16] = xor_out[20][7][16] + xor_out[21][7][16] + xor_out[22][7][16] + xor_out[23][7][16] + xor_out[24][7][16];
assign sum_out[5][7][16] = xor_out[25][7][16] + xor_out[26][7][16] + xor_out[27][7][16] + xor_out[28][7][16] + xor_out[29][7][16];
assign sum_out[6][7][16] = xor_out[30][7][16] + xor_out[31][7][16] + xor_out[32][7][16] + xor_out[33][7][16] + xor_out[34][7][16];
assign sum_out[7][7][16] = xor_out[35][7][16] + xor_out[36][7][16] + xor_out[37][7][16] + xor_out[38][7][16] + xor_out[39][7][16];
assign sum_out[8][7][16] = xor_out[40][7][16] + xor_out[41][7][16] + xor_out[42][7][16] + xor_out[43][7][16] + xor_out[44][7][16];
assign sum_out[9][7][16] = xor_out[45][7][16] + xor_out[46][7][16] + xor_out[47][7][16] + xor_out[48][7][16] + xor_out[49][7][16];
assign sum_out[10][7][16] = xor_out[50][7][16] + xor_out[51][7][16] + xor_out[52][7][16] + xor_out[53][7][16] + xor_out[54][7][16];
assign sum_out[11][7][16] = xor_out[55][7][16] + xor_out[56][7][16] + xor_out[57][7][16] + xor_out[58][7][16] + xor_out[59][7][16];
assign sum_out[12][7][16] = xor_out[60][7][16] + xor_out[61][7][16] + xor_out[62][7][16] + xor_out[63][7][16] + xor_out[64][7][16];
assign sum_out[13][7][16] = xor_out[65][7][16] + xor_out[66][7][16] + xor_out[67][7][16] + xor_out[68][7][16] + xor_out[69][7][16];
assign sum_out[14][7][16] = xor_out[70][7][16] + xor_out[71][7][16] + xor_out[72][7][16] + xor_out[73][7][16] + xor_out[74][7][16];
assign sum_out[15][7][16] = xor_out[75][7][16] + xor_out[76][7][16] + xor_out[77][7][16] + xor_out[78][7][16] + xor_out[79][7][16];
assign sum_out[16][7][16] = xor_out[80][7][16] + xor_out[81][7][16] + xor_out[82][7][16] + xor_out[83][7][16] + xor_out[84][7][16];
assign sum_out[17][7][16] = xor_out[85][7][16] + xor_out[86][7][16] + xor_out[87][7][16] + xor_out[88][7][16] + xor_out[89][7][16];
assign sum_out[18][7][16] = xor_out[90][7][16] + xor_out[91][7][16] + xor_out[92][7][16] + xor_out[93][7][16] + xor_out[94][7][16];
assign sum_out[19][7][16] = xor_out[95][7][16] + xor_out[96][7][16] + xor_out[97][7][16] + xor_out[98][7][16] + xor_out[99][7][16];

assign sum_out[0][7][17] = xor_out[0][7][17] + xor_out[1][7][17] + xor_out[2][7][17] + xor_out[3][7][17] + xor_out[4][7][17];
assign sum_out[1][7][17] = xor_out[5][7][17] + xor_out[6][7][17] + xor_out[7][7][17] + xor_out[8][7][17] + xor_out[9][7][17];
assign sum_out[2][7][17] = xor_out[10][7][17] + xor_out[11][7][17] + xor_out[12][7][17] + xor_out[13][7][17] + xor_out[14][7][17];
assign sum_out[3][7][17] = xor_out[15][7][17] + xor_out[16][7][17] + xor_out[17][7][17] + xor_out[18][7][17] + xor_out[19][7][17];
assign sum_out[4][7][17] = xor_out[20][7][17] + xor_out[21][7][17] + xor_out[22][7][17] + xor_out[23][7][17] + xor_out[24][7][17];
assign sum_out[5][7][17] = xor_out[25][7][17] + xor_out[26][7][17] + xor_out[27][7][17] + xor_out[28][7][17] + xor_out[29][7][17];
assign sum_out[6][7][17] = xor_out[30][7][17] + xor_out[31][7][17] + xor_out[32][7][17] + xor_out[33][7][17] + xor_out[34][7][17];
assign sum_out[7][7][17] = xor_out[35][7][17] + xor_out[36][7][17] + xor_out[37][7][17] + xor_out[38][7][17] + xor_out[39][7][17];
assign sum_out[8][7][17] = xor_out[40][7][17] + xor_out[41][7][17] + xor_out[42][7][17] + xor_out[43][7][17] + xor_out[44][7][17];
assign sum_out[9][7][17] = xor_out[45][7][17] + xor_out[46][7][17] + xor_out[47][7][17] + xor_out[48][7][17] + xor_out[49][7][17];
assign sum_out[10][7][17] = xor_out[50][7][17] + xor_out[51][7][17] + xor_out[52][7][17] + xor_out[53][7][17] + xor_out[54][7][17];
assign sum_out[11][7][17] = xor_out[55][7][17] + xor_out[56][7][17] + xor_out[57][7][17] + xor_out[58][7][17] + xor_out[59][7][17];
assign sum_out[12][7][17] = xor_out[60][7][17] + xor_out[61][7][17] + xor_out[62][7][17] + xor_out[63][7][17] + xor_out[64][7][17];
assign sum_out[13][7][17] = xor_out[65][7][17] + xor_out[66][7][17] + xor_out[67][7][17] + xor_out[68][7][17] + xor_out[69][7][17];
assign sum_out[14][7][17] = xor_out[70][7][17] + xor_out[71][7][17] + xor_out[72][7][17] + xor_out[73][7][17] + xor_out[74][7][17];
assign sum_out[15][7][17] = xor_out[75][7][17] + xor_out[76][7][17] + xor_out[77][7][17] + xor_out[78][7][17] + xor_out[79][7][17];
assign sum_out[16][7][17] = xor_out[80][7][17] + xor_out[81][7][17] + xor_out[82][7][17] + xor_out[83][7][17] + xor_out[84][7][17];
assign sum_out[17][7][17] = xor_out[85][7][17] + xor_out[86][7][17] + xor_out[87][7][17] + xor_out[88][7][17] + xor_out[89][7][17];
assign sum_out[18][7][17] = xor_out[90][7][17] + xor_out[91][7][17] + xor_out[92][7][17] + xor_out[93][7][17] + xor_out[94][7][17];
assign sum_out[19][7][17] = xor_out[95][7][17] + xor_out[96][7][17] + xor_out[97][7][17] + xor_out[98][7][17] + xor_out[99][7][17];

assign sum_out[0][7][18] = xor_out[0][7][18] + xor_out[1][7][18] + xor_out[2][7][18] + xor_out[3][7][18] + xor_out[4][7][18];
assign sum_out[1][7][18] = xor_out[5][7][18] + xor_out[6][7][18] + xor_out[7][7][18] + xor_out[8][7][18] + xor_out[9][7][18];
assign sum_out[2][7][18] = xor_out[10][7][18] + xor_out[11][7][18] + xor_out[12][7][18] + xor_out[13][7][18] + xor_out[14][7][18];
assign sum_out[3][7][18] = xor_out[15][7][18] + xor_out[16][7][18] + xor_out[17][7][18] + xor_out[18][7][18] + xor_out[19][7][18];
assign sum_out[4][7][18] = xor_out[20][7][18] + xor_out[21][7][18] + xor_out[22][7][18] + xor_out[23][7][18] + xor_out[24][7][18];
assign sum_out[5][7][18] = xor_out[25][7][18] + xor_out[26][7][18] + xor_out[27][7][18] + xor_out[28][7][18] + xor_out[29][7][18];
assign sum_out[6][7][18] = xor_out[30][7][18] + xor_out[31][7][18] + xor_out[32][7][18] + xor_out[33][7][18] + xor_out[34][7][18];
assign sum_out[7][7][18] = xor_out[35][7][18] + xor_out[36][7][18] + xor_out[37][7][18] + xor_out[38][7][18] + xor_out[39][7][18];
assign sum_out[8][7][18] = xor_out[40][7][18] + xor_out[41][7][18] + xor_out[42][7][18] + xor_out[43][7][18] + xor_out[44][7][18];
assign sum_out[9][7][18] = xor_out[45][7][18] + xor_out[46][7][18] + xor_out[47][7][18] + xor_out[48][7][18] + xor_out[49][7][18];
assign sum_out[10][7][18] = xor_out[50][7][18] + xor_out[51][7][18] + xor_out[52][7][18] + xor_out[53][7][18] + xor_out[54][7][18];
assign sum_out[11][7][18] = xor_out[55][7][18] + xor_out[56][7][18] + xor_out[57][7][18] + xor_out[58][7][18] + xor_out[59][7][18];
assign sum_out[12][7][18] = xor_out[60][7][18] + xor_out[61][7][18] + xor_out[62][7][18] + xor_out[63][7][18] + xor_out[64][7][18];
assign sum_out[13][7][18] = xor_out[65][7][18] + xor_out[66][7][18] + xor_out[67][7][18] + xor_out[68][7][18] + xor_out[69][7][18];
assign sum_out[14][7][18] = xor_out[70][7][18] + xor_out[71][7][18] + xor_out[72][7][18] + xor_out[73][7][18] + xor_out[74][7][18];
assign sum_out[15][7][18] = xor_out[75][7][18] + xor_out[76][7][18] + xor_out[77][7][18] + xor_out[78][7][18] + xor_out[79][7][18];
assign sum_out[16][7][18] = xor_out[80][7][18] + xor_out[81][7][18] + xor_out[82][7][18] + xor_out[83][7][18] + xor_out[84][7][18];
assign sum_out[17][7][18] = xor_out[85][7][18] + xor_out[86][7][18] + xor_out[87][7][18] + xor_out[88][7][18] + xor_out[89][7][18];
assign sum_out[18][7][18] = xor_out[90][7][18] + xor_out[91][7][18] + xor_out[92][7][18] + xor_out[93][7][18] + xor_out[94][7][18];
assign sum_out[19][7][18] = xor_out[95][7][18] + xor_out[96][7][18] + xor_out[97][7][18] + xor_out[98][7][18] + xor_out[99][7][18];

assign sum_out[0][7][19] = xor_out[0][7][19] + xor_out[1][7][19] + xor_out[2][7][19] + xor_out[3][7][19] + xor_out[4][7][19];
assign sum_out[1][7][19] = xor_out[5][7][19] + xor_out[6][7][19] + xor_out[7][7][19] + xor_out[8][7][19] + xor_out[9][7][19];
assign sum_out[2][7][19] = xor_out[10][7][19] + xor_out[11][7][19] + xor_out[12][7][19] + xor_out[13][7][19] + xor_out[14][7][19];
assign sum_out[3][7][19] = xor_out[15][7][19] + xor_out[16][7][19] + xor_out[17][7][19] + xor_out[18][7][19] + xor_out[19][7][19];
assign sum_out[4][7][19] = xor_out[20][7][19] + xor_out[21][7][19] + xor_out[22][7][19] + xor_out[23][7][19] + xor_out[24][7][19];
assign sum_out[5][7][19] = xor_out[25][7][19] + xor_out[26][7][19] + xor_out[27][7][19] + xor_out[28][7][19] + xor_out[29][7][19];
assign sum_out[6][7][19] = xor_out[30][7][19] + xor_out[31][7][19] + xor_out[32][7][19] + xor_out[33][7][19] + xor_out[34][7][19];
assign sum_out[7][7][19] = xor_out[35][7][19] + xor_out[36][7][19] + xor_out[37][7][19] + xor_out[38][7][19] + xor_out[39][7][19];
assign sum_out[8][7][19] = xor_out[40][7][19] + xor_out[41][7][19] + xor_out[42][7][19] + xor_out[43][7][19] + xor_out[44][7][19];
assign sum_out[9][7][19] = xor_out[45][7][19] + xor_out[46][7][19] + xor_out[47][7][19] + xor_out[48][7][19] + xor_out[49][7][19];
assign sum_out[10][7][19] = xor_out[50][7][19] + xor_out[51][7][19] + xor_out[52][7][19] + xor_out[53][7][19] + xor_out[54][7][19];
assign sum_out[11][7][19] = xor_out[55][7][19] + xor_out[56][7][19] + xor_out[57][7][19] + xor_out[58][7][19] + xor_out[59][7][19];
assign sum_out[12][7][19] = xor_out[60][7][19] + xor_out[61][7][19] + xor_out[62][7][19] + xor_out[63][7][19] + xor_out[64][7][19];
assign sum_out[13][7][19] = xor_out[65][7][19] + xor_out[66][7][19] + xor_out[67][7][19] + xor_out[68][7][19] + xor_out[69][7][19];
assign sum_out[14][7][19] = xor_out[70][7][19] + xor_out[71][7][19] + xor_out[72][7][19] + xor_out[73][7][19] + xor_out[74][7][19];
assign sum_out[15][7][19] = xor_out[75][7][19] + xor_out[76][7][19] + xor_out[77][7][19] + xor_out[78][7][19] + xor_out[79][7][19];
assign sum_out[16][7][19] = xor_out[80][7][19] + xor_out[81][7][19] + xor_out[82][7][19] + xor_out[83][7][19] + xor_out[84][7][19];
assign sum_out[17][7][19] = xor_out[85][7][19] + xor_out[86][7][19] + xor_out[87][7][19] + xor_out[88][7][19] + xor_out[89][7][19];
assign sum_out[18][7][19] = xor_out[90][7][19] + xor_out[91][7][19] + xor_out[92][7][19] + xor_out[93][7][19] + xor_out[94][7][19];
assign sum_out[19][7][19] = xor_out[95][7][19] + xor_out[96][7][19] + xor_out[97][7][19] + xor_out[98][7][19] + xor_out[99][7][19];

assign sum_out[0][7][20] = xor_out[0][7][20] + xor_out[1][7][20] + xor_out[2][7][20] + xor_out[3][7][20] + xor_out[4][7][20];
assign sum_out[1][7][20] = xor_out[5][7][20] + xor_out[6][7][20] + xor_out[7][7][20] + xor_out[8][7][20] + xor_out[9][7][20];
assign sum_out[2][7][20] = xor_out[10][7][20] + xor_out[11][7][20] + xor_out[12][7][20] + xor_out[13][7][20] + xor_out[14][7][20];
assign sum_out[3][7][20] = xor_out[15][7][20] + xor_out[16][7][20] + xor_out[17][7][20] + xor_out[18][7][20] + xor_out[19][7][20];
assign sum_out[4][7][20] = xor_out[20][7][20] + xor_out[21][7][20] + xor_out[22][7][20] + xor_out[23][7][20] + xor_out[24][7][20];
assign sum_out[5][7][20] = xor_out[25][7][20] + xor_out[26][7][20] + xor_out[27][7][20] + xor_out[28][7][20] + xor_out[29][7][20];
assign sum_out[6][7][20] = xor_out[30][7][20] + xor_out[31][7][20] + xor_out[32][7][20] + xor_out[33][7][20] + xor_out[34][7][20];
assign sum_out[7][7][20] = xor_out[35][7][20] + xor_out[36][7][20] + xor_out[37][7][20] + xor_out[38][7][20] + xor_out[39][7][20];
assign sum_out[8][7][20] = xor_out[40][7][20] + xor_out[41][7][20] + xor_out[42][7][20] + xor_out[43][7][20] + xor_out[44][7][20];
assign sum_out[9][7][20] = xor_out[45][7][20] + xor_out[46][7][20] + xor_out[47][7][20] + xor_out[48][7][20] + xor_out[49][7][20];
assign sum_out[10][7][20] = xor_out[50][7][20] + xor_out[51][7][20] + xor_out[52][7][20] + xor_out[53][7][20] + xor_out[54][7][20];
assign sum_out[11][7][20] = xor_out[55][7][20] + xor_out[56][7][20] + xor_out[57][7][20] + xor_out[58][7][20] + xor_out[59][7][20];
assign sum_out[12][7][20] = xor_out[60][7][20] + xor_out[61][7][20] + xor_out[62][7][20] + xor_out[63][7][20] + xor_out[64][7][20];
assign sum_out[13][7][20] = xor_out[65][7][20] + xor_out[66][7][20] + xor_out[67][7][20] + xor_out[68][7][20] + xor_out[69][7][20];
assign sum_out[14][7][20] = xor_out[70][7][20] + xor_out[71][7][20] + xor_out[72][7][20] + xor_out[73][7][20] + xor_out[74][7][20];
assign sum_out[15][7][20] = xor_out[75][7][20] + xor_out[76][7][20] + xor_out[77][7][20] + xor_out[78][7][20] + xor_out[79][7][20];
assign sum_out[16][7][20] = xor_out[80][7][20] + xor_out[81][7][20] + xor_out[82][7][20] + xor_out[83][7][20] + xor_out[84][7][20];
assign sum_out[17][7][20] = xor_out[85][7][20] + xor_out[86][7][20] + xor_out[87][7][20] + xor_out[88][7][20] + xor_out[89][7][20];
assign sum_out[18][7][20] = xor_out[90][7][20] + xor_out[91][7][20] + xor_out[92][7][20] + xor_out[93][7][20] + xor_out[94][7][20];
assign sum_out[19][7][20] = xor_out[95][7][20] + xor_out[96][7][20] + xor_out[97][7][20] + xor_out[98][7][20] + xor_out[99][7][20];

assign sum_out[0][7][21] = xor_out[0][7][21] + xor_out[1][7][21] + xor_out[2][7][21] + xor_out[3][7][21] + xor_out[4][7][21];
assign sum_out[1][7][21] = xor_out[5][7][21] + xor_out[6][7][21] + xor_out[7][7][21] + xor_out[8][7][21] + xor_out[9][7][21];
assign sum_out[2][7][21] = xor_out[10][7][21] + xor_out[11][7][21] + xor_out[12][7][21] + xor_out[13][7][21] + xor_out[14][7][21];
assign sum_out[3][7][21] = xor_out[15][7][21] + xor_out[16][7][21] + xor_out[17][7][21] + xor_out[18][7][21] + xor_out[19][7][21];
assign sum_out[4][7][21] = xor_out[20][7][21] + xor_out[21][7][21] + xor_out[22][7][21] + xor_out[23][7][21] + xor_out[24][7][21];
assign sum_out[5][7][21] = xor_out[25][7][21] + xor_out[26][7][21] + xor_out[27][7][21] + xor_out[28][7][21] + xor_out[29][7][21];
assign sum_out[6][7][21] = xor_out[30][7][21] + xor_out[31][7][21] + xor_out[32][7][21] + xor_out[33][7][21] + xor_out[34][7][21];
assign sum_out[7][7][21] = xor_out[35][7][21] + xor_out[36][7][21] + xor_out[37][7][21] + xor_out[38][7][21] + xor_out[39][7][21];
assign sum_out[8][7][21] = xor_out[40][7][21] + xor_out[41][7][21] + xor_out[42][7][21] + xor_out[43][7][21] + xor_out[44][7][21];
assign sum_out[9][7][21] = xor_out[45][7][21] + xor_out[46][7][21] + xor_out[47][7][21] + xor_out[48][7][21] + xor_out[49][7][21];
assign sum_out[10][7][21] = xor_out[50][7][21] + xor_out[51][7][21] + xor_out[52][7][21] + xor_out[53][7][21] + xor_out[54][7][21];
assign sum_out[11][7][21] = xor_out[55][7][21] + xor_out[56][7][21] + xor_out[57][7][21] + xor_out[58][7][21] + xor_out[59][7][21];
assign sum_out[12][7][21] = xor_out[60][7][21] + xor_out[61][7][21] + xor_out[62][7][21] + xor_out[63][7][21] + xor_out[64][7][21];
assign sum_out[13][7][21] = xor_out[65][7][21] + xor_out[66][7][21] + xor_out[67][7][21] + xor_out[68][7][21] + xor_out[69][7][21];
assign sum_out[14][7][21] = xor_out[70][7][21] + xor_out[71][7][21] + xor_out[72][7][21] + xor_out[73][7][21] + xor_out[74][7][21];
assign sum_out[15][7][21] = xor_out[75][7][21] + xor_out[76][7][21] + xor_out[77][7][21] + xor_out[78][7][21] + xor_out[79][7][21];
assign sum_out[16][7][21] = xor_out[80][7][21] + xor_out[81][7][21] + xor_out[82][7][21] + xor_out[83][7][21] + xor_out[84][7][21];
assign sum_out[17][7][21] = xor_out[85][7][21] + xor_out[86][7][21] + xor_out[87][7][21] + xor_out[88][7][21] + xor_out[89][7][21];
assign sum_out[18][7][21] = xor_out[90][7][21] + xor_out[91][7][21] + xor_out[92][7][21] + xor_out[93][7][21] + xor_out[94][7][21];
assign sum_out[19][7][21] = xor_out[95][7][21] + xor_out[96][7][21] + xor_out[97][7][21] + xor_out[98][7][21] + xor_out[99][7][21];

assign sum_out[0][7][22] = xor_out[0][7][22] + xor_out[1][7][22] + xor_out[2][7][22] + xor_out[3][7][22] + xor_out[4][7][22];
assign sum_out[1][7][22] = xor_out[5][7][22] + xor_out[6][7][22] + xor_out[7][7][22] + xor_out[8][7][22] + xor_out[9][7][22];
assign sum_out[2][7][22] = xor_out[10][7][22] + xor_out[11][7][22] + xor_out[12][7][22] + xor_out[13][7][22] + xor_out[14][7][22];
assign sum_out[3][7][22] = xor_out[15][7][22] + xor_out[16][7][22] + xor_out[17][7][22] + xor_out[18][7][22] + xor_out[19][7][22];
assign sum_out[4][7][22] = xor_out[20][7][22] + xor_out[21][7][22] + xor_out[22][7][22] + xor_out[23][7][22] + xor_out[24][7][22];
assign sum_out[5][7][22] = xor_out[25][7][22] + xor_out[26][7][22] + xor_out[27][7][22] + xor_out[28][7][22] + xor_out[29][7][22];
assign sum_out[6][7][22] = xor_out[30][7][22] + xor_out[31][7][22] + xor_out[32][7][22] + xor_out[33][7][22] + xor_out[34][7][22];
assign sum_out[7][7][22] = xor_out[35][7][22] + xor_out[36][7][22] + xor_out[37][7][22] + xor_out[38][7][22] + xor_out[39][7][22];
assign sum_out[8][7][22] = xor_out[40][7][22] + xor_out[41][7][22] + xor_out[42][7][22] + xor_out[43][7][22] + xor_out[44][7][22];
assign sum_out[9][7][22] = xor_out[45][7][22] + xor_out[46][7][22] + xor_out[47][7][22] + xor_out[48][7][22] + xor_out[49][7][22];
assign sum_out[10][7][22] = xor_out[50][7][22] + xor_out[51][7][22] + xor_out[52][7][22] + xor_out[53][7][22] + xor_out[54][7][22];
assign sum_out[11][7][22] = xor_out[55][7][22] + xor_out[56][7][22] + xor_out[57][7][22] + xor_out[58][7][22] + xor_out[59][7][22];
assign sum_out[12][7][22] = xor_out[60][7][22] + xor_out[61][7][22] + xor_out[62][7][22] + xor_out[63][7][22] + xor_out[64][7][22];
assign sum_out[13][7][22] = xor_out[65][7][22] + xor_out[66][7][22] + xor_out[67][7][22] + xor_out[68][7][22] + xor_out[69][7][22];
assign sum_out[14][7][22] = xor_out[70][7][22] + xor_out[71][7][22] + xor_out[72][7][22] + xor_out[73][7][22] + xor_out[74][7][22];
assign sum_out[15][7][22] = xor_out[75][7][22] + xor_out[76][7][22] + xor_out[77][7][22] + xor_out[78][7][22] + xor_out[79][7][22];
assign sum_out[16][7][22] = xor_out[80][7][22] + xor_out[81][7][22] + xor_out[82][7][22] + xor_out[83][7][22] + xor_out[84][7][22];
assign sum_out[17][7][22] = xor_out[85][7][22] + xor_out[86][7][22] + xor_out[87][7][22] + xor_out[88][7][22] + xor_out[89][7][22];
assign sum_out[18][7][22] = xor_out[90][7][22] + xor_out[91][7][22] + xor_out[92][7][22] + xor_out[93][7][22] + xor_out[94][7][22];
assign sum_out[19][7][22] = xor_out[95][7][22] + xor_out[96][7][22] + xor_out[97][7][22] + xor_out[98][7][22] + xor_out[99][7][22];

assign sum_out[0][7][23] = xor_out[0][7][23] + xor_out[1][7][23] + xor_out[2][7][23] + xor_out[3][7][23] + xor_out[4][7][23];
assign sum_out[1][7][23] = xor_out[5][7][23] + xor_out[6][7][23] + xor_out[7][7][23] + xor_out[8][7][23] + xor_out[9][7][23];
assign sum_out[2][7][23] = xor_out[10][7][23] + xor_out[11][7][23] + xor_out[12][7][23] + xor_out[13][7][23] + xor_out[14][7][23];
assign sum_out[3][7][23] = xor_out[15][7][23] + xor_out[16][7][23] + xor_out[17][7][23] + xor_out[18][7][23] + xor_out[19][7][23];
assign sum_out[4][7][23] = xor_out[20][7][23] + xor_out[21][7][23] + xor_out[22][7][23] + xor_out[23][7][23] + xor_out[24][7][23];
assign sum_out[5][7][23] = xor_out[25][7][23] + xor_out[26][7][23] + xor_out[27][7][23] + xor_out[28][7][23] + xor_out[29][7][23];
assign sum_out[6][7][23] = xor_out[30][7][23] + xor_out[31][7][23] + xor_out[32][7][23] + xor_out[33][7][23] + xor_out[34][7][23];
assign sum_out[7][7][23] = xor_out[35][7][23] + xor_out[36][7][23] + xor_out[37][7][23] + xor_out[38][7][23] + xor_out[39][7][23];
assign sum_out[8][7][23] = xor_out[40][7][23] + xor_out[41][7][23] + xor_out[42][7][23] + xor_out[43][7][23] + xor_out[44][7][23];
assign sum_out[9][7][23] = xor_out[45][7][23] + xor_out[46][7][23] + xor_out[47][7][23] + xor_out[48][7][23] + xor_out[49][7][23];
assign sum_out[10][7][23] = xor_out[50][7][23] + xor_out[51][7][23] + xor_out[52][7][23] + xor_out[53][7][23] + xor_out[54][7][23];
assign sum_out[11][7][23] = xor_out[55][7][23] + xor_out[56][7][23] + xor_out[57][7][23] + xor_out[58][7][23] + xor_out[59][7][23];
assign sum_out[12][7][23] = xor_out[60][7][23] + xor_out[61][7][23] + xor_out[62][7][23] + xor_out[63][7][23] + xor_out[64][7][23];
assign sum_out[13][7][23] = xor_out[65][7][23] + xor_out[66][7][23] + xor_out[67][7][23] + xor_out[68][7][23] + xor_out[69][7][23];
assign sum_out[14][7][23] = xor_out[70][7][23] + xor_out[71][7][23] + xor_out[72][7][23] + xor_out[73][7][23] + xor_out[74][7][23];
assign sum_out[15][7][23] = xor_out[75][7][23] + xor_out[76][7][23] + xor_out[77][7][23] + xor_out[78][7][23] + xor_out[79][7][23];
assign sum_out[16][7][23] = xor_out[80][7][23] + xor_out[81][7][23] + xor_out[82][7][23] + xor_out[83][7][23] + xor_out[84][7][23];
assign sum_out[17][7][23] = xor_out[85][7][23] + xor_out[86][7][23] + xor_out[87][7][23] + xor_out[88][7][23] + xor_out[89][7][23];
assign sum_out[18][7][23] = xor_out[90][7][23] + xor_out[91][7][23] + xor_out[92][7][23] + xor_out[93][7][23] + xor_out[94][7][23];
assign sum_out[19][7][23] = xor_out[95][7][23] + xor_out[96][7][23] + xor_out[97][7][23] + xor_out[98][7][23] + xor_out[99][7][23];

assign sum_out[0][8][0] = xor_out[0][8][0] + xor_out[1][8][0] + xor_out[2][8][0] + xor_out[3][8][0] + xor_out[4][8][0];
assign sum_out[1][8][0] = xor_out[5][8][0] + xor_out[6][8][0] + xor_out[7][8][0] + xor_out[8][8][0] + xor_out[9][8][0];
assign sum_out[2][8][0] = xor_out[10][8][0] + xor_out[11][8][0] + xor_out[12][8][0] + xor_out[13][8][0] + xor_out[14][8][0];
assign sum_out[3][8][0] = xor_out[15][8][0] + xor_out[16][8][0] + xor_out[17][8][0] + xor_out[18][8][0] + xor_out[19][8][0];
assign sum_out[4][8][0] = xor_out[20][8][0] + xor_out[21][8][0] + xor_out[22][8][0] + xor_out[23][8][0] + xor_out[24][8][0];
assign sum_out[5][8][0] = xor_out[25][8][0] + xor_out[26][8][0] + xor_out[27][8][0] + xor_out[28][8][0] + xor_out[29][8][0];
assign sum_out[6][8][0] = xor_out[30][8][0] + xor_out[31][8][0] + xor_out[32][8][0] + xor_out[33][8][0] + xor_out[34][8][0];
assign sum_out[7][8][0] = xor_out[35][8][0] + xor_out[36][8][0] + xor_out[37][8][0] + xor_out[38][8][0] + xor_out[39][8][0];
assign sum_out[8][8][0] = xor_out[40][8][0] + xor_out[41][8][0] + xor_out[42][8][0] + xor_out[43][8][0] + xor_out[44][8][0];
assign sum_out[9][8][0] = xor_out[45][8][0] + xor_out[46][8][0] + xor_out[47][8][0] + xor_out[48][8][0] + xor_out[49][8][0];
assign sum_out[10][8][0] = xor_out[50][8][0] + xor_out[51][8][0] + xor_out[52][8][0] + xor_out[53][8][0] + xor_out[54][8][0];
assign sum_out[11][8][0] = xor_out[55][8][0] + xor_out[56][8][0] + xor_out[57][8][0] + xor_out[58][8][0] + xor_out[59][8][0];
assign sum_out[12][8][0] = xor_out[60][8][0] + xor_out[61][8][0] + xor_out[62][8][0] + xor_out[63][8][0] + xor_out[64][8][0];
assign sum_out[13][8][0] = xor_out[65][8][0] + xor_out[66][8][0] + xor_out[67][8][0] + xor_out[68][8][0] + xor_out[69][8][0];
assign sum_out[14][8][0] = xor_out[70][8][0] + xor_out[71][8][0] + xor_out[72][8][0] + xor_out[73][8][0] + xor_out[74][8][0];
assign sum_out[15][8][0] = xor_out[75][8][0] + xor_out[76][8][0] + xor_out[77][8][0] + xor_out[78][8][0] + xor_out[79][8][0];
assign sum_out[16][8][0] = xor_out[80][8][0] + xor_out[81][8][0] + xor_out[82][8][0] + xor_out[83][8][0] + xor_out[84][8][0];
assign sum_out[17][8][0] = xor_out[85][8][0] + xor_out[86][8][0] + xor_out[87][8][0] + xor_out[88][8][0] + xor_out[89][8][0];
assign sum_out[18][8][0] = xor_out[90][8][0] + xor_out[91][8][0] + xor_out[92][8][0] + xor_out[93][8][0] + xor_out[94][8][0];
assign sum_out[19][8][0] = xor_out[95][8][0] + xor_out[96][8][0] + xor_out[97][8][0] + xor_out[98][8][0] + xor_out[99][8][0];

assign sum_out[0][8][1] = xor_out[0][8][1] + xor_out[1][8][1] + xor_out[2][8][1] + xor_out[3][8][1] + xor_out[4][8][1];
assign sum_out[1][8][1] = xor_out[5][8][1] + xor_out[6][8][1] + xor_out[7][8][1] + xor_out[8][8][1] + xor_out[9][8][1];
assign sum_out[2][8][1] = xor_out[10][8][1] + xor_out[11][8][1] + xor_out[12][8][1] + xor_out[13][8][1] + xor_out[14][8][1];
assign sum_out[3][8][1] = xor_out[15][8][1] + xor_out[16][8][1] + xor_out[17][8][1] + xor_out[18][8][1] + xor_out[19][8][1];
assign sum_out[4][8][1] = xor_out[20][8][1] + xor_out[21][8][1] + xor_out[22][8][1] + xor_out[23][8][1] + xor_out[24][8][1];
assign sum_out[5][8][1] = xor_out[25][8][1] + xor_out[26][8][1] + xor_out[27][8][1] + xor_out[28][8][1] + xor_out[29][8][1];
assign sum_out[6][8][1] = xor_out[30][8][1] + xor_out[31][8][1] + xor_out[32][8][1] + xor_out[33][8][1] + xor_out[34][8][1];
assign sum_out[7][8][1] = xor_out[35][8][1] + xor_out[36][8][1] + xor_out[37][8][1] + xor_out[38][8][1] + xor_out[39][8][1];
assign sum_out[8][8][1] = xor_out[40][8][1] + xor_out[41][8][1] + xor_out[42][8][1] + xor_out[43][8][1] + xor_out[44][8][1];
assign sum_out[9][8][1] = xor_out[45][8][1] + xor_out[46][8][1] + xor_out[47][8][1] + xor_out[48][8][1] + xor_out[49][8][1];
assign sum_out[10][8][1] = xor_out[50][8][1] + xor_out[51][8][1] + xor_out[52][8][1] + xor_out[53][8][1] + xor_out[54][8][1];
assign sum_out[11][8][1] = xor_out[55][8][1] + xor_out[56][8][1] + xor_out[57][8][1] + xor_out[58][8][1] + xor_out[59][8][1];
assign sum_out[12][8][1] = xor_out[60][8][1] + xor_out[61][8][1] + xor_out[62][8][1] + xor_out[63][8][1] + xor_out[64][8][1];
assign sum_out[13][8][1] = xor_out[65][8][1] + xor_out[66][8][1] + xor_out[67][8][1] + xor_out[68][8][1] + xor_out[69][8][1];
assign sum_out[14][8][1] = xor_out[70][8][1] + xor_out[71][8][1] + xor_out[72][8][1] + xor_out[73][8][1] + xor_out[74][8][1];
assign sum_out[15][8][1] = xor_out[75][8][1] + xor_out[76][8][1] + xor_out[77][8][1] + xor_out[78][8][1] + xor_out[79][8][1];
assign sum_out[16][8][1] = xor_out[80][8][1] + xor_out[81][8][1] + xor_out[82][8][1] + xor_out[83][8][1] + xor_out[84][8][1];
assign sum_out[17][8][1] = xor_out[85][8][1] + xor_out[86][8][1] + xor_out[87][8][1] + xor_out[88][8][1] + xor_out[89][8][1];
assign sum_out[18][8][1] = xor_out[90][8][1] + xor_out[91][8][1] + xor_out[92][8][1] + xor_out[93][8][1] + xor_out[94][8][1];
assign sum_out[19][8][1] = xor_out[95][8][1] + xor_out[96][8][1] + xor_out[97][8][1] + xor_out[98][8][1] + xor_out[99][8][1];

assign sum_out[0][8][2] = xor_out[0][8][2] + xor_out[1][8][2] + xor_out[2][8][2] + xor_out[3][8][2] + xor_out[4][8][2];
assign sum_out[1][8][2] = xor_out[5][8][2] + xor_out[6][8][2] + xor_out[7][8][2] + xor_out[8][8][2] + xor_out[9][8][2];
assign sum_out[2][8][2] = xor_out[10][8][2] + xor_out[11][8][2] + xor_out[12][8][2] + xor_out[13][8][2] + xor_out[14][8][2];
assign sum_out[3][8][2] = xor_out[15][8][2] + xor_out[16][8][2] + xor_out[17][8][2] + xor_out[18][8][2] + xor_out[19][8][2];
assign sum_out[4][8][2] = xor_out[20][8][2] + xor_out[21][8][2] + xor_out[22][8][2] + xor_out[23][8][2] + xor_out[24][8][2];
assign sum_out[5][8][2] = xor_out[25][8][2] + xor_out[26][8][2] + xor_out[27][8][2] + xor_out[28][8][2] + xor_out[29][8][2];
assign sum_out[6][8][2] = xor_out[30][8][2] + xor_out[31][8][2] + xor_out[32][8][2] + xor_out[33][8][2] + xor_out[34][8][2];
assign sum_out[7][8][2] = xor_out[35][8][2] + xor_out[36][8][2] + xor_out[37][8][2] + xor_out[38][8][2] + xor_out[39][8][2];
assign sum_out[8][8][2] = xor_out[40][8][2] + xor_out[41][8][2] + xor_out[42][8][2] + xor_out[43][8][2] + xor_out[44][8][2];
assign sum_out[9][8][2] = xor_out[45][8][2] + xor_out[46][8][2] + xor_out[47][8][2] + xor_out[48][8][2] + xor_out[49][8][2];
assign sum_out[10][8][2] = xor_out[50][8][2] + xor_out[51][8][2] + xor_out[52][8][2] + xor_out[53][8][2] + xor_out[54][8][2];
assign sum_out[11][8][2] = xor_out[55][8][2] + xor_out[56][8][2] + xor_out[57][8][2] + xor_out[58][8][2] + xor_out[59][8][2];
assign sum_out[12][8][2] = xor_out[60][8][2] + xor_out[61][8][2] + xor_out[62][8][2] + xor_out[63][8][2] + xor_out[64][8][2];
assign sum_out[13][8][2] = xor_out[65][8][2] + xor_out[66][8][2] + xor_out[67][8][2] + xor_out[68][8][2] + xor_out[69][8][2];
assign sum_out[14][8][2] = xor_out[70][8][2] + xor_out[71][8][2] + xor_out[72][8][2] + xor_out[73][8][2] + xor_out[74][8][2];
assign sum_out[15][8][2] = xor_out[75][8][2] + xor_out[76][8][2] + xor_out[77][8][2] + xor_out[78][8][2] + xor_out[79][8][2];
assign sum_out[16][8][2] = xor_out[80][8][2] + xor_out[81][8][2] + xor_out[82][8][2] + xor_out[83][8][2] + xor_out[84][8][2];
assign sum_out[17][8][2] = xor_out[85][8][2] + xor_out[86][8][2] + xor_out[87][8][2] + xor_out[88][8][2] + xor_out[89][8][2];
assign sum_out[18][8][2] = xor_out[90][8][2] + xor_out[91][8][2] + xor_out[92][8][2] + xor_out[93][8][2] + xor_out[94][8][2];
assign sum_out[19][8][2] = xor_out[95][8][2] + xor_out[96][8][2] + xor_out[97][8][2] + xor_out[98][8][2] + xor_out[99][8][2];

assign sum_out[0][8][3] = xor_out[0][8][3] + xor_out[1][8][3] + xor_out[2][8][3] + xor_out[3][8][3] + xor_out[4][8][3];
assign sum_out[1][8][3] = xor_out[5][8][3] + xor_out[6][8][3] + xor_out[7][8][3] + xor_out[8][8][3] + xor_out[9][8][3];
assign sum_out[2][8][3] = xor_out[10][8][3] + xor_out[11][8][3] + xor_out[12][8][3] + xor_out[13][8][3] + xor_out[14][8][3];
assign sum_out[3][8][3] = xor_out[15][8][3] + xor_out[16][8][3] + xor_out[17][8][3] + xor_out[18][8][3] + xor_out[19][8][3];
assign sum_out[4][8][3] = xor_out[20][8][3] + xor_out[21][8][3] + xor_out[22][8][3] + xor_out[23][8][3] + xor_out[24][8][3];
assign sum_out[5][8][3] = xor_out[25][8][3] + xor_out[26][8][3] + xor_out[27][8][3] + xor_out[28][8][3] + xor_out[29][8][3];
assign sum_out[6][8][3] = xor_out[30][8][3] + xor_out[31][8][3] + xor_out[32][8][3] + xor_out[33][8][3] + xor_out[34][8][3];
assign sum_out[7][8][3] = xor_out[35][8][3] + xor_out[36][8][3] + xor_out[37][8][3] + xor_out[38][8][3] + xor_out[39][8][3];
assign sum_out[8][8][3] = xor_out[40][8][3] + xor_out[41][8][3] + xor_out[42][8][3] + xor_out[43][8][3] + xor_out[44][8][3];
assign sum_out[9][8][3] = xor_out[45][8][3] + xor_out[46][8][3] + xor_out[47][8][3] + xor_out[48][8][3] + xor_out[49][8][3];
assign sum_out[10][8][3] = xor_out[50][8][3] + xor_out[51][8][3] + xor_out[52][8][3] + xor_out[53][8][3] + xor_out[54][8][3];
assign sum_out[11][8][3] = xor_out[55][8][3] + xor_out[56][8][3] + xor_out[57][8][3] + xor_out[58][8][3] + xor_out[59][8][3];
assign sum_out[12][8][3] = xor_out[60][8][3] + xor_out[61][8][3] + xor_out[62][8][3] + xor_out[63][8][3] + xor_out[64][8][3];
assign sum_out[13][8][3] = xor_out[65][8][3] + xor_out[66][8][3] + xor_out[67][8][3] + xor_out[68][8][3] + xor_out[69][8][3];
assign sum_out[14][8][3] = xor_out[70][8][3] + xor_out[71][8][3] + xor_out[72][8][3] + xor_out[73][8][3] + xor_out[74][8][3];
assign sum_out[15][8][3] = xor_out[75][8][3] + xor_out[76][8][3] + xor_out[77][8][3] + xor_out[78][8][3] + xor_out[79][8][3];
assign sum_out[16][8][3] = xor_out[80][8][3] + xor_out[81][8][3] + xor_out[82][8][3] + xor_out[83][8][3] + xor_out[84][8][3];
assign sum_out[17][8][3] = xor_out[85][8][3] + xor_out[86][8][3] + xor_out[87][8][3] + xor_out[88][8][3] + xor_out[89][8][3];
assign sum_out[18][8][3] = xor_out[90][8][3] + xor_out[91][8][3] + xor_out[92][8][3] + xor_out[93][8][3] + xor_out[94][8][3];
assign sum_out[19][8][3] = xor_out[95][8][3] + xor_out[96][8][3] + xor_out[97][8][3] + xor_out[98][8][3] + xor_out[99][8][3];

assign sum_out[0][8][4] = xor_out[0][8][4] + xor_out[1][8][4] + xor_out[2][8][4] + xor_out[3][8][4] + xor_out[4][8][4];
assign sum_out[1][8][4] = xor_out[5][8][4] + xor_out[6][8][4] + xor_out[7][8][4] + xor_out[8][8][4] + xor_out[9][8][4];
assign sum_out[2][8][4] = xor_out[10][8][4] + xor_out[11][8][4] + xor_out[12][8][4] + xor_out[13][8][4] + xor_out[14][8][4];
assign sum_out[3][8][4] = xor_out[15][8][4] + xor_out[16][8][4] + xor_out[17][8][4] + xor_out[18][8][4] + xor_out[19][8][4];
assign sum_out[4][8][4] = xor_out[20][8][4] + xor_out[21][8][4] + xor_out[22][8][4] + xor_out[23][8][4] + xor_out[24][8][4];
assign sum_out[5][8][4] = xor_out[25][8][4] + xor_out[26][8][4] + xor_out[27][8][4] + xor_out[28][8][4] + xor_out[29][8][4];
assign sum_out[6][8][4] = xor_out[30][8][4] + xor_out[31][8][4] + xor_out[32][8][4] + xor_out[33][8][4] + xor_out[34][8][4];
assign sum_out[7][8][4] = xor_out[35][8][4] + xor_out[36][8][4] + xor_out[37][8][4] + xor_out[38][8][4] + xor_out[39][8][4];
assign sum_out[8][8][4] = xor_out[40][8][4] + xor_out[41][8][4] + xor_out[42][8][4] + xor_out[43][8][4] + xor_out[44][8][4];
assign sum_out[9][8][4] = xor_out[45][8][4] + xor_out[46][8][4] + xor_out[47][8][4] + xor_out[48][8][4] + xor_out[49][8][4];
assign sum_out[10][8][4] = xor_out[50][8][4] + xor_out[51][8][4] + xor_out[52][8][4] + xor_out[53][8][4] + xor_out[54][8][4];
assign sum_out[11][8][4] = xor_out[55][8][4] + xor_out[56][8][4] + xor_out[57][8][4] + xor_out[58][8][4] + xor_out[59][8][4];
assign sum_out[12][8][4] = xor_out[60][8][4] + xor_out[61][8][4] + xor_out[62][8][4] + xor_out[63][8][4] + xor_out[64][8][4];
assign sum_out[13][8][4] = xor_out[65][8][4] + xor_out[66][8][4] + xor_out[67][8][4] + xor_out[68][8][4] + xor_out[69][8][4];
assign sum_out[14][8][4] = xor_out[70][8][4] + xor_out[71][8][4] + xor_out[72][8][4] + xor_out[73][8][4] + xor_out[74][8][4];
assign sum_out[15][8][4] = xor_out[75][8][4] + xor_out[76][8][4] + xor_out[77][8][4] + xor_out[78][8][4] + xor_out[79][8][4];
assign sum_out[16][8][4] = xor_out[80][8][4] + xor_out[81][8][4] + xor_out[82][8][4] + xor_out[83][8][4] + xor_out[84][8][4];
assign sum_out[17][8][4] = xor_out[85][8][4] + xor_out[86][8][4] + xor_out[87][8][4] + xor_out[88][8][4] + xor_out[89][8][4];
assign sum_out[18][8][4] = xor_out[90][8][4] + xor_out[91][8][4] + xor_out[92][8][4] + xor_out[93][8][4] + xor_out[94][8][4];
assign sum_out[19][8][4] = xor_out[95][8][4] + xor_out[96][8][4] + xor_out[97][8][4] + xor_out[98][8][4] + xor_out[99][8][4];

assign sum_out[0][8][5] = xor_out[0][8][5] + xor_out[1][8][5] + xor_out[2][8][5] + xor_out[3][8][5] + xor_out[4][8][5];
assign sum_out[1][8][5] = xor_out[5][8][5] + xor_out[6][8][5] + xor_out[7][8][5] + xor_out[8][8][5] + xor_out[9][8][5];
assign sum_out[2][8][5] = xor_out[10][8][5] + xor_out[11][8][5] + xor_out[12][8][5] + xor_out[13][8][5] + xor_out[14][8][5];
assign sum_out[3][8][5] = xor_out[15][8][5] + xor_out[16][8][5] + xor_out[17][8][5] + xor_out[18][8][5] + xor_out[19][8][5];
assign sum_out[4][8][5] = xor_out[20][8][5] + xor_out[21][8][5] + xor_out[22][8][5] + xor_out[23][8][5] + xor_out[24][8][5];
assign sum_out[5][8][5] = xor_out[25][8][5] + xor_out[26][8][5] + xor_out[27][8][5] + xor_out[28][8][5] + xor_out[29][8][5];
assign sum_out[6][8][5] = xor_out[30][8][5] + xor_out[31][8][5] + xor_out[32][8][5] + xor_out[33][8][5] + xor_out[34][8][5];
assign sum_out[7][8][5] = xor_out[35][8][5] + xor_out[36][8][5] + xor_out[37][8][5] + xor_out[38][8][5] + xor_out[39][8][5];
assign sum_out[8][8][5] = xor_out[40][8][5] + xor_out[41][8][5] + xor_out[42][8][5] + xor_out[43][8][5] + xor_out[44][8][5];
assign sum_out[9][8][5] = xor_out[45][8][5] + xor_out[46][8][5] + xor_out[47][8][5] + xor_out[48][8][5] + xor_out[49][8][5];
assign sum_out[10][8][5] = xor_out[50][8][5] + xor_out[51][8][5] + xor_out[52][8][5] + xor_out[53][8][5] + xor_out[54][8][5];
assign sum_out[11][8][5] = xor_out[55][8][5] + xor_out[56][8][5] + xor_out[57][8][5] + xor_out[58][8][5] + xor_out[59][8][5];
assign sum_out[12][8][5] = xor_out[60][8][5] + xor_out[61][8][5] + xor_out[62][8][5] + xor_out[63][8][5] + xor_out[64][8][5];
assign sum_out[13][8][5] = xor_out[65][8][5] + xor_out[66][8][5] + xor_out[67][8][5] + xor_out[68][8][5] + xor_out[69][8][5];
assign sum_out[14][8][5] = xor_out[70][8][5] + xor_out[71][8][5] + xor_out[72][8][5] + xor_out[73][8][5] + xor_out[74][8][5];
assign sum_out[15][8][5] = xor_out[75][8][5] + xor_out[76][8][5] + xor_out[77][8][5] + xor_out[78][8][5] + xor_out[79][8][5];
assign sum_out[16][8][5] = xor_out[80][8][5] + xor_out[81][8][5] + xor_out[82][8][5] + xor_out[83][8][5] + xor_out[84][8][5];
assign sum_out[17][8][5] = xor_out[85][8][5] + xor_out[86][8][5] + xor_out[87][8][5] + xor_out[88][8][5] + xor_out[89][8][5];
assign sum_out[18][8][5] = xor_out[90][8][5] + xor_out[91][8][5] + xor_out[92][8][5] + xor_out[93][8][5] + xor_out[94][8][5];
assign sum_out[19][8][5] = xor_out[95][8][5] + xor_out[96][8][5] + xor_out[97][8][5] + xor_out[98][8][5] + xor_out[99][8][5];

assign sum_out[0][8][6] = xor_out[0][8][6] + xor_out[1][8][6] + xor_out[2][8][6] + xor_out[3][8][6] + xor_out[4][8][6];
assign sum_out[1][8][6] = xor_out[5][8][6] + xor_out[6][8][6] + xor_out[7][8][6] + xor_out[8][8][6] + xor_out[9][8][6];
assign sum_out[2][8][6] = xor_out[10][8][6] + xor_out[11][8][6] + xor_out[12][8][6] + xor_out[13][8][6] + xor_out[14][8][6];
assign sum_out[3][8][6] = xor_out[15][8][6] + xor_out[16][8][6] + xor_out[17][8][6] + xor_out[18][8][6] + xor_out[19][8][6];
assign sum_out[4][8][6] = xor_out[20][8][6] + xor_out[21][8][6] + xor_out[22][8][6] + xor_out[23][8][6] + xor_out[24][8][6];
assign sum_out[5][8][6] = xor_out[25][8][6] + xor_out[26][8][6] + xor_out[27][8][6] + xor_out[28][8][6] + xor_out[29][8][6];
assign sum_out[6][8][6] = xor_out[30][8][6] + xor_out[31][8][6] + xor_out[32][8][6] + xor_out[33][8][6] + xor_out[34][8][6];
assign sum_out[7][8][6] = xor_out[35][8][6] + xor_out[36][8][6] + xor_out[37][8][6] + xor_out[38][8][6] + xor_out[39][8][6];
assign sum_out[8][8][6] = xor_out[40][8][6] + xor_out[41][8][6] + xor_out[42][8][6] + xor_out[43][8][6] + xor_out[44][8][6];
assign sum_out[9][8][6] = xor_out[45][8][6] + xor_out[46][8][6] + xor_out[47][8][6] + xor_out[48][8][6] + xor_out[49][8][6];
assign sum_out[10][8][6] = xor_out[50][8][6] + xor_out[51][8][6] + xor_out[52][8][6] + xor_out[53][8][6] + xor_out[54][8][6];
assign sum_out[11][8][6] = xor_out[55][8][6] + xor_out[56][8][6] + xor_out[57][8][6] + xor_out[58][8][6] + xor_out[59][8][6];
assign sum_out[12][8][6] = xor_out[60][8][6] + xor_out[61][8][6] + xor_out[62][8][6] + xor_out[63][8][6] + xor_out[64][8][6];
assign sum_out[13][8][6] = xor_out[65][8][6] + xor_out[66][8][6] + xor_out[67][8][6] + xor_out[68][8][6] + xor_out[69][8][6];
assign sum_out[14][8][6] = xor_out[70][8][6] + xor_out[71][8][6] + xor_out[72][8][6] + xor_out[73][8][6] + xor_out[74][8][6];
assign sum_out[15][8][6] = xor_out[75][8][6] + xor_out[76][8][6] + xor_out[77][8][6] + xor_out[78][8][6] + xor_out[79][8][6];
assign sum_out[16][8][6] = xor_out[80][8][6] + xor_out[81][8][6] + xor_out[82][8][6] + xor_out[83][8][6] + xor_out[84][8][6];
assign sum_out[17][8][6] = xor_out[85][8][6] + xor_out[86][8][6] + xor_out[87][8][6] + xor_out[88][8][6] + xor_out[89][8][6];
assign sum_out[18][8][6] = xor_out[90][8][6] + xor_out[91][8][6] + xor_out[92][8][6] + xor_out[93][8][6] + xor_out[94][8][6];
assign sum_out[19][8][6] = xor_out[95][8][6] + xor_out[96][8][6] + xor_out[97][8][6] + xor_out[98][8][6] + xor_out[99][8][6];

assign sum_out[0][8][7] = xor_out[0][8][7] + xor_out[1][8][7] + xor_out[2][8][7] + xor_out[3][8][7] + xor_out[4][8][7];
assign sum_out[1][8][7] = xor_out[5][8][7] + xor_out[6][8][7] + xor_out[7][8][7] + xor_out[8][8][7] + xor_out[9][8][7];
assign sum_out[2][8][7] = xor_out[10][8][7] + xor_out[11][8][7] + xor_out[12][8][7] + xor_out[13][8][7] + xor_out[14][8][7];
assign sum_out[3][8][7] = xor_out[15][8][7] + xor_out[16][8][7] + xor_out[17][8][7] + xor_out[18][8][7] + xor_out[19][8][7];
assign sum_out[4][8][7] = xor_out[20][8][7] + xor_out[21][8][7] + xor_out[22][8][7] + xor_out[23][8][7] + xor_out[24][8][7];
assign sum_out[5][8][7] = xor_out[25][8][7] + xor_out[26][8][7] + xor_out[27][8][7] + xor_out[28][8][7] + xor_out[29][8][7];
assign sum_out[6][8][7] = xor_out[30][8][7] + xor_out[31][8][7] + xor_out[32][8][7] + xor_out[33][8][7] + xor_out[34][8][7];
assign sum_out[7][8][7] = xor_out[35][8][7] + xor_out[36][8][7] + xor_out[37][8][7] + xor_out[38][8][7] + xor_out[39][8][7];
assign sum_out[8][8][7] = xor_out[40][8][7] + xor_out[41][8][7] + xor_out[42][8][7] + xor_out[43][8][7] + xor_out[44][8][7];
assign sum_out[9][8][7] = xor_out[45][8][7] + xor_out[46][8][7] + xor_out[47][8][7] + xor_out[48][8][7] + xor_out[49][8][7];
assign sum_out[10][8][7] = xor_out[50][8][7] + xor_out[51][8][7] + xor_out[52][8][7] + xor_out[53][8][7] + xor_out[54][8][7];
assign sum_out[11][8][7] = xor_out[55][8][7] + xor_out[56][8][7] + xor_out[57][8][7] + xor_out[58][8][7] + xor_out[59][8][7];
assign sum_out[12][8][7] = xor_out[60][8][7] + xor_out[61][8][7] + xor_out[62][8][7] + xor_out[63][8][7] + xor_out[64][8][7];
assign sum_out[13][8][7] = xor_out[65][8][7] + xor_out[66][8][7] + xor_out[67][8][7] + xor_out[68][8][7] + xor_out[69][8][7];
assign sum_out[14][8][7] = xor_out[70][8][7] + xor_out[71][8][7] + xor_out[72][8][7] + xor_out[73][8][7] + xor_out[74][8][7];
assign sum_out[15][8][7] = xor_out[75][8][7] + xor_out[76][8][7] + xor_out[77][8][7] + xor_out[78][8][7] + xor_out[79][8][7];
assign sum_out[16][8][7] = xor_out[80][8][7] + xor_out[81][8][7] + xor_out[82][8][7] + xor_out[83][8][7] + xor_out[84][8][7];
assign sum_out[17][8][7] = xor_out[85][8][7] + xor_out[86][8][7] + xor_out[87][8][7] + xor_out[88][8][7] + xor_out[89][8][7];
assign sum_out[18][8][7] = xor_out[90][8][7] + xor_out[91][8][7] + xor_out[92][8][7] + xor_out[93][8][7] + xor_out[94][8][7];
assign sum_out[19][8][7] = xor_out[95][8][7] + xor_out[96][8][7] + xor_out[97][8][7] + xor_out[98][8][7] + xor_out[99][8][7];

assign sum_out[0][8][8] = xor_out[0][8][8] + xor_out[1][8][8] + xor_out[2][8][8] + xor_out[3][8][8] + xor_out[4][8][8];
assign sum_out[1][8][8] = xor_out[5][8][8] + xor_out[6][8][8] + xor_out[7][8][8] + xor_out[8][8][8] + xor_out[9][8][8];
assign sum_out[2][8][8] = xor_out[10][8][8] + xor_out[11][8][8] + xor_out[12][8][8] + xor_out[13][8][8] + xor_out[14][8][8];
assign sum_out[3][8][8] = xor_out[15][8][8] + xor_out[16][8][8] + xor_out[17][8][8] + xor_out[18][8][8] + xor_out[19][8][8];
assign sum_out[4][8][8] = xor_out[20][8][8] + xor_out[21][8][8] + xor_out[22][8][8] + xor_out[23][8][8] + xor_out[24][8][8];
assign sum_out[5][8][8] = xor_out[25][8][8] + xor_out[26][8][8] + xor_out[27][8][8] + xor_out[28][8][8] + xor_out[29][8][8];
assign sum_out[6][8][8] = xor_out[30][8][8] + xor_out[31][8][8] + xor_out[32][8][8] + xor_out[33][8][8] + xor_out[34][8][8];
assign sum_out[7][8][8] = xor_out[35][8][8] + xor_out[36][8][8] + xor_out[37][8][8] + xor_out[38][8][8] + xor_out[39][8][8];
assign sum_out[8][8][8] = xor_out[40][8][8] + xor_out[41][8][8] + xor_out[42][8][8] + xor_out[43][8][8] + xor_out[44][8][8];
assign sum_out[9][8][8] = xor_out[45][8][8] + xor_out[46][8][8] + xor_out[47][8][8] + xor_out[48][8][8] + xor_out[49][8][8];
assign sum_out[10][8][8] = xor_out[50][8][8] + xor_out[51][8][8] + xor_out[52][8][8] + xor_out[53][8][8] + xor_out[54][8][8];
assign sum_out[11][8][8] = xor_out[55][8][8] + xor_out[56][8][8] + xor_out[57][8][8] + xor_out[58][8][8] + xor_out[59][8][8];
assign sum_out[12][8][8] = xor_out[60][8][8] + xor_out[61][8][8] + xor_out[62][8][8] + xor_out[63][8][8] + xor_out[64][8][8];
assign sum_out[13][8][8] = xor_out[65][8][8] + xor_out[66][8][8] + xor_out[67][8][8] + xor_out[68][8][8] + xor_out[69][8][8];
assign sum_out[14][8][8] = xor_out[70][8][8] + xor_out[71][8][8] + xor_out[72][8][8] + xor_out[73][8][8] + xor_out[74][8][8];
assign sum_out[15][8][8] = xor_out[75][8][8] + xor_out[76][8][8] + xor_out[77][8][8] + xor_out[78][8][8] + xor_out[79][8][8];
assign sum_out[16][8][8] = xor_out[80][8][8] + xor_out[81][8][8] + xor_out[82][8][8] + xor_out[83][8][8] + xor_out[84][8][8];
assign sum_out[17][8][8] = xor_out[85][8][8] + xor_out[86][8][8] + xor_out[87][8][8] + xor_out[88][8][8] + xor_out[89][8][8];
assign sum_out[18][8][8] = xor_out[90][8][8] + xor_out[91][8][8] + xor_out[92][8][8] + xor_out[93][8][8] + xor_out[94][8][8];
assign sum_out[19][8][8] = xor_out[95][8][8] + xor_out[96][8][8] + xor_out[97][8][8] + xor_out[98][8][8] + xor_out[99][8][8];

assign sum_out[0][8][9] = xor_out[0][8][9] + xor_out[1][8][9] + xor_out[2][8][9] + xor_out[3][8][9] + xor_out[4][8][9];
assign sum_out[1][8][9] = xor_out[5][8][9] + xor_out[6][8][9] + xor_out[7][8][9] + xor_out[8][8][9] + xor_out[9][8][9];
assign sum_out[2][8][9] = xor_out[10][8][9] + xor_out[11][8][9] + xor_out[12][8][9] + xor_out[13][8][9] + xor_out[14][8][9];
assign sum_out[3][8][9] = xor_out[15][8][9] + xor_out[16][8][9] + xor_out[17][8][9] + xor_out[18][8][9] + xor_out[19][8][9];
assign sum_out[4][8][9] = xor_out[20][8][9] + xor_out[21][8][9] + xor_out[22][8][9] + xor_out[23][8][9] + xor_out[24][8][9];
assign sum_out[5][8][9] = xor_out[25][8][9] + xor_out[26][8][9] + xor_out[27][8][9] + xor_out[28][8][9] + xor_out[29][8][9];
assign sum_out[6][8][9] = xor_out[30][8][9] + xor_out[31][8][9] + xor_out[32][8][9] + xor_out[33][8][9] + xor_out[34][8][9];
assign sum_out[7][8][9] = xor_out[35][8][9] + xor_out[36][8][9] + xor_out[37][8][9] + xor_out[38][8][9] + xor_out[39][8][9];
assign sum_out[8][8][9] = xor_out[40][8][9] + xor_out[41][8][9] + xor_out[42][8][9] + xor_out[43][8][9] + xor_out[44][8][9];
assign sum_out[9][8][9] = xor_out[45][8][9] + xor_out[46][8][9] + xor_out[47][8][9] + xor_out[48][8][9] + xor_out[49][8][9];
assign sum_out[10][8][9] = xor_out[50][8][9] + xor_out[51][8][9] + xor_out[52][8][9] + xor_out[53][8][9] + xor_out[54][8][9];
assign sum_out[11][8][9] = xor_out[55][8][9] + xor_out[56][8][9] + xor_out[57][8][9] + xor_out[58][8][9] + xor_out[59][8][9];
assign sum_out[12][8][9] = xor_out[60][8][9] + xor_out[61][8][9] + xor_out[62][8][9] + xor_out[63][8][9] + xor_out[64][8][9];
assign sum_out[13][8][9] = xor_out[65][8][9] + xor_out[66][8][9] + xor_out[67][8][9] + xor_out[68][8][9] + xor_out[69][8][9];
assign sum_out[14][8][9] = xor_out[70][8][9] + xor_out[71][8][9] + xor_out[72][8][9] + xor_out[73][8][9] + xor_out[74][8][9];
assign sum_out[15][8][9] = xor_out[75][8][9] + xor_out[76][8][9] + xor_out[77][8][9] + xor_out[78][8][9] + xor_out[79][8][9];
assign sum_out[16][8][9] = xor_out[80][8][9] + xor_out[81][8][9] + xor_out[82][8][9] + xor_out[83][8][9] + xor_out[84][8][9];
assign sum_out[17][8][9] = xor_out[85][8][9] + xor_out[86][8][9] + xor_out[87][8][9] + xor_out[88][8][9] + xor_out[89][8][9];
assign sum_out[18][8][9] = xor_out[90][8][9] + xor_out[91][8][9] + xor_out[92][8][9] + xor_out[93][8][9] + xor_out[94][8][9];
assign sum_out[19][8][9] = xor_out[95][8][9] + xor_out[96][8][9] + xor_out[97][8][9] + xor_out[98][8][9] + xor_out[99][8][9];

assign sum_out[0][8][10] = xor_out[0][8][10] + xor_out[1][8][10] + xor_out[2][8][10] + xor_out[3][8][10] + xor_out[4][8][10];
assign sum_out[1][8][10] = xor_out[5][8][10] + xor_out[6][8][10] + xor_out[7][8][10] + xor_out[8][8][10] + xor_out[9][8][10];
assign sum_out[2][8][10] = xor_out[10][8][10] + xor_out[11][8][10] + xor_out[12][8][10] + xor_out[13][8][10] + xor_out[14][8][10];
assign sum_out[3][8][10] = xor_out[15][8][10] + xor_out[16][8][10] + xor_out[17][8][10] + xor_out[18][8][10] + xor_out[19][8][10];
assign sum_out[4][8][10] = xor_out[20][8][10] + xor_out[21][8][10] + xor_out[22][8][10] + xor_out[23][8][10] + xor_out[24][8][10];
assign sum_out[5][8][10] = xor_out[25][8][10] + xor_out[26][8][10] + xor_out[27][8][10] + xor_out[28][8][10] + xor_out[29][8][10];
assign sum_out[6][8][10] = xor_out[30][8][10] + xor_out[31][8][10] + xor_out[32][8][10] + xor_out[33][8][10] + xor_out[34][8][10];
assign sum_out[7][8][10] = xor_out[35][8][10] + xor_out[36][8][10] + xor_out[37][8][10] + xor_out[38][8][10] + xor_out[39][8][10];
assign sum_out[8][8][10] = xor_out[40][8][10] + xor_out[41][8][10] + xor_out[42][8][10] + xor_out[43][8][10] + xor_out[44][8][10];
assign sum_out[9][8][10] = xor_out[45][8][10] + xor_out[46][8][10] + xor_out[47][8][10] + xor_out[48][8][10] + xor_out[49][8][10];
assign sum_out[10][8][10] = xor_out[50][8][10] + xor_out[51][8][10] + xor_out[52][8][10] + xor_out[53][8][10] + xor_out[54][8][10];
assign sum_out[11][8][10] = xor_out[55][8][10] + xor_out[56][8][10] + xor_out[57][8][10] + xor_out[58][8][10] + xor_out[59][8][10];
assign sum_out[12][8][10] = xor_out[60][8][10] + xor_out[61][8][10] + xor_out[62][8][10] + xor_out[63][8][10] + xor_out[64][8][10];
assign sum_out[13][8][10] = xor_out[65][8][10] + xor_out[66][8][10] + xor_out[67][8][10] + xor_out[68][8][10] + xor_out[69][8][10];
assign sum_out[14][8][10] = xor_out[70][8][10] + xor_out[71][8][10] + xor_out[72][8][10] + xor_out[73][8][10] + xor_out[74][8][10];
assign sum_out[15][8][10] = xor_out[75][8][10] + xor_out[76][8][10] + xor_out[77][8][10] + xor_out[78][8][10] + xor_out[79][8][10];
assign sum_out[16][8][10] = xor_out[80][8][10] + xor_out[81][8][10] + xor_out[82][8][10] + xor_out[83][8][10] + xor_out[84][8][10];
assign sum_out[17][8][10] = xor_out[85][8][10] + xor_out[86][8][10] + xor_out[87][8][10] + xor_out[88][8][10] + xor_out[89][8][10];
assign sum_out[18][8][10] = xor_out[90][8][10] + xor_out[91][8][10] + xor_out[92][8][10] + xor_out[93][8][10] + xor_out[94][8][10];
assign sum_out[19][8][10] = xor_out[95][8][10] + xor_out[96][8][10] + xor_out[97][8][10] + xor_out[98][8][10] + xor_out[99][8][10];

assign sum_out[0][8][11] = xor_out[0][8][11] + xor_out[1][8][11] + xor_out[2][8][11] + xor_out[3][8][11] + xor_out[4][8][11];
assign sum_out[1][8][11] = xor_out[5][8][11] + xor_out[6][8][11] + xor_out[7][8][11] + xor_out[8][8][11] + xor_out[9][8][11];
assign sum_out[2][8][11] = xor_out[10][8][11] + xor_out[11][8][11] + xor_out[12][8][11] + xor_out[13][8][11] + xor_out[14][8][11];
assign sum_out[3][8][11] = xor_out[15][8][11] + xor_out[16][8][11] + xor_out[17][8][11] + xor_out[18][8][11] + xor_out[19][8][11];
assign sum_out[4][8][11] = xor_out[20][8][11] + xor_out[21][8][11] + xor_out[22][8][11] + xor_out[23][8][11] + xor_out[24][8][11];
assign sum_out[5][8][11] = xor_out[25][8][11] + xor_out[26][8][11] + xor_out[27][8][11] + xor_out[28][8][11] + xor_out[29][8][11];
assign sum_out[6][8][11] = xor_out[30][8][11] + xor_out[31][8][11] + xor_out[32][8][11] + xor_out[33][8][11] + xor_out[34][8][11];
assign sum_out[7][8][11] = xor_out[35][8][11] + xor_out[36][8][11] + xor_out[37][8][11] + xor_out[38][8][11] + xor_out[39][8][11];
assign sum_out[8][8][11] = xor_out[40][8][11] + xor_out[41][8][11] + xor_out[42][8][11] + xor_out[43][8][11] + xor_out[44][8][11];
assign sum_out[9][8][11] = xor_out[45][8][11] + xor_out[46][8][11] + xor_out[47][8][11] + xor_out[48][8][11] + xor_out[49][8][11];
assign sum_out[10][8][11] = xor_out[50][8][11] + xor_out[51][8][11] + xor_out[52][8][11] + xor_out[53][8][11] + xor_out[54][8][11];
assign sum_out[11][8][11] = xor_out[55][8][11] + xor_out[56][8][11] + xor_out[57][8][11] + xor_out[58][8][11] + xor_out[59][8][11];
assign sum_out[12][8][11] = xor_out[60][8][11] + xor_out[61][8][11] + xor_out[62][8][11] + xor_out[63][8][11] + xor_out[64][8][11];
assign sum_out[13][8][11] = xor_out[65][8][11] + xor_out[66][8][11] + xor_out[67][8][11] + xor_out[68][8][11] + xor_out[69][8][11];
assign sum_out[14][8][11] = xor_out[70][8][11] + xor_out[71][8][11] + xor_out[72][8][11] + xor_out[73][8][11] + xor_out[74][8][11];
assign sum_out[15][8][11] = xor_out[75][8][11] + xor_out[76][8][11] + xor_out[77][8][11] + xor_out[78][8][11] + xor_out[79][8][11];
assign sum_out[16][8][11] = xor_out[80][8][11] + xor_out[81][8][11] + xor_out[82][8][11] + xor_out[83][8][11] + xor_out[84][8][11];
assign sum_out[17][8][11] = xor_out[85][8][11] + xor_out[86][8][11] + xor_out[87][8][11] + xor_out[88][8][11] + xor_out[89][8][11];
assign sum_out[18][8][11] = xor_out[90][8][11] + xor_out[91][8][11] + xor_out[92][8][11] + xor_out[93][8][11] + xor_out[94][8][11];
assign sum_out[19][8][11] = xor_out[95][8][11] + xor_out[96][8][11] + xor_out[97][8][11] + xor_out[98][8][11] + xor_out[99][8][11];

assign sum_out[0][8][12] = xor_out[0][8][12] + xor_out[1][8][12] + xor_out[2][8][12] + xor_out[3][8][12] + xor_out[4][8][12];
assign sum_out[1][8][12] = xor_out[5][8][12] + xor_out[6][8][12] + xor_out[7][8][12] + xor_out[8][8][12] + xor_out[9][8][12];
assign sum_out[2][8][12] = xor_out[10][8][12] + xor_out[11][8][12] + xor_out[12][8][12] + xor_out[13][8][12] + xor_out[14][8][12];
assign sum_out[3][8][12] = xor_out[15][8][12] + xor_out[16][8][12] + xor_out[17][8][12] + xor_out[18][8][12] + xor_out[19][8][12];
assign sum_out[4][8][12] = xor_out[20][8][12] + xor_out[21][8][12] + xor_out[22][8][12] + xor_out[23][8][12] + xor_out[24][8][12];
assign sum_out[5][8][12] = xor_out[25][8][12] + xor_out[26][8][12] + xor_out[27][8][12] + xor_out[28][8][12] + xor_out[29][8][12];
assign sum_out[6][8][12] = xor_out[30][8][12] + xor_out[31][8][12] + xor_out[32][8][12] + xor_out[33][8][12] + xor_out[34][8][12];
assign sum_out[7][8][12] = xor_out[35][8][12] + xor_out[36][8][12] + xor_out[37][8][12] + xor_out[38][8][12] + xor_out[39][8][12];
assign sum_out[8][8][12] = xor_out[40][8][12] + xor_out[41][8][12] + xor_out[42][8][12] + xor_out[43][8][12] + xor_out[44][8][12];
assign sum_out[9][8][12] = xor_out[45][8][12] + xor_out[46][8][12] + xor_out[47][8][12] + xor_out[48][8][12] + xor_out[49][8][12];
assign sum_out[10][8][12] = xor_out[50][8][12] + xor_out[51][8][12] + xor_out[52][8][12] + xor_out[53][8][12] + xor_out[54][8][12];
assign sum_out[11][8][12] = xor_out[55][8][12] + xor_out[56][8][12] + xor_out[57][8][12] + xor_out[58][8][12] + xor_out[59][8][12];
assign sum_out[12][8][12] = xor_out[60][8][12] + xor_out[61][8][12] + xor_out[62][8][12] + xor_out[63][8][12] + xor_out[64][8][12];
assign sum_out[13][8][12] = xor_out[65][8][12] + xor_out[66][8][12] + xor_out[67][8][12] + xor_out[68][8][12] + xor_out[69][8][12];
assign sum_out[14][8][12] = xor_out[70][8][12] + xor_out[71][8][12] + xor_out[72][8][12] + xor_out[73][8][12] + xor_out[74][8][12];
assign sum_out[15][8][12] = xor_out[75][8][12] + xor_out[76][8][12] + xor_out[77][8][12] + xor_out[78][8][12] + xor_out[79][8][12];
assign sum_out[16][8][12] = xor_out[80][8][12] + xor_out[81][8][12] + xor_out[82][8][12] + xor_out[83][8][12] + xor_out[84][8][12];
assign sum_out[17][8][12] = xor_out[85][8][12] + xor_out[86][8][12] + xor_out[87][8][12] + xor_out[88][8][12] + xor_out[89][8][12];
assign sum_out[18][8][12] = xor_out[90][8][12] + xor_out[91][8][12] + xor_out[92][8][12] + xor_out[93][8][12] + xor_out[94][8][12];
assign sum_out[19][8][12] = xor_out[95][8][12] + xor_out[96][8][12] + xor_out[97][8][12] + xor_out[98][8][12] + xor_out[99][8][12];

assign sum_out[0][8][13] = xor_out[0][8][13] + xor_out[1][8][13] + xor_out[2][8][13] + xor_out[3][8][13] + xor_out[4][8][13];
assign sum_out[1][8][13] = xor_out[5][8][13] + xor_out[6][8][13] + xor_out[7][8][13] + xor_out[8][8][13] + xor_out[9][8][13];
assign sum_out[2][8][13] = xor_out[10][8][13] + xor_out[11][8][13] + xor_out[12][8][13] + xor_out[13][8][13] + xor_out[14][8][13];
assign sum_out[3][8][13] = xor_out[15][8][13] + xor_out[16][8][13] + xor_out[17][8][13] + xor_out[18][8][13] + xor_out[19][8][13];
assign sum_out[4][8][13] = xor_out[20][8][13] + xor_out[21][8][13] + xor_out[22][8][13] + xor_out[23][8][13] + xor_out[24][8][13];
assign sum_out[5][8][13] = xor_out[25][8][13] + xor_out[26][8][13] + xor_out[27][8][13] + xor_out[28][8][13] + xor_out[29][8][13];
assign sum_out[6][8][13] = xor_out[30][8][13] + xor_out[31][8][13] + xor_out[32][8][13] + xor_out[33][8][13] + xor_out[34][8][13];
assign sum_out[7][8][13] = xor_out[35][8][13] + xor_out[36][8][13] + xor_out[37][8][13] + xor_out[38][8][13] + xor_out[39][8][13];
assign sum_out[8][8][13] = xor_out[40][8][13] + xor_out[41][8][13] + xor_out[42][8][13] + xor_out[43][8][13] + xor_out[44][8][13];
assign sum_out[9][8][13] = xor_out[45][8][13] + xor_out[46][8][13] + xor_out[47][8][13] + xor_out[48][8][13] + xor_out[49][8][13];
assign sum_out[10][8][13] = xor_out[50][8][13] + xor_out[51][8][13] + xor_out[52][8][13] + xor_out[53][8][13] + xor_out[54][8][13];
assign sum_out[11][8][13] = xor_out[55][8][13] + xor_out[56][8][13] + xor_out[57][8][13] + xor_out[58][8][13] + xor_out[59][8][13];
assign sum_out[12][8][13] = xor_out[60][8][13] + xor_out[61][8][13] + xor_out[62][8][13] + xor_out[63][8][13] + xor_out[64][8][13];
assign sum_out[13][8][13] = xor_out[65][8][13] + xor_out[66][8][13] + xor_out[67][8][13] + xor_out[68][8][13] + xor_out[69][8][13];
assign sum_out[14][8][13] = xor_out[70][8][13] + xor_out[71][8][13] + xor_out[72][8][13] + xor_out[73][8][13] + xor_out[74][8][13];
assign sum_out[15][8][13] = xor_out[75][8][13] + xor_out[76][8][13] + xor_out[77][8][13] + xor_out[78][8][13] + xor_out[79][8][13];
assign sum_out[16][8][13] = xor_out[80][8][13] + xor_out[81][8][13] + xor_out[82][8][13] + xor_out[83][8][13] + xor_out[84][8][13];
assign sum_out[17][8][13] = xor_out[85][8][13] + xor_out[86][8][13] + xor_out[87][8][13] + xor_out[88][8][13] + xor_out[89][8][13];
assign sum_out[18][8][13] = xor_out[90][8][13] + xor_out[91][8][13] + xor_out[92][8][13] + xor_out[93][8][13] + xor_out[94][8][13];
assign sum_out[19][8][13] = xor_out[95][8][13] + xor_out[96][8][13] + xor_out[97][8][13] + xor_out[98][8][13] + xor_out[99][8][13];

assign sum_out[0][8][14] = xor_out[0][8][14] + xor_out[1][8][14] + xor_out[2][8][14] + xor_out[3][8][14] + xor_out[4][8][14];
assign sum_out[1][8][14] = xor_out[5][8][14] + xor_out[6][8][14] + xor_out[7][8][14] + xor_out[8][8][14] + xor_out[9][8][14];
assign sum_out[2][8][14] = xor_out[10][8][14] + xor_out[11][8][14] + xor_out[12][8][14] + xor_out[13][8][14] + xor_out[14][8][14];
assign sum_out[3][8][14] = xor_out[15][8][14] + xor_out[16][8][14] + xor_out[17][8][14] + xor_out[18][8][14] + xor_out[19][8][14];
assign sum_out[4][8][14] = xor_out[20][8][14] + xor_out[21][8][14] + xor_out[22][8][14] + xor_out[23][8][14] + xor_out[24][8][14];
assign sum_out[5][8][14] = xor_out[25][8][14] + xor_out[26][8][14] + xor_out[27][8][14] + xor_out[28][8][14] + xor_out[29][8][14];
assign sum_out[6][8][14] = xor_out[30][8][14] + xor_out[31][8][14] + xor_out[32][8][14] + xor_out[33][8][14] + xor_out[34][8][14];
assign sum_out[7][8][14] = xor_out[35][8][14] + xor_out[36][8][14] + xor_out[37][8][14] + xor_out[38][8][14] + xor_out[39][8][14];
assign sum_out[8][8][14] = xor_out[40][8][14] + xor_out[41][8][14] + xor_out[42][8][14] + xor_out[43][8][14] + xor_out[44][8][14];
assign sum_out[9][8][14] = xor_out[45][8][14] + xor_out[46][8][14] + xor_out[47][8][14] + xor_out[48][8][14] + xor_out[49][8][14];
assign sum_out[10][8][14] = xor_out[50][8][14] + xor_out[51][8][14] + xor_out[52][8][14] + xor_out[53][8][14] + xor_out[54][8][14];
assign sum_out[11][8][14] = xor_out[55][8][14] + xor_out[56][8][14] + xor_out[57][8][14] + xor_out[58][8][14] + xor_out[59][8][14];
assign sum_out[12][8][14] = xor_out[60][8][14] + xor_out[61][8][14] + xor_out[62][8][14] + xor_out[63][8][14] + xor_out[64][8][14];
assign sum_out[13][8][14] = xor_out[65][8][14] + xor_out[66][8][14] + xor_out[67][8][14] + xor_out[68][8][14] + xor_out[69][8][14];
assign sum_out[14][8][14] = xor_out[70][8][14] + xor_out[71][8][14] + xor_out[72][8][14] + xor_out[73][8][14] + xor_out[74][8][14];
assign sum_out[15][8][14] = xor_out[75][8][14] + xor_out[76][8][14] + xor_out[77][8][14] + xor_out[78][8][14] + xor_out[79][8][14];
assign sum_out[16][8][14] = xor_out[80][8][14] + xor_out[81][8][14] + xor_out[82][8][14] + xor_out[83][8][14] + xor_out[84][8][14];
assign sum_out[17][8][14] = xor_out[85][8][14] + xor_out[86][8][14] + xor_out[87][8][14] + xor_out[88][8][14] + xor_out[89][8][14];
assign sum_out[18][8][14] = xor_out[90][8][14] + xor_out[91][8][14] + xor_out[92][8][14] + xor_out[93][8][14] + xor_out[94][8][14];
assign sum_out[19][8][14] = xor_out[95][8][14] + xor_out[96][8][14] + xor_out[97][8][14] + xor_out[98][8][14] + xor_out[99][8][14];

assign sum_out[0][8][15] = xor_out[0][8][15] + xor_out[1][8][15] + xor_out[2][8][15] + xor_out[3][8][15] + xor_out[4][8][15];
assign sum_out[1][8][15] = xor_out[5][8][15] + xor_out[6][8][15] + xor_out[7][8][15] + xor_out[8][8][15] + xor_out[9][8][15];
assign sum_out[2][8][15] = xor_out[10][8][15] + xor_out[11][8][15] + xor_out[12][8][15] + xor_out[13][8][15] + xor_out[14][8][15];
assign sum_out[3][8][15] = xor_out[15][8][15] + xor_out[16][8][15] + xor_out[17][8][15] + xor_out[18][8][15] + xor_out[19][8][15];
assign sum_out[4][8][15] = xor_out[20][8][15] + xor_out[21][8][15] + xor_out[22][8][15] + xor_out[23][8][15] + xor_out[24][8][15];
assign sum_out[5][8][15] = xor_out[25][8][15] + xor_out[26][8][15] + xor_out[27][8][15] + xor_out[28][8][15] + xor_out[29][8][15];
assign sum_out[6][8][15] = xor_out[30][8][15] + xor_out[31][8][15] + xor_out[32][8][15] + xor_out[33][8][15] + xor_out[34][8][15];
assign sum_out[7][8][15] = xor_out[35][8][15] + xor_out[36][8][15] + xor_out[37][8][15] + xor_out[38][8][15] + xor_out[39][8][15];
assign sum_out[8][8][15] = xor_out[40][8][15] + xor_out[41][8][15] + xor_out[42][8][15] + xor_out[43][8][15] + xor_out[44][8][15];
assign sum_out[9][8][15] = xor_out[45][8][15] + xor_out[46][8][15] + xor_out[47][8][15] + xor_out[48][8][15] + xor_out[49][8][15];
assign sum_out[10][8][15] = xor_out[50][8][15] + xor_out[51][8][15] + xor_out[52][8][15] + xor_out[53][8][15] + xor_out[54][8][15];
assign sum_out[11][8][15] = xor_out[55][8][15] + xor_out[56][8][15] + xor_out[57][8][15] + xor_out[58][8][15] + xor_out[59][8][15];
assign sum_out[12][8][15] = xor_out[60][8][15] + xor_out[61][8][15] + xor_out[62][8][15] + xor_out[63][8][15] + xor_out[64][8][15];
assign sum_out[13][8][15] = xor_out[65][8][15] + xor_out[66][8][15] + xor_out[67][8][15] + xor_out[68][8][15] + xor_out[69][8][15];
assign sum_out[14][8][15] = xor_out[70][8][15] + xor_out[71][8][15] + xor_out[72][8][15] + xor_out[73][8][15] + xor_out[74][8][15];
assign sum_out[15][8][15] = xor_out[75][8][15] + xor_out[76][8][15] + xor_out[77][8][15] + xor_out[78][8][15] + xor_out[79][8][15];
assign sum_out[16][8][15] = xor_out[80][8][15] + xor_out[81][8][15] + xor_out[82][8][15] + xor_out[83][8][15] + xor_out[84][8][15];
assign sum_out[17][8][15] = xor_out[85][8][15] + xor_out[86][8][15] + xor_out[87][8][15] + xor_out[88][8][15] + xor_out[89][8][15];
assign sum_out[18][8][15] = xor_out[90][8][15] + xor_out[91][8][15] + xor_out[92][8][15] + xor_out[93][8][15] + xor_out[94][8][15];
assign sum_out[19][8][15] = xor_out[95][8][15] + xor_out[96][8][15] + xor_out[97][8][15] + xor_out[98][8][15] + xor_out[99][8][15];

assign sum_out[0][8][16] = xor_out[0][8][16] + xor_out[1][8][16] + xor_out[2][8][16] + xor_out[3][8][16] + xor_out[4][8][16];
assign sum_out[1][8][16] = xor_out[5][8][16] + xor_out[6][8][16] + xor_out[7][8][16] + xor_out[8][8][16] + xor_out[9][8][16];
assign sum_out[2][8][16] = xor_out[10][8][16] + xor_out[11][8][16] + xor_out[12][8][16] + xor_out[13][8][16] + xor_out[14][8][16];
assign sum_out[3][8][16] = xor_out[15][8][16] + xor_out[16][8][16] + xor_out[17][8][16] + xor_out[18][8][16] + xor_out[19][8][16];
assign sum_out[4][8][16] = xor_out[20][8][16] + xor_out[21][8][16] + xor_out[22][8][16] + xor_out[23][8][16] + xor_out[24][8][16];
assign sum_out[5][8][16] = xor_out[25][8][16] + xor_out[26][8][16] + xor_out[27][8][16] + xor_out[28][8][16] + xor_out[29][8][16];
assign sum_out[6][8][16] = xor_out[30][8][16] + xor_out[31][8][16] + xor_out[32][8][16] + xor_out[33][8][16] + xor_out[34][8][16];
assign sum_out[7][8][16] = xor_out[35][8][16] + xor_out[36][8][16] + xor_out[37][8][16] + xor_out[38][8][16] + xor_out[39][8][16];
assign sum_out[8][8][16] = xor_out[40][8][16] + xor_out[41][8][16] + xor_out[42][8][16] + xor_out[43][8][16] + xor_out[44][8][16];
assign sum_out[9][8][16] = xor_out[45][8][16] + xor_out[46][8][16] + xor_out[47][8][16] + xor_out[48][8][16] + xor_out[49][8][16];
assign sum_out[10][8][16] = xor_out[50][8][16] + xor_out[51][8][16] + xor_out[52][8][16] + xor_out[53][8][16] + xor_out[54][8][16];
assign sum_out[11][8][16] = xor_out[55][8][16] + xor_out[56][8][16] + xor_out[57][8][16] + xor_out[58][8][16] + xor_out[59][8][16];
assign sum_out[12][8][16] = xor_out[60][8][16] + xor_out[61][8][16] + xor_out[62][8][16] + xor_out[63][8][16] + xor_out[64][8][16];
assign sum_out[13][8][16] = xor_out[65][8][16] + xor_out[66][8][16] + xor_out[67][8][16] + xor_out[68][8][16] + xor_out[69][8][16];
assign sum_out[14][8][16] = xor_out[70][8][16] + xor_out[71][8][16] + xor_out[72][8][16] + xor_out[73][8][16] + xor_out[74][8][16];
assign sum_out[15][8][16] = xor_out[75][8][16] + xor_out[76][8][16] + xor_out[77][8][16] + xor_out[78][8][16] + xor_out[79][8][16];
assign sum_out[16][8][16] = xor_out[80][8][16] + xor_out[81][8][16] + xor_out[82][8][16] + xor_out[83][8][16] + xor_out[84][8][16];
assign sum_out[17][8][16] = xor_out[85][8][16] + xor_out[86][8][16] + xor_out[87][8][16] + xor_out[88][8][16] + xor_out[89][8][16];
assign sum_out[18][8][16] = xor_out[90][8][16] + xor_out[91][8][16] + xor_out[92][8][16] + xor_out[93][8][16] + xor_out[94][8][16];
assign sum_out[19][8][16] = xor_out[95][8][16] + xor_out[96][8][16] + xor_out[97][8][16] + xor_out[98][8][16] + xor_out[99][8][16];

assign sum_out[0][8][17] = xor_out[0][8][17] + xor_out[1][8][17] + xor_out[2][8][17] + xor_out[3][8][17] + xor_out[4][8][17];
assign sum_out[1][8][17] = xor_out[5][8][17] + xor_out[6][8][17] + xor_out[7][8][17] + xor_out[8][8][17] + xor_out[9][8][17];
assign sum_out[2][8][17] = xor_out[10][8][17] + xor_out[11][8][17] + xor_out[12][8][17] + xor_out[13][8][17] + xor_out[14][8][17];
assign sum_out[3][8][17] = xor_out[15][8][17] + xor_out[16][8][17] + xor_out[17][8][17] + xor_out[18][8][17] + xor_out[19][8][17];
assign sum_out[4][8][17] = xor_out[20][8][17] + xor_out[21][8][17] + xor_out[22][8][17] + xor_out[23][8][17] + xor_out[24][8][17];
assign sum_out[5][8][17] = xor_out[25][8][17] + xor_out[26][8][17] + xor_out[27][8][17] + xor_out[28][8][17] + xor_out[29][8][17];
assign sum_out[6][8][17] = xor_out[30][8][17] + xor_out[31][8][17] + xor_out[32][8][17] + xor_out[33][8][17] + xor_out[34][8][17];
assign sum_out[7][8][17] = xor_out[35][8][17] + xor_out[36][8][17] + xor_out[37][8][17] + xor_out[38][8][17] + xor_out[39][8][17];
assign sum_out[8][8][17] = xor_out[40][8][17] + xor_out[41][8][17] + xor_out[42][8][17] + xor_out[43][8][17] + xor_out[44][8][17];
assign sum_out[9][8][17] = xor_out[45][8][17] + xor_out[46][8][17] + xor_out[47][8][17] + xor_out[48][8][17] + xor_out[49][8][17];
assign sum_out[10][8][17] = xor_out[50][8][17] + xor_out[51][8][17] + xor_out[52][8][17] + xor_out[53][8][17] + xor_out[54][8][17];
assign sum_out[11][8][17] = xor_out[55][8][17] + xor_out[56][8][17] + xor_out[57][8][17] + xor_out[58][8][17] + xor_out[59][8][17];
assign sum_out[12][8][17] = xor_out[60][8][17] + xor_out[61][8][17] + xor_out[62][8][17] + xor_out[63][8][17] + xor_out[64][8][17];
assign sum_out[13][8][17] = xor_out[65][8][17] + xor_out[66][8][17] + xor_out[67][8][17] + xor_out[68][8][17] + xor_out[69][8][17];
assign sum_out[14][8][17] = xor_out[70][8][17] + xor_out[71][8][17] + xor_out[72][8][17] + xor_out[73][8][17] + xor_out[74][8][17];
assign sum_out[15][8][17] = xor_out[75][8][17] + xor_out[76][8][17] + xor_out[77][8][17] + xor_out[78][8][17] + xor_out[79][8][17];
assign sum_out[16][8][17] = xor_out[80][8][17] + xor_out[81][8][17] + xor_out[82][8][17] + xor_out[83][8][17] + xor_out[84][8][17];
assign sum_out[17][8][17] = xor_out[85][8][17] + xor_out[86][8][17] + xor_out[87][8][17] + xor_out[88][8][17] + xor_out[89][8][17];
assign sum_out[18][8][17] = xor_out[90][8][17] + xor_out[91][8][17] + xor_out[92][8][17] + xor_out[93][8][17] + xor_out[94][8][17];
assign sum_out[19][8][17] = xor_out[95][8][17] + xor_out[96][8][17] + xor_out[97][8][17] + xor_out[98][8][17] + xor_out[99][8][17];

assign sum_out[0][8][18] = xor_out[0][8][18] + xor_out[1][8][18] + xor_out[2][8][18] + xor_out[3][8][18] + xor_out[4][8][18];
assign sum_out[1][8][18] = xor_out[5][8][18] + xor_out[6][8][18] + xor_out[7][8][18] + xor_out[8][8][18] + xor_out[9][8][18];
assign sum_out[2][8][18] = xor_out[10][8][18] + xor_out[11][8][18] + xor_out[12][8][18] + xor_out[13][8][18] + xor_out[14][8][18];
assign sum_out[3][8][18] = xor_out[15][8][18] + xor_out[16][8][18] + xor_out[17][8][18] + xor_out[18][8][18] + xor_out[19][8][18];
assign sum_out[4][8][18] = xor_out[20][8][18] + xor_out[21][8][18] + xor_out[22][8][18] + xor_out[23][8][18] + xor_out[24][8][18];
assign sum_out[5][8][18] = xor_out[25][8][18] + xor_out[26][8][18] + xor_out[27][8][18] + xor_out[28][8][18] + xor_out[29][8][18];
assign sum_out[6][8][18] = xor_out[30][8][18] + xor_out[31][8][18] + xor_out[32][8][18] + xor_out[33][8][18] + xor_out[34][8][18];
assign sum_out[7][8][18] = xor_out[35][8][18] + xor_out[36][8][18] + xor_out[37][8][18] + xor_out[38][8][18] + xor_out[39][8][18];
assign sum_out[8][8][18] = xor_out[40][8][18] + xor_out[41][8][18] + xor_out[42][8][18] + xor_out[43][8][18] + xor_out[44][8][18];
assign sum_out[9][8][18] = xor_out[45][8][18] + xor_out[46][8][18] + xor_out[47][8][18] + xor_out[48][8][18] + xor_out[49][8][18];
assign sum_out[10][8][18] = xor_out[50][8][18] + xor_out[51][8][18] + xor_out[52][8][18] + xor_out[53][8][18] + xor_out[54][8][18];
assign sum_out[11][8][18] = xor_out[55][8][18] + xor_out[56][8][18] + xor_out[57][8][18] + xor_out[58][8][18] + xor_out[59][8][18];
assign sum_out[12][8][18] = xor_out[60][8][18] + xor_out[61][8][18] + xor_out[62][8][18] + xor_out[63][8][18] + xor_out[64][8][18];
assign sum_out[13][8][18] = xor_out[65][8][18] + xor_out[66][8][18] + xor_out[67][8][18] + xor_out[68][8][18] + xor_out[69][8][18];
assign sum_out[14][8][18] = xor_out[70][8][18] + xor_out[71][8][18] + xor_out[72][8][18] + xor_out[73][8][18] + xor_out[74][8][18];
assign sum_out[15][8][18] = xor_out[75][8][18] + xor_out[76][8][18] + xor_out[77][8][18] + xor_out[78][8][18] + xor_out[79][8][18];
assign sum_out[16][8][18] = xor_out[80][8][18] + xor_out[81][8][18] + xor_out[82][8][18] + xor_out[83][8][18] + xor_out[84][8][18];
assign sum_out[17][8][18] = xor_out[85][8][18] + xor_out[86][8][18] + xor_out[87][8][18] + xor_out[88][8][18] + xor_out[89][8][18];
assign sum_out[18][8][18] = xor_out[90][8][18] + xor_out[91][8][18] + xor_out[92][8][18] + xor_out[93][8][18] + xor_out[94][8][18];
assign sum_out[19][8][18] = xor_out[95][8][18] + xor_out[96][8][18] + xor_out[97][8][18] + xor_out[98][8][18] + xor_out[99][8][18];

assign sum_out[0][8][19] = xor_out[0][8][19] + xor_out[1][8][19] + xor_out[2][8][19] + xor_out[3][8][19] + xor_out[4][8][19];
assign sum_out[1][8][19] = xor_out[5][8][19] + xor_out[6][8][19] + xor_out[7][8][19] + xor_out[8][8][19] + xor_out[9][8][19];
assign sum_out[2][8][19] = xor_out[10][8][19] + xor_out[11][8][19] + xor_out[12][8][19] + xor_out[13][8][19] + xor_out[14][8][19];
assign sum_out[3][8][19] = xor_out[15][8][19] + xor_out[16][8][19] + xor_out[17][8][19] + xor_out[18][8][19] + xor_out[19][8][19];
assign sum_out[4][8][19] = xor_out[20][8][19] + xor_out[21][8][19] + xor_out[22][8][19] + xor_out[23][8][19] + xor_out[24][8][19];
assign sum_out[5][8][19] = xor_out[25][8][19] + xor_out[26][8][19] + xor_out[27][8][19] + xor_out[28][8][19] + xor_out[29][8][19];
assign sum_out[6][8][19] = xor_out[30][8][19] + xor_out[31][8][19] + xor_out[32][8][19] + xor_out[33][8][19] + xor_out[34][8][19];
assign sum_out[7][8][19] = xor_out[35][8][19] + xor_out[36][8][19] + xor_out[37][8][19] + xor_out[38][8][19] + xor_out[39][8][19];
assign sum_out[8][8][19] = xor_out[40][8][19] + xor_out[41][8][19] + xor_out[42][8][19] + xor_out[43][8][19] + xor_out[44][8][19];
assign sum_out[9][8][19] = xor_out[45][8][19] + xor_out[46][8][19] + xor_out[47][8][19] + xor_out[48][8][19] + xor_out[49][8][19];
assign sum_out[10][8][19] = xor_out[50][8][19] + xor_out[51][8][19] + xor_out[52][8][19] + xor_out[53][8][19] + xor_out[54][8][19];
assign sum_out[11][8][19] = xor_out[55][8][19] + xor_out[56][8][19] + xor_out[57][8][19] + xor_out[58][8][19] + xor_out[59][8][19];
assign sum_out[12][8][19] = xor_out[60][8][19] + xor_out[61][8][19] + xor_out[62][8][19] + xor_out[63][8][19] + xor_out[64][8][19];
assign sum_out[13][8][19] = xor_out[65][8][19] + xor_out[66][8][19] + xor_out[67][8][19] + xor_out[68][8][19] + xor_out[69][8][19];
assign sum_out[14][8][19] = xor_out[70][8][19] + xor_out[71][8][19] + xor_out[72][8][19] + xor_out[73][8][19] + xor_out[74][8][19];
assign sum_out[15][8][19] = xor_out[75][8][19] + xor_out[76][8][19] + xor_out[77][8][19] + xor_out[78][8][19] + xor_out[79][8][19];
assign sum_out[16][8][19] = xor_out[80][8][19] + xor_out[81][8][19] + xor_out[82][8][19] + xor_out[83][8][19] + xor_out[84][8][19];
assign sum_out[17][8][19] = xor_out[85][8][19] + xor_out[86][8][19] + xor_out[87][8][19] + xor_out[88][8][19] + xor_out[89][8][19];
assign sum_out[18][8][19] = xor_out[90][8][19] + xor_out[91][8][19] + xor_out[92][8][19] + xor_out[93][8][19] + xor_out[94][8][19];
assign sum_out[19][8][19] = xor_out[95][8][19] + xor_out[96][8][19] + xor_out[97][8][19] + xor_out[98][8][19] + xor_out[99][8][19];

assign sum_out[0][8][20] = xor_out[0][8][20] + xor_out[1][8][20] + xor_out[2][8][20] + xor_out[3][8][20] + xor_out[4][8][20];
assign sum_out[1][8][20] = xor_out[5][8][20] + xor_out[6][8][20] + xor_out[7][8][20] + xor_out[8][8][20] + xor_out[9][8][20];
assign sum_out[2][8][20] = xor_out[10][8][20] + xor_out[11][8][20] + xor_out[12][8][20] + xor_out[13][8][20] + xor_out[14][8][20];
assign sum_out[3][8][20] = xor_out[15][8][20] + xor_out[16][8][20] + xor_out[17][8][20] + xor_out[18][8][20] + xor_out[19][8][20];
assign sum_out[4][8][20] = xor_out[20][8][20] + xor_out[21][8][20] + xor_out[22][8][20] + xor_out[23][8][20] + xor_out[24][8][20];
assign sum_out[5][8][20] = xor_out[25][8][20] + xor_out[26][8][20] + xor_out[27][8][20] + xor_out[28][8][20] + xor_out[29][8][20];
assign sum_out[6][8][20] = xor_out[30][8][20] + xor_out[31][8][20] + xor_out[32][8][20] + xor_out[33][8][20] + xor_out[34][8][20];
assign sum_out[7][8][20] = xor_out[35][8][20] + xor_out[36][8][20] + xor_out[37][8][20] + xor_out[38][8][20] + xor_out[39][8][20];
assign sum_out[8][8][20] = xor_out[40][8][20] + xor_out[41][8][20] + xor_out[42][8][20] + xor_out[43][8][20] + xor_out[44][8][20];
assign sum_out[9][8][20] = xor_out[45][8][20] + xor_out[46][8][20] + xor_out[47][8][20] + xor_out[48][8][20] + xor_out[49][8][20];
assign sum_out[10][8][20] = xor_out[50][8][20] + xor_out[51][8][20] + xor_out[52][8][20] + xor_out[53][8][20] + xor_out[54][8][20];
assign sum_out[11][8][20] = xor_out[55][8][20] + xor_out[56][8][20] + xor_out[57][8][20] + xor_out[58][8][20] + xor_out[59][8][20];
assign sum_out[12][8][20] = xor_out[60][8][20] + xor_out[61][8][20] + xor_out[62][8][20] + xor_out[63][8][20] + xor_out[64][8][20];
assign sum_out[13][8][20] = xor_out[65][8][20] + xor_out[66][8][20] + xor_out[67][8][20] + xor_out[68][8][20] + xor_out[69][8][20];
assign sum_out[14][8][20] = xor_out[70][8][20] + xor_out[71][8][20] + xor_out[72][8][20] + xor_out[73][8][20] + xor_out[74][8][20];
assign sum_out[15][8][20] = xor_out[75][8][20] + xor_out[76][8][20] + xor_out[77][8][20] + xor_out[78][8][20] + xor_out[79][8][20];
assign sum_out[16][8][20] = xor_out[80][8][20] + xor_out[81][8][20] + xor_out[82][8][20] + xor_out[83][8][20] + xor_out[84][8][20];
assign sum_out[17][8][20] = xor_out[85][8][20] + xor_out[86][8][20] + xor_out[87][8][20] + xor_out[88][8][20] + xor_out[89][8][20];
assign sum_out[18][8][20] = xor_out[90][8][20] + xor_out[91][8][20] + xor_out[92][8][20] + xor_out[93][8][20] + xor_out[94][8][20];
assign sum_out[19][8][20] = xor_out[95][8][20] + xor_out[96][8][20] + xor_out[97][8][20] + xor_out[98][8][20] + xor_out[99][8][20];

assign sum_out[0][8][21] = xor_out[0][8][21] + xor_out[1][8][21] + xor_out[2][8][21] + xor_out[3][8][21] + xor_out[4][8][21];
assign sum_out[1][8][21] = xor_out[5][8][21] + xor_out[6][8][21] + xor_out[7][8][21] + xor_out[8][8][21] + xor_out[9][8][21];
assign sum_out[2][8][21] = xor_out[10][8][21] + xor_out[11][8][21] + xor_out[12][8][21] + xor_out[13][8][21] + xor_out[14][8][21];
assign sum_out[3][8][21] = xor_out[15][8][21] + xor_out[16][8][21] + xor_out[17][8][21] + xor_out[18][8][21] + xor_out[19][8][21];
assign sum_out[4][8][21] = xor_out[20][8][21] + xor_out[21][8][21] + xor_out[22][8][21] + xor_out[23][8][21] + xor_out[24][8][21];
assign sum_out[5][8][21] = xor_out[25][8][21] + xor_out[26][8][21] + xor_out[27][8][21] + xor_out[28][8][21] + xor_out[29][8][21];
assign sum_out[6][8][21] = xor_out[30][8][21] + xor_out[31][8][21] + xor_out[32][8][21] + xor_out[33][8][21] + xor_out[34][8][21];
assign sum_out[7][8][21] = xor_out[35][8][21] + xor_out[36][8][21] + xor_out[37][8][21] + xor_out[38][8][21] + xor_out[39][8][21];
assign sum_out[8][8][21] = xor_out[40][8][21] + xor_out[41][8][21] + xor_out[42][8][21] + xor_out[43][8][21] + xor_out[44][8][21];
assign sum_out[9][8][21] = xor_out[45][8][21] + xor_out[46][8][21] + xor_out[47][8][21] + xor_out[48][8][21] + xor_out[49][8][21];
assign sum_out[10][8][21] = xor_out[50][8][21] + xor_out[51][8][21] + xor_out[52][8][21] + xor_out[53][8][21] + xor_out[54][8][21];
assign sum_out[11][8][21] = xor_out[55][8][21] + xor_out[56][8][21] + xor_out[57][8][21] + xor_out[58][8][21] + xor_out[59][8][21];
assign sum_out[12][8][21] = xor_out[60][8][21] + xor_out[61][8][21] + xor_out[62][8][21] + xor_out[63][8][21] + xor_out[64][8][21];
assign sum_out[13][8][21] = xor_out[65][8][21] + xor_out[66][8][21] + xor_out[67][8][21] + xor_out[68][8][21] + xor_out[69][8][21];
assign sum_out[14][8][21] = xor_out[70][8][21] + xor_out[71][8][21] + xor_out[72][8][21] + xor_out[73][8][21] + xor_out[74][8][21];
assign sum_out[15][8][21] = xor_out[75][8][21] + xor_out[76][8][21] + xor_out[77][8][21] + xor_out[78][8][21] + xor_out[79][8][21];
assign sum_out[16][8][21] = xor_out[80][8][21] + xor_out[81][8][21] + xor_out[82][8][21] + xor_out[83][8][21] + xor_out[84][8][21];
assign sum_out[17][8][21] = xor_out[85][8][21] + xor_out[86][8][21] + xor_out[87][8][21] + xor_out[88][8][21] + xor_out[89][8][21];
assign sum_out[18][8][21] = xor_out[90][8][21] + xor_out[91][8][21] + xor_out[92][8][21] + xor_out[93][8][21] + xor_out[94][8][21];
assign sum_out[19][8][21] = xor_out[95][8][21] + xor_out[96][8][21] + xor_out[97][8][21] + xor_out[98][8][21] + xor_out[99][8][21];

assign sum_out[0][8][22] = xor_out[0][8][22] + xor_out[1][8][22] + xor_out[2][8][22] + xor_out[3][8][22] + xor_out[4][8][22];
assign sum_out[1][8][22] = xor_out[5][8][22] + xor_out[6][8][22] + xor_out[7][8][22] + xor_out[8][8][22] + xor_out[9][8][22];
assign sum_out[2][8][22] = xor_out[10][8][22] + xor_out[11][8][22] + xor_out[12][8][22] + xor_out[13][8][22] + xor_out[14][8][22];
assign sum_out[3][8][22] = xor_out[15][8][22] + xor_out[16][8][22] + xor_out[17][8][22] + xor_out[18][8][22] + xor_out[19][8][22];
assign sum_out[4][8][22] = xor_out[20][8][22] + xor_out[21][8][22] + xor_out[22][8][22] + xor_out[23][8][22] + xor_out[24][8][22];
assign sum_out[5][8][22] = xor_out[25][8][22] + xor_out[26][8][22] + xor_out[27][8][22] + xor_out[28][8][22] + xor_out[29][8][22];
assign sum_out[6][8][22] = xor_out[30][8][22] + xor_out[31][8][22] + xor_out[32][8][22] + xor_out[33][8][22] + xor_out[34][8][22];
assign sum_out[7][8][22] = xor_out[35][8][22] + xor_out[36][8][22] + xor_out[37][8][22] + xor_out[38][8][22] + xor_out[39][8][22];
assign sum_out[8][8][22] = xor_out[40][8][22] + xor_out[41][8][22] + xor_out[42][8][22] + xor_out[43][8][22] + xor_out[44][8][22];
assign sum_out[9][8][22] = xor_out[45][8][22] + xor_out[46][8][22] + xor_out[47][8][22] + xor_out[48][8][22] + xor_out[49][8][22];
assign sum_out[10][8][22] = xor_out[50][8][22] + xor_out[51][8][22] + xor_out[52][8][22] + xor_out[53][8][22] + xor_out[54][8][22];
assign sum_out[11][8][22] = xor_out[55][8][22] + xor_out[56][8][22] + xor_out[57][8][22] + xor_out[58][8][22] + xor_out[59][8][22];
assign sum_out[12][8][22] = xor_out[60][8][22] + xor_out[61][8][22] + xor_out[62][8][22] + xor_out[63][8][22] + xor_out[64][8][22];
assign sum_out[13][8][22] = xor_out[65][8][22] + xor_out[66][8][22] + xor_out[67][8][22] + xor_out[68][8][22] + xor_out[69][8][22];
assign sum_out[14][8][22] = xor_out[70][8][22] + xor_out[71][8][22] + xor_out[72][8][22] + xor_out[73][8][22] + xor_out[74][8][22];
assign sum_out[15][8][22] = xor_out[75][8][22] + xor_out[76][8][22] + xor_out[77][8][22] + xor_out[78][8][22] + xor_out[79][8][22];
assign sum_out[16][8][22] = xor_out[80][8][22] + xor_out[81][8][22] + xor_out[82][8][22] + xor_out[83][8][22] + xor_out[84][8][22];
assign sum_out[17][8][22] = xor_out[85][8][22] + xor_out[86][8][22] + xor_out[87][8][22] + xor_out[88][8][22] + xor_out[89][8][22];
assign sum_out[18][8][22] = xor_out[90][8][22] + xor_out[91][8][22] + xor_out[92][8][22] + xor_out[93][8][22] + xor_out[94][8][22];
assign sum_out[19][8][22] = xor_out[95][8][22] + xor_out[96][8][22] + xor_out[97][8][22] + xor_out[98][8][22] + xor_out[99][8][22];

assign sum_out[0][8][23] = xor_out[0][8][23] + xor_out[1][8][23] + xor_out[2][8][23] + xor_out[3][8][23] + xor_out[4][8][23];
assign sum_out[1][8][23] = xor_out[5][8][23] + xor_out[6][8][23] + xor_out[7][8][23] + xor_out[8][8][23] + xor_out[9][8][23];
assign sum_out[2][8][23] = xor_out[10][8][23] + xor_out[11][8][23] + xor_out[12][8][23] + xor_out[13][8][23] + xor_out[14][8][23];
assign sum_out[3][8][23] = xor_out[15][8][23] + xor_out[16][8][23] + xor_out[17][8][23] + xor_out[18][8][23] + xor_out[19][8][23];
assign sum_out[4][8][23] = xor_out[20][8][23] + xor_out[21][8][23] + xor_out[22][8][23] + xor_out[23][8][23] + xor_out[24][8][23];
assign sum_out[5][8][23] = xor_out[25][8][23] + xor_out[26][8][23] + xor_out[27][8][23] + xor_out[28][8][23] + xor_out[29][8][23];
assign sum_out[6][8][23] = xor_out[30][8][23] + xor_out[31][8][23] + xor_out[32][8][23] + xor_out[33][8][23] + xor_out[34][8][23];
assign sum_out[7][8][23] = xor_out[35][8][23] + xor_out[36][8][23] + xor_out[37][8][23] + xor_out[38][8][23] + xor_out[39][8][23];
assign sum_out[8][8][23] = xor_out[40][8][23] + xor_out[41][8][23] + xor_out[42][8][23] + xor_out[43][8][23] + xor_out[44][8][23];
assign sum_out[9][8][23] = xor_out[45][8][23] + xor_out[46][8][23] + xor_out[47][8][23] + xor_out[48][8][23] + xor_out[49][8][23];
assign sum_out[10][8][23] = xor_out[50][8][23] + xor_out[51][8][23] + xor_out[52][8][23] + xor_out[53][8][23] + xor_out[54][8][23];
assign sum_out[11][8][23] = xor_out[55][8][23] + xor_out[56][8][23] + xor_out[57][8][23] + xor_out[58][8][23] + xor_out[59][8][23];
assign sum_out[12][8][23] = xor_out[60][8][23] + xor_out[61][8][23] + xor_out[62][8][23] + xor_out[63][8][23] + xor_out[64][8][23];
assign sum_out[13][8][23] = xor_out[65][8][23] + xor_out[66][8][23] + xor_out[67][8][23] + xor_out[68][8][23] + xor_out[69][8][23];
assign sum_out[14][8][23] = xor_out[70][8][23] + xor_out[71][8][23] + xor_out[72][8][23] + xor_out[73][8][23] + xor_out[74][8][23];
assign sum_out[15][8][23] = xor_out[75][8][23] + xor_out[76][8][23] + xor_out[77][8][23] + xor_out[78][8][23] + xor_out[79][8][23];
assign sum_out[16][8][23] = xor_out[80][8][23] + xor_out[81][8][23] + xor_out[82][8][23] + xor_out[83][8][23] + xor_out[84][8][23];
assign sum_out[17][8][23] = xor_out[85][8][23] + xor_out[86][8][23] + xor_out[87][8][23] + xor_out[88][8][23] + xor_out[89][8][23];
assign sum_out[18][8][23] = xor_out[90][8][23] + xor_out[91][8][23] + xor_out[92][8][23] + xor_out[93][8][23] + xor_out[94][8][23];
assign sum_out[19][8][23] = xor_out[95][8][23] + xor_out[96][8][23] + xor_out[97][8][23] + xor_out[98][8][23] + xor_out[99][8][23];

assign sum_out[0][9][0] = xor_out[0][9][0] + xor_out[1][9][0] + xor_out[2][9][0] + xor_out[3][9][0] + xor_out[4][9][0];
assign sum_out[1][9][0] = xor_out[5][9][0] + xor_out[6][9][0] + xor_out[7][9][0] + xor_out[8][9][0] + xor_out[9][9][0];
assign sum_out[2][9][0] = xor_out[10][9][0] + xor_out[11][9][0] + xor_out[12][9][0] + xor_out[13][9][0] + xor_out[14][9][0];
assign sum_out[3][9][0] = xor_out[15][9][0] + xor_out[16][9][0] + xor_out[17][9][0] + xor_out[18][9][0] + xor_out[19][9][0];
assign sum_out[4][9][0] = xor_out[20][9][0] + xor_out[21][9][0] + xor_out[22][9][0] + xor_out[23][9][0] + xor_out[24][9][0];
assign sum_out[5][9][0] = xor_out[25][9][0] + xor_out[26][9][0] + xor_out[27][9][0] + xor_out[28][9][0] + xor_out[29][9][0];
assign sum_out[6][9][0] = xor_out[30][9][0] + xor_out[31][9][0] + xor_out[32][9][0] + xor_out[33][9][0] + xor_out[34][9][0];
assign sum_out[7][9][0] = xor_out[35][9][0] + xor_out[36][9][0] + xor_out[37][9][0] + xor_out[38][9][0] + xor_out[39][9][0];
assign sum_out[8][9][0] = xor_out[40][9][0] + xor_out[41][9][0] + xor_out[42][9][0] + xor_out[43][9][0] + xor_out[44][9][0];
assign sum_out[9][9][0] = xor_out[45][9][0] + xor_out[46][9][0] + xor_out[47][9][0] + xor_out[48][9][0] + xor_out[49][9][0];
assign sum_out[10][9][0] = xor_out[50][9][0] + xor_out[51][9][0] + xor_out[52][9][0] + xor_out[53][9][0] + xor_out[54][9][0];
assign sum_out[11][9][0] = xor_out[55][9][0] + xor_out[56][9][0] + xor_out[57][9][0] + xor_out[58][9][0] + xor_out[59][9][0];
assign sum_out[12][9][0] = xor_out[60][9][0] + xor_out[61][9][0] + xor_out[62][9][0] + xor_out[63][9][0] + xor_out[64][9][0];
assign sum_out[13][9][0] = xor_out[65][9][0] + xor_out[66][9][0] + xor_out[67][9][0] + xor_out[68][9][0] + xor_out[69][9][0];
assign sum_out[14][9][0] = xor_out[70][9][0] + xor_out[71][9][0] + xor_out[72][9][0] + xor_out[73][9][0] + xor_out[74][9][0];
assign sum_out[15][9][0] = xor_out[75][9][0] + xor_out[76][9][0] + xor_out[77][9][0] + xor_out[78][9][0] + xor_out[79][9][0];
assign sum_out[16][9][0] = xor_out[80][9][0] + xor_out[81][9][0] + xor_out[82][9][0] + xor_out[83][9][0] + xor_out[84][9][0];
assign sum_out[17][9][0] = xor_out[85][9][0] + xor_out[86][9][0] + xor_out[87][9][0] + xor_out[88][9][0] + xor_out[89][9][0];
assign sum_out[18][9][0] = xor_out[90][9][0] + xor_out[91][9][0] + xor_out[92][9][0] + xor_out[93][9][0] + xor_out[94][9][0];
assign sum_out[19][9][0] = xor_out[95][9][0] + xor_out[96][9][0] + xor_out[97][9][0] + xor_out[98][9][0] + xor_out[99][9][0];

assign sum_out[0][9][1] = xor_out[0][9][1] + xor_out[1][9][1] + xor_out[2][9][1] + xor_out[3][9][1] + xor_out[4][9][1];
assign sum_out[1][9][1] = xor_out[5][9][1] + xor_out[6][9][1] + xor_out[7][9][1] + xor_out[8][9][1] + xor_out[9][9][1];
assign sum_out[2][9][1] = xor_out[10][9][1] + xor_out[11][9][1] + xor_out[12][9][1] + xor_out[13][9][1] + xor_out[14][9][1];
assign sum_out[3][9][1] = xor_out[15][9][1] + xor_out[16][9][1] + xor_out[17][9][1] + xor_out[18][9][1] + xor_out[19][9][1];
assign sum_out[4][9][1] = xor_out[20][9][1] + xor_out[21][9][1] + xor_out[22][9][1] + xor_out[23][9][1] + xor_out[24][9][1];
assign sum_out[5][9][1] = xor_out[25][9][1] + xor_out[26][9][1] + xor_out[27][9][1] + xor_out[28][9][1] + xor_out[29][9][1];
assign sum_out[6][9][1] = xor_out[30][9][1] + xor_out[31][9][1] + xor_out[32][9][1] + xor_out[33][9][1] + xor_out[34][9][1];
assign sum_out[7][9][1] = xor_out[35][9][1] + xor_out[36][9][1] + xor_out[37][9][1] + xor_out[38][9][1] + xor_out[39][9][1];
assign sum_out[8][9][1] = xor_out[40][9][1] + xor_out[41][9][1] + xor_out[42][9][1] + xor_out[43][9][1] + xor_out[44][9][1];
assign sum_out[9][9][1] = xor_out[45][9][1] + xor_out[46][9][1] + xor_out[47][9][1] + xor_out[48][9][1] + xor_out[49][9][1];
assign sum_out[10][9][1] = xor_out[50][9][1] + xor_out[51][9][1] + xor_out[52][9][1] + xor_out[53][9][1] + xor_out[54][9][1];
assign sum_out[11][9][1] = xor_out[55][9][1] + xor_out[56][9][1] + xor_out[57][9][1] + xor_out[58][9][1] + xor_out[59][9][1];
assign sum_out[12][9][1] = xor_out[60][9][1] + xor_out[61][9][1] + xor_out[62][9][1] + xor_out[63][9][1] + xor_out[64][9][1];
assign sum_out[13][9][1] = xor_out[65][9][1] + xor_out[66][9][1] + xor_out[67][9][1] + xor_out[68][9][1] + xor_out[69][9][1];
assign sum_out[14][9][1] = xor_out[70][9][1] + xor_out[71][9][1] + xor_out[72][9][1] + xor_out[73][9][1] + xor_out[74][9][1];
assign sum_out[15][9][1] = xor_out[75][9][1] + xor_out[76][9][1] + xor_out[77][9][1] + xor_out[78][9][1] + xor_out[79][9][1];
assign sum_out[16][9][1] = xor_out[80][9][1] + xor_out[81][9][1] + xor_out[82][9][1] + xor_out[83][9][1] + xor_out[84][9][1];
assign sum_out[17][9][1] = xor_out[85][9][1] + xor_out[86][9][1] + xor_out[87][9][1] + xor_out[88][9][1] + xor_out[89][9][1];
assign sum_out[18][9][1] = xor_out[90][9][1] + xor_out[91][9][1] + xor_out[92][9][1] + xor_out[93][9][1] + xor_out[94][9][1];
assign sum_out[19][9][1] = xor_out[95][9][1] + xor_out[96][9][1] + xor_out[97][9][1] + xor_out[98][9][1] + xor_out[99][9][1];

assign sum_out[0][9][2] = xor_out[0][9][2] + xor_out[1][9][2] + xor_out[2][9][2] + xor_out[3][9][2] + xor_out[4][9][2];
assign sum_out[1][9][2] = xor_out[5][9][2] + xor_out[6][9][2] + xor_out[7][9][2] + xor_out[8][9][2] + xor_out[9][9][2];
assign sum_out[2][9][2] = xor_out[10][9][2] + xor_out[11][9][2] + xor_out[12][9][2] + xor_out[13][9][2] + xor_out[14][9][2];
assign sum_out[3][9][2] = xor_out[15][9][2] + xor_out[16][9][2] + xor_out[17][9][2] + xor_out[18][9][2] + xor_out[19][9][2];
assign sum_out[4][9][2] = xor_out[20][9][2] + xor_out[21][9][2] + xor_out[22][9][2] + xor_out[23][9][2] + xor_out[24][9][2];
assign sum_out[5][9][2] = xor_out[25][9][2] + xor_out[26][9][2] + xor_out[27][9][2] + xor_out[28][9][2] + xor_out[29][9][2];
assign sum_out[6][9][2] = xor_out[30][9][2] + xor_out[31][9][2] + xor_out[32][9][2] + xor_out[33][9][2] + xor_out[34][9][2];
assign sum_out[7][9][2] = xor_out[35][9][2] + xor_out[36][9][2] + xor_out[37][9][2] + xor_out[38][9][2] + xor_out[39][9][2];
assign sum_out[8][9][2] = xor_out[40][9][2] + xor_out[41][9][2] + xor_out[42][9][2] + xor_out[43][9][2] + xor_out[44][9][2];
assign sum_out[9][9][2] = xor_out[45][9][2] + xor_out[46][9][2] + xor_out[47][9][2] + xor_out[48][9][2] + xor_out[49][9][2];
assign sum_out[10][9][2] = xor_out[50][9][2] + xor_out[51][9][2] + xor_out[52][9][2] + xor_out[53][9][2] + xor_out[54][9][2];
assign sum_out[11][9][2] = xor_out[55][9][2] + xor_out[56][9][2] + xor_out[57][9][2] + xor_out[58][9][2] + xor_out[59][9][2];
assign sum_out[12][9][2] = xor_out[60][9][2] + xor_out[61][9][2] + xor_out[62][9][2] + xor_out[63][9][2] + xor_out[64][9][2];
assign sum_out[13][9][2] = xor_out[65][9][2] + xor_out[66][9][2] + xor_out[67][9][2] + xor_out[68][9][2] + xor_out[69][9][2];
assign sum_out[14][9][2] = xor_out[70][9][2] + xor_out[71][9][2] + xor_out[72][9][2] + xor_out[73][9][2] + xor_out[74][9][2];
assign sum_out[15][9][2] = xor_out[75][9][2] + xor_out[76][9][2] + xor_out[77][9][2] + xor_out[78][9][2] + xor_out[79][9][2];
assign sum_out[16][9][2] = xor_out[80][9][2] + xor_out[81][9][2] + xor_out[82][9][2] + xor_out[83][9][2] + xor_out[84][9][2];
assign sum_out[17][9][2] = xor_out[85][9][2] + xor_out[86][9][2] + xor_out[87][9][2] + xor_out[88][9][2] + xor_out[89][9][2];
assign sum_out[18][9][2] = xor_out[90][9][2] + xor_out[91][9][2] + xor_out[92][9][2] + xor_out[93][9][2] + xor_out[94][9][2];
assign sum_out[19][9][2] = xor_out[95][9][2] + xor_out[96][9][2] + xor_out[97][9][2] + xor_out[98][9][2] + xor_out[99][9][2];

assign sum_out[0][9][3] = xor_out[0][9][3] + xor_out[1][9][3] + xor_out[2][9][3] + xor_out[3][9][3] + xor_out[4][9][3];
assign sum_out[1][9][3] = xor_out[5][9][3] + xor_out[6][9][3] + xor_out[7][9][3] + xor_out[8][9][3] + xor_out[9][9][3];
assign sum_out[2][9][3] = xor_out[10][9][3] + xor_out[11][9][3] + xor_out[12][9][3] + xor_out[13][9][3] + xor_out[14][9][3];
assign sum_out[3][9][3] = xor_out[15][9][3] + xor_out[16][9][3] + xor_out[17][9][3] + xor_out[18][9][3] + xor_out[19][9][3];
assign sum_out[4][9][3] = xor_out[20][9][3] + xor_out[21][9][3] + xor_out[22][9][3] + xor_out[23][9][3] + xor_out[24][9][3];
assign sum_out[5][9][3] = xor_out[25][9][3] + xor_out[26][9][3] + xor_out[27][9][3] + xor_out[28][9][3] + xor_out[29][9][3];
assign sum_out[6][9][3] = xor_out[30][9][3] + xor_out[31][9][3] + xor_out[32][9][3] + xor_out[33][9][3] + xor_out[34][9][3];
assign sum_out[7][9][3] = xor_out[35][9][3] + xor_out[36][9][3] + xor_out[37][9][3] + xor_out[38][9][3] + xor_out[39][9][3];
assign sum_out[8][9][3] = xor_out[40][9][3] + xor_out[41][9][3] + xor_out[42][9][3] + xor_out[43][9][3] + xor_out[44][9][3];
assign sum_out[9][9][3] = xor_out[45][9][3] + xor_out[46][9][3] + xor_out[47][9][3] + xor_out[48][9][3] + xor_out[49][9][3];
assign sum_out[10][9][3] = xor_out[50][9][3] + xor_out[51][9][3] + xor_out[52][9][3] + xor_out[53][9][3] + xor_out[54][9][3];
assign sum_out[11][9][3] = xor_out[55][9][3] + xor_out[56][9][3] + xor_out[57][9][3] + xor_out[58][9][3] + xor_out[59][9][3];
assign sum_out[12][9][3] = xor_out[60][9][3] + xor_out[61][9][3] + xor_out[62][9][3] + xor_out[63][9][3] + xor_out[64][9][3];
assign sum_out[13][9][3] = xor_out[65][9][3] + xor_out[66][9][3] + xor_out[67][9][3] + xor_out[68][9][3] + xor_out[69][9][3];
assign sum_out[14][9][3] = xor_out[70][9][3] + xor_out[71][9][3] + xor_out[72][9][3] + xor_out[73][9][3] + xor_out[74][9][3];
assign sum_out[15][9][3] = xor_out[75][9][3] + xor_out[76][9][3] + xor_out[77][9][3] + xor_out[78][9][3] + xor_out[79][9][3];
assign sum_out[16][9][3] = xor_out[80][9][3] + xor_out[81][9][3] + xor_out[82][9][3] + xor_out[83][9][3] + xor_out[84][9][3];
assign sum_out[17][9][3] = xor_out[85][9][3] + xor_out[86][9][3] + xor_out[87][9][3] + xor_out[88][9][3] + xor_out[89][9][3];
assign sum_out[18][9][3] = xor_out[90][9][3] + xor_out[91][9][3] + xor_out[92][9][3] + xor_out[93][9][3] + xor_out[94][9][3];
assign sum_out[19][9][3] = xor_out[95][9][3] + xor_out[96][9][3] + xor_out[97][9][3] + xor_out[98][9][3] + xor_out[99][9][3];

assign sum_out[0][9][4] = xor_out[0][9][4] + xor_out[1][9][4] + xor_out[2][9][4] + xor_out[3][9][4] + xor_out[4][9][4];
assign sum_out[1][9][4] = xor_out[5][9][4] + xor_out[6][9][4] + xor_out[7][9][4] + xor_out[8][9][4] + xor_out[9][9][4];
assign sum_out[2][9][4] = xor_out[10][9][4] + xor_out[11][9][4] + xor_out[12][9][4] + xor_out[13][9][4] + xor_out[14][9][4];
assign sum_out[3][9][4] = xor_out[15][9][4] + xor_out[16][9][4] + xor_out[17][9][4] + xor_out[18][9][4] + xor_out[19][9][4];
assign sum_out[4][9][4] = xor_out[20][9][4] + xor_out[21][9][4] + xor_out[22][9][4] + xor_out[23][9][4] + xor_out[24][9][4];
assign sum_out[5][9][4] = xor_out[25][9][4] + xor_out[26][9][4] + xor_out[27][9][4] + xor_out[28][9][4] + xor_out[29][9][4];
assign sum_out[6][9][4] = xor_out[30][9][4] + xor_out[31][9][4] + xor_out[32][9][4] + xor_out[33][9][4] + xor_out[34][9][4];
assign sum_out[7][9][4] = xor_out[35][9][4] + xor_out[36][9][4] + xor_out[37][9][4] + xor_out[38][9][4] + xor_out[39][9][4];
assign sum_out[8][9][4] = xor_out[40][9][4] + xor_out[41][9][4] + xor_out[42][9][4] + xor_out[43][9][4] + xor_out[44][9][4];
assign sum_out[9][9][4] = xor_out[45][9][4] + xor_out[46][9][4] + xor_out[47][9][4] + xor_out[48][9][4] + xor_out[49][9][4];
assign sum_out[10][9][4] = xor_out[50][9][4] + xor_out[51][9][4] + xor_out[52][9][4] + xor_out[53][9][4] + xor_out[54][9][4];
assign sum_out[11][9][4] = xor_out[55][9][4] + xor_out[56][9][4] + xor_out[57][9][4] + xor_out[58][9][4] + xor_out[59][9][4];
assign sum_out[12][9][4] = xor_out[60][9][4] + xor_out[61][9][4] + xor_out[62][9][4] + xor_out[63][9][4] + xor_out[64][9][4];
assign sum_out[13][9][4] = xor_out[65][9][4] + xor_out[66][9][4] + xor_out[67][9][4] + xor_out[68][9][4] + xor_out[69][9][4];
assign sum_out[14][9][4] = xor_out[70][9][4] + xor_out[71][9][4] + xor_out[72][9][4] + xor_out[73][9][4] + xor_out[74][9][4];
assign sum_out[15][9][4] = xor_out[75][9][4] + xor_out[76][9][4] + xor_out[77][9][4] + xor_out[78][9][4] + xor_out[79][9][4];
assign sum_out[16][9][4] = xor_out[80][9][4] + xor_out[81][9][4] + xor_out[82][9][4] + xor_out[83][9][4] + xor_out[84][9][4];
assign sum_out[17][9][4] = xor_out[85][9][4] + xor_out[86][9][4] + xor_out[87][9][4] + xor_out[88][9][4] + xor_out[89][9][4];
assign sum_out[18][9][4] = xor_out[90][9][4] + xor_out[91][9][4] + xor_out[92][9][4] + xor_out[93][9][4] + xor_out[94][9][4];
assign sum_out[19][9][4] = xor_out[95][9][4] + xor_out[96][9][4] + xor_out[97][9][4] + xor_out[98][9][4] + xor_out[99][9][4];

assign sum_out[0][9][5] = xor_out[0][9][5] + xor_out[1][9][5] + xor_out[2][9][5] + xor_out[3][9][5] + xor_out[4][9][5];
assign sum_out[1][9][5] = xor_out[5][9][5] + xor_out[6][9][5] + xor_out[7][9][5] + xor_out[8][9][5] + xor_out[9][9][5];
assign sum_out[2][9][5] = xor_out[10][9][5] + xor_out[11][9][5] + xor_out[12][9][5] + xor_out[13][9][5] + xor_out[14][9][5];
assign sum_out[3][9][5] = xor_out[15][9][5] + xor_out[16][9][5] + xor_out[17][9][5] + xor_out[18][9][5] + xor_out[19][9][5];
assign sum_out[4][9][5] = xor_out[20][9][5] + xor_out[21][9][5] + xor_out[22][9][5] + xor_out[23][9][5] + xor_out[24][9][5];
assign sum_out[5][9][5] = xor_out[25][9][5] + xor_out[26][9][5] + xor_out[27][9][5] + xor_out[28][9][5] + xor_out[29][9][5];
assign sum_out[6][9][5] = xor_out[30][9][5] + xor_out[31][9][5] + xor_out[32][9][5] + xor_out[33][9][5] + xor_out[34][9][5];
assign sum_out[7][9][5] = xor_out[35][9][5] + xor_out[36][9][5] + xor_out[37][9][5] + xor_out[38][9][5] + xor_out[39][9][5];
assign sum_out[8][9][5] = xor_out[40][9][5] + xor_out[41][9][5] + xor_out[42][9][5] + xor_out[43][9][5] + xor_out[44][9][5];
assign sum_out[9][9][5] = xor_out[45][9][5] + xor_out[46][9][5] + xor_out[47][9][5] + xor_out[48][9][5] + xor_out[49][9][5];
assign sum_out[10][9][5] = xor_out[50][9][5] + xor_out[51][9][5] + xor_out[52][9][5] + xor_out[53][9][5] + xor_out[54][9][5];
assign sum_out[11][9][5] = xor_out[55][9][5] + xor_out[56][9][5] + xor_out[57][9][5] + xor_out[58][9][5] + xor_out[59][9][5];
assign sum_out[12][9][5] = xor_out[60][9][5] + xor_out[61][9][5] + xor_out[62][9][5] + xor_out[63][9][5] + xor_out[64][9][5];
assign sum_out[13][9][5] = xor_out[65][9][5] + xor_out[66][9][5] + xor_out[67][9][5] + xor_out[68][9][5] + xor_out[69][9][5];
assign sum_out[14][9][5] = xor_out[70][9][5] + xor_out[71][9][5] + xor_out[72][9][5] + xor_out[73][9][5] + xor_out[74][9][5];
assign sum_out[15][9][5] = xor_out[75][9][5] + xor_out[76][9][5] + xor_out[77][9][5] + xor_out[78][9][5] + xor_out[79][9][5];
assign sum_out[16][9][5] = xor_out[80][9][5] + xor_out[81][9][5] + xor_out[82][9][5] + xor_out[83][9][5] + xor_out[84][9][5];
assign sum_out[17][9][5] = xor_out[85][9][5] + xor_out[86][9][5] + xor_out[87][9][5] + xor_out[88][9][5] + xor_out[89][9][5];
assign sum_out[18][9][5] = xor_out[90][9][5] + xor_out[91][9][5] + xor_out[92][9][5] + xor_out[93][9][5] + xor_out[94][9][5];
assign sum_out[19][9][5] = xor_out[95][9][5] + xor_out[96][9][5] + xor_out[97][9][5] + xor_out[98][9][5] + xor_out[99][9][5];

assign sum_out[0][9][6] = xor_out[0][9][6] + xor_out[1][9][6] + xor_out[2][9][6] + xor_out[3][9][6] + xor_out[4][9][6];
assign sum_out[1][9][6] = xor_out[5][9][6] + xor_out[6][9][6] + xor_out[7][9][6] + xor_out[8][9][6] + xor_out[9][9][6];
assign sum_out[2][9][6] = xor_out[10][9][6] + xor_out[11][9][6] + xor_out[12][9][6] + xor_out[13][9][6] + xor_out[14][9][6];
assign sum_out[3][9][6] = xor_out[15][9][6] + xor_out[16][9][6] + xor_out[17][9][6] + xor_out[18][9][6] + xor_out[19][9][6];
assign sum_out[4][9][6] = xor_out[20][9][6] + xor_out[21][9][6] + xor_out[22][9][6] + xor_out[23][9][6] + xor_out[24][9][6];
assign sum_out[5][9][6] = xor_out[25][9][6] + xor_out[26][9][6] + xor_out[27][9][6] + xor_out[28][9][6] + xor_out[29][9][6];
assign sum_out[6][9][6] = xor_out[30][9][6] + xor_out[31][9][6] + xor_out[32][9][6] + xor_out[33][9][6] + xor_out[34][9][6];
assign sum_out[7][9][6] = xor_out[35][9][6] + xor_out[36][9][6] + xor_out[37][9][6] + xor_out[38][9][6] + xor_out[39][9][6];
assign sum_out[8][9][6] = xor_out[40][9][6] + xor_out[41][9][6] + xor_out[42][9][6] + xor_out[43][9][6] + xor_out[44][9][6];
assign sum_out[9][9][6] = xor_out[45][9][6] + xor_out[46][9][6] + xor_out[47][9][6] + xor_out[48][9][6] + xor_out[49][9][6];
assign sum_out[10][9][6] = xor_out[50][9][6] + xor_out[51][9][6] + xor_out[52][9][6] + xor_out[53][9][6] + xor_out[54][9][6];
assign sum_out[11][9][6] = xor_out[55][9][6] + xor_out[56][9][6] + xor_out[57][9][6] + xor_out[58][9][6] + xor_out[59][9][6];
assign sum_out[12][9][6] = xor_out[60][9][6] + xor_out[61][9][6] + xor_out[62][9][6] + xor_out[63][9][6] + xor_out[64][9][6];
assign sum_out[13][9][6] = xor_out[65][9][6] + xor_out[66][9][6] + xor_out[67][9][6] + xor_out[68][9][6] + xor_out[69][9][6];
assign sum_out[14][9][6] = xor_out[70][9][6] + xor_out[71][9][6] + xor_out[72][9][6] + xor_out[73][9][6] + xor_out[74][9][6];
assign sum_out[15][9][6] = xor_out[75][9][6] + xor_out[76][9][6] + xor_out[77][9][6] + xor_out[78][9][6] + xor_out[79][9][6];
assign sum_out[16][9][6] = xor_out[80][9][6] + xor_out[81][9][6] + xor_out[82][9][6] + xor_out[83][9][6] + xor_out[84][9][6];
assign sum_out[17][9][6] = xor_out[85][9][6] + xor_out[86][9][6] + xor_out[87][9][6] + xor_out[88][9][6] + xor_out[89][9][6];
assign sum_out[18][9][6] = xor_out[90][9][6] + xor_out[91][9][6] + xor_out[92][9][6] + xor_out[93][9][6] + xor_out[94][9][6];
assign sum_out[19][9][6] = xor_out[95][9][6] + xor_out[96][9][6] + xor_out[97][9][6] + xor_out[98][9][6] + xor_out[99][9][6];

assign sum_out[0][9][7] = xor_out[0][9][7] + xor_out[1][9][7] + xor_out[2][9][7] + xor_out[3][9][7] + xor_out[4][9][7];
assign sum_out[1][9][7] = xor_out[5][9][7] + xor_out[6][9][7] + xor_out[7][9][7] + xor_out[8][9][7] + xor_out[9][9][7];
assign sum_out[2][9][7] = xor_out[10][9][7] + xor_out[11][9][7] + xor_out[12][9][7] + xor_out[13][9][7] + xor_out[14][9][7];
assign sum_out[3][9][7] = xor_out[15][9][7] + xor_out[16][9][7] + xor_out[17][9][7] + xor_out[18][9][7] + xor_out[19][9][7];
assign sum_out[4][9][7] = xor_out[20][9][7] + xor_out[21][9][7] + xor_out[22][9][7] + xor_out[23][9][7] + xor_out[24][9][7];
assign sum_out[5][9][7] = xor_out[25][9][7] + xor_out[26][9][7] + xor_out[27][9][7] + xor_out[28][9][7] + xor_out[29][9][7];
assign sum_out[6][9][7] = xor_out[30][9][7] + xor_out[31][9][7] + xor_out[32][9][7] + xor_out[33][9][7] + xor_out[34][9][7];
assign sum_out[7][9][7] = xor_out[35][9][7] + xor_out[36][9][7] + xor_out[37][9][7] + xor_out[38][9][7] + xor_out[39][9][7];
assign sum_out[8][9][7] = xor_out[40][9][7] + xor_out[41][9][7] + xor_out[42][9][7] + xor_out[43][9][7] + xor_out[44][9][7];
assign sum_out[9][9][7] = xor_out[45][9][7] + xor_out[46][9][7] + xor_out[47][9][7] + xor_out[48][9][7] + xor_out[49][9][7];
assign sum_out[10][9][7] = xor_out[50][9][7] + xor_out[51][9][7] + xor_out[52][9][7] + xor_out[53][9][7] + xor_out[54][9][7];
assign sum_out[11][9][7] = xor_out[55][9][7] + xor_out[56][9][7] + xor_out[57][9][7] + xor_out[58][9][7] + xor_out[59][9][7];
assign sum_out[12][9][7] = xor_out[60][9][7] + xor_out[61][9][7] + xor_out[62][9][7] + xor_out[63][9][7] + xor_out[64][9][7];
assign sum_out[13][9][7] = xor_out[65][9][7] + xor_out[66][9][7] + xor_out[67][9][7] + xor_out[68][9][7] + xor_out[69][9][7];
assign sum_out[14][9][7] = xor_out[70][9][7] + xor_out[71][9][7] + xor_out[72][9][7] + xor_out[73][9][7] + xor_out[74][9][7];
assign sum_out[15][9][7] = xor_out[75][9][7] + xor_out[76][9][7] + xor_out[77][9][7] + xor_out[78][9][7] + xor_out[79][9][7];
assign sum_out[16][9][7] = xor_out[80][9][7] + xor_out[81][9][7] + xor_out[82][9][7] + xor_out[83][9][7] + xor_out[84][9][7];
assign sum_out[17][9][7] = xor_out[85][9][7] + xor_out[86][9][7] + xor_out[87][9][7] + xor_out[88][9][7] + xor_out[89][9][7];
assign sum_out[18][9][7] = xor_out[90][9][7] + xor_out[91][9][7] + xor_out[92][9][7] + xor_out[93][9][7] + xor_out[94][9][7];
assign sum_out[19][9][7] = xor_out[95][9][7] + xor_out[96][9][7] + xor_out[97][9][7] + xor_out[98][9][7] + xor_out[99][9][7];

assign sum_out[0][9][8] = xor_out[0][9][8] + xor_out[1][9][8] + xor_out[2][9][8] + xor_out[3][9][8] + xor_out[4][9][8];
assign sum_out[1][9][8] = xor_out[5][9][8] + xor_out[6][9][8] + xor_out[7][9][8] + xor_out[8][9][8] + xor_out[9][9][8];
assign sum_out[2][9][8] = xor_out[10][9][8] + xor_out[11][9][8] + xor_out[12][9][8] + xor_out[13][9][8] + xor_out[14][9][8];
assign sum_out[3][9][8] = xor_out[15][9][8] + xor_out[16][9][8] + xor_out[17][9][8] + xor_out[18][9][8] + xor_out[19][9][8];
assign sum_out[4][9][8] = xor_out[20][9][8] + xor_out[21][9][8] + xor_out[22][9][8] + xor_out[23][9][8] + xor_out[24][9][8];
assign sum_out[5][9][8] = xor_out[25][9][8] + xor_out[26][9][8] + xor_out[27][9][8] + xor_out[28][9][8] + xor_out[29][9][8];
assign sum_out[6][9][8] = xor_out[30][9][8] + xor_out[31][9][8] + xor_out[32][9][8] + xor_out[33][9][8] + xor_out[34][9][8];
assign sum_out[7][9][8] = xor_out[35][9][8] + xor_out[36][9][8] + xor_out[37][9][8] + xor_out[38][9][8] + xor_out[39][9][8];
assign sum_out[8][9][8] = xor_out[40][9][8] + xor_out[41][9][8] + xor_out[42][9][8] + xor_out[43][9][8] + xor_out[44][9][8];
assign sum_out[9][9][8] = xor_out[45][9][8] + xor_out[46][9][8] + xor_out[47][9][8] + xor_out[48][9][8] + xor_out[49][9][8];
assign sum_out[10][9][8] = xor_out[50][9][8] + xor_out[51][9][8] + xor_out[52][9][8] + xor_out[53][9][8] + xor_out[54][9][8];
assign sum_out[11][9][8] = xor_out[55][9][8] + xor_out[56][9][8] + xor_out[57][9][8] + xor_out[58][9][8] + xor_out[59][9][8];
assign sum_out[12][9][8] = xor_out[60][9][8] + xor_out[61][9][8] + xor_out[62][9][8] + xor_out[63][9][8] + xor_out[64][9][8];
assign sum_out[13][9][8] = xor_out[65][9][8] + xor_out[66][9][8] + xor_out[67][9][8] + xor_out[68][9][8] + xor_out[69][9][8];
assign sum_out[14][9][8] = xor_out[70][9][8] + xor_out[71][9][8] + xor_out[72][9][8] + xor_out[73][9][8] + xor_out[74][9][8];
assign sum_out[15][9][8] = xor_out[75][9][8] + xor_out[76][9][8] + xor_out[77][9][8] + xor_out[78][9][8] + xor_out[79][9][8];
assign sum_out[16][9][8] = xor_out[80][9][8] + xor_out[81][9][8] + xor_out[82][9][8] + xor_out[83][9][8] + xor_out[84][9][8];
assign sum_out[17][9][8] = xor_out[85][9][8] + xor_out[86][9][8] + xor_out[87][9][8] + xor_out[88][9][8] + xor_out[89][9][8];
assign sum_out[18][9][8] = xor_out[90][9][8] + xor_out[91][9][8] + xor_out[92][9][8] + xor_out[93][9][8] + xor_out[94][9][8];
assign sum_out[19][9][8] = xor_out[95][9][8] + xor_out[96][9][8] + xor_out[97][9][8] + xor_out[98][9][8] + xor_out[99][9][8];

assign sum_out[0][9][9] = xor_out[0][9][9] + xor_out[1][9][9] + xor_out[2][9][9] + xor_out[3][9][9] + xor_out[4][9][9];
assign sum_out[1][9][9] = xor_out[5][9][9] + xor_out[6][9][9] + xor_out[7][9][9] + xor_out[8][9][9] + xor_out[9][9][9];
assign sum_out[2][9][9] = xor_out[10][9][9] + xor_out[11][9][9] + xor_out[12][9][9] + xor_out[13][9][9] + xor_out[14][9][9];
assign sum_out[3][9][9] = xor_out[15][9][9] + xor_out[16][9][9] + xor_out[17][9][9] + xor_out[18][9][9] + xor_out[19][9][9];
assign sum_out[4][9][9] = xor_out[20][9][9] + xor_out[21][9][9] + xor_out[22][9][9] + xor_out[23][9][9] + xor_out[24][9][9];
assign sum_out[5][9][9] = xor_out[25][9][9] + xor_out[26][9][9] + xor_out[27][9][9] + xor_out[28][9][9] + xor_out[29][9][9];
assign sum_out[6][9][9] = xor_out[30][9][9] + xor_out[31][9][9] + xor_out[32][9][9] + xor_out[33][9][9] + xor_out[34][9][9];
assign sum_out[7][9][9] = xor_out[35][9][9] + xor_out[36][9][9] + xor_out[37][9][9] + xor_out[38][9][9] + xor_out[39][9][9];
assign sum_out[8][9][9] = xor_out[40][9][9] + xor_out[41][9][9] + xor_out[42][9][9] + xor_out[43][9][9] + xor_out[44][9][9];
assign sum_out[9][9][9] = xor_out[45][9][9] + xor_out[46][9][9] + xor_out[47][9][9] + xor_out[48][9][9] + xor_out[49][9][9];
assign sum_out[10][9][9] = xor_out[50][9][9] + xor_out[51][9][9] + xor_out[52][9][9] + xor_out[53][9][9] + xor_out[54][9][9];
assign sum_out[11][9][9] = xor_out[55][9][9] + xor_out[56][9][9] + xor_out[57][9][9] + xor_out[58][9][9] + xor_out[59][9][9];
assign sum_out[12][9][9] = xor_out[60][9][9] + xor_out[61][9][9] + xor_out[62][9][9] + xor_out[63][9][9] + xor_out[64][9][9];
assign sum_out[13][9][9] = xor_out[65][9][9] + xor_out[66][9][9] + xor_out[67][9][9] + xor_out[68][9][9] + xor_out[69][9][9];
assign sum_out[14][9][9] = xor_out[70][9][9] + xor_out[71][9][9] + xor_out[72][9][9] + xor_out[73][9][9] + xor_out[74][9][9];
assign sum_out[15][9][9] = xor_out[75][9][9] + xor_out[76][9][9] + xor_out[77][9][9] + xor_out[78][9][9] + xor_out[79][9][9];
assign sum_out[16][9][9] = xor_out[80][9][9] + xor_out[81][9][9] + xor_out[82][9][9] + xor_out[83][9][9] + xor_out[84][9][9];
assign sum_out[17][9][9] = xor_out[85][9][9] + xor_out[86][9][9] + xor_out[87][9][9] + xor_out[88][9][9] + xor_out[89][9][9];
assign sum_out[18][9][9] = xor_out[90][9][9] + xor_out[91][9][9] + xor_out[92][9][9] + xor_out[93][9][9] + xor_out[94][9][9];
assign sum_out[19][9][9] = xor_out[95][9][9] + xor_out[96][9][9] + xor_out[97][9][9] + xor_out[98][9][9] + xor_out[99][9][9];

assign sum_out[0][9][10] = xor_out[0][9][10] + xor_out[1][9][10] + xor_out[2][9][10] + xor_out[3][9][10] + xor_out[4][9][10];
assign sum_out[1][9][10] = xor_out[5][9][10] + xor_out[6][9][10] + xor_out[7][9][10] + xor_out[8][9][10] + xor_out[9][9][10];
assign sum_out[2][9][10] = xor_out[10][9][10] + xor_out[11][9][10] + xor_out[12][9][10] + xor_out[13][9][10] + xor_out[14][9][10];
assign sum_out[3][9][10] = xor_out[15][9][10] + xor_out[16][9][10] + xor_out[17][9][10] + xor_out[18][9][10] + xor_out[19][9][10];
assign sum_out[4][9][10] = xor_out[20][9][10] + xor_out[21][9][10] + xor_out[22][9][10] + xor_out[23][9][10] + xor_out[24][9][10];
assign sum_out[5][9][10] = xor_out[25][9][10] + xor_out[26][9][10] + xor_out[27][9][10] + xor_out[28][9][10] + xor_out[29][9][10];
assign sum_out[6][9][10] = xor_out[30][9][10] + xor_out[31][9][10] + xor_out[32][9][10] + xor_out[33][9][10] + xor_out[34][9][10];
assign sum_out[7][9][10] = xor_out[35][9][10] + xor_out[36][9][10] + xor_out[37][9][10] + xor_out[38][9][10] + xor_out[39][9][10];
assign sum_out[8][9][10] = xor_out[40][9][10] + xor_out[41][9][10] + xor_out[42][9][10] + xor_out[43][9][10] + xor_out[44][9][10];
assign sum_out[9][9][10] = xor_out[45][9][10] + xor_out[46][9][10] + xor_out[47][9][10] + xor_out[48][9][10] + xor_out[49][9][10];
assign sum_out[10][9][10] = xor_out[50][9][10] + xor_out[51][9][10] + xor_out[52][9][10] + xor_out[53][9][10] + xor_out[54][9][10];
assign sum_out[11][9][10] = xor_out[55][9][10] + xor_out[56][9][10] + xor_out[57][9][10] + xor_out[58][9][10] + xor_out[59][9][10];
assign sum_out[12][9][10] = xor_out[60][9][10] + xor_out[61][9][10] + xor_out[62][9][10] + xor_out[63][9][10] + xor_out[64][9][10];
assign sum_out[13][9][10] = xor_out[65][9][10] + xor_out[66][9][10] + xor_out[67][9][10] + xor_out[68][9][10] + xor_out[69][9][10];
assign sum_out[14][9][10] = xor_out[70][9][10] + xor_out[71][9][10] + xor_out[72][9][10] + xor_out[73][9][10] + xor_out[74][9][10];
assign sum_out[15][9][10] = xor_out[75][9][10] + xor_out[76][9][10] + xor_out[77][9][10] + xor_out[78][9][10] + xor_out[79][9][10];
assign sum_out[16][9][10] = xor_out[80][9][10] + xor_out[81][9][10] + xor_out[82][9][10] + xor_out[83][9][10] + xor_out[84][9][10];
assign sum_out[17][9][10] = xor_out[85][9][10] + xor_out[86][9][10] + xor_out[87][9][10] + xor_out[88][9][10] + xor_out[89][9][10];
assign sum_out[18][9][10] = xor_out[90][9][10] + xor_out[91][9][10] + xor_out[92][9][10] + xor_out[93][9][10] + xor_out[94][9][10];
assign sum_out[19][9][10] = xor_out[95][9][10] + xor_out[96][9][10] + xor_out[97][9][10] + xor_out[98][9][10] + xor_out[99][9][10];

assign sum_out[0][9][11] = xor_out[0][9][11] + xor_out[1][9][11] + xor_out[2][9][11] + xor_out[3][9][11] + xor_out[4][9][11];
assign sum_out[1][9][11] = xor_out[5][9][11] + xor_out[6][9][11] + xor_out[7][9][11] + xor_out[8][9][11] + xor_out[9][9][11];
assign sum_out[2][9][11] = xor_out[10][9][11] + xor_out[11][9][11] + xor_out[12][9][11] + xor_out[13][9][11] + xor_out[14][9][11];
assign sum_out[3][9][11] = xor_out[15][9][11] + xor_out[16][9][11] + xor_out[17][9][11] + xor_out[18][9][11] + xor_out[19][9][11];
assign sum_out[4][9][11] = xor_out[20][9][11] + xor_out[21][9][11] + xor_out[22][9][11] + xor_out[23][9][11] + xor_out[24][9][11];
assign sum_out[5][9][11] = xor_out[25][9][11] + xor_out[26][9][11] + xor_out[27][9][11] + xor_out[28][9][11] + xor_out[29][9][11];
assign sum_out[6][9][11] = xor_out[30][9][11] + xor_out[31][9][11] + xor_out[32][9][11] + xor_out[33][9][11] + xor_out[34][9][11];
assign sum_out[7][9][11] = xor_out[35][9][11] + xor_out[36][9][11] + xor_out[37][9][11] + xor_out[38][9][11] + xor_out[39][9][11];
assign sum_out[8][9][11] = xor_out[40][9][11] + xor_out[41][9][11] + xor_out[42][9][11] + xor_out[43][9][11] + xor_out[44][9][11];
assign sum_out[9][9][11] = xor_out[45][9][11] + xor_out[46][9][11] + xor_out[47][9][11] + xor_out[48][9][11] + xor_out[49][9][11];
assign sum_out[10][9][11] = xor_out[50][9][11] + xor_out[51][9][11] + xor_out[52][9][11] + xor_out[53][9][11] + xor_out[54][9][11];
assign sum_out[11][9][11] = xor_out[55][9][11] + xor_out[56][9][11] + xor_out[57][9][11] + xor_out[58][9][11] + xor_out[59][9][11];
assign sum_out[12][9][11] = xor_out[60][9][11] + xor_out[61][9][11] + xor_out[62][9][11] + xor_out[63][9][11] + xor_out[64][9][11];
assign sum_out[13][9][11] = xor_out[65][9][11] + xor_out[66][9][11] + xor_out[67][9][11] + xor_out[68][9][11] + xor_out[69][9][11];
assign sum_out[14][9][11] = xor_out[70][9][11] + xor_out[71][9][11] + xor_out[72][9][11] + xor_out[73][9][11] + xor_out[74][9][11];
assign sum_out[15][9][11] = xor_out[75][9][11] + xor_out[76][9][11] + xor_out[77][9][11] + xor_out[78][9][11] + xor_out[79][9][11];
assign sum_out[16][9][11] = xor_out[80][9][11] + xor_out[81][9][11] + xor_out[82][9][11] + xor_out[83][9][11] + xor_out[84][9][11];
assign sum_out[17][9][11] = xor_out[85][9][11] + xor_out[86][9][11] + xor_out[87][9][11] + xor_out[88][9][11] + xor_out[89][9][11];
assign sum_out[18][9][11] = xor_out[90][9][11] + xor_out[91][9][11] + xor_out[92][9][11] + xor_out[93][9][11] + xor_out[94][9][11];
assign sum_out[19][9][11] = xor_out[95][9][11] + xor_out[96][9][11] + xor_out[97][9][11] + xor_out[98][9][11] + xor_out[99][9][11];

assign sum_out[0][9][12] = xor_out[0][9][12] + xor_out[1][9][12] + xor_out[2][9][12] + xor_out[3][9][12] + xor_out[4][9][12];
assign sum_out[1][9][12] = xor_out[5][9][12] + xor_out[6][9][12] + xor_out[7][9][12] + xor_out[8][9][12] + xor_out[9][9][12];
assign sum_out[2][9][12] = xor_out[10][9][12] + xor_out[11][9][12] + xor_out[12][9][12] + xor_out[13][9][12] + xor_out[14][9][12];
assign sum_out[3][9][12] = xor_out[15][9][12] + xor_out[16][9][12] + xor_out[17][9][12] + xor_out[18][9][12] + xor_out[19][9][12];
assign sum_out[4][9][12] = xor_out[20][9][12] + xor_out[21][9][12] + xor_out[22][9][12] + xor_out[23][9][12] + xor_out[24][9][12];
assign sum_out[5][9][12] = xor_out[25][9][12] + xor_out[26][9][12] + xor_out[27][9][12] + xor_out[28][9][12] + xor_out[29][9][12];
assign sum_out[6][9][12] = xor_out[30][9][12] + xor_out[31][9][12] + xor_out[32][9][12] + xor_out[33][9][12] + xor_out[34][9][12];
assign sum_out[7][9][12] = xor_out[35][9][12] + xor_out[36][9][12] + xor_out[37][9][12] + xor_out[38][9][12] + xor_out[39][9][12];
assign sum_out[8][9][12] = xor_out[40][9][12] + xor_out[41][9][12] + xor_out[42][9][12] + xor_out[43][9][12] + xor_out[44][9][12];
assign sum_out[9][9][12] = xor_out[45][9][12] + xor_out[46][9][12] + xor_out[47][9][12] + xor_out[48][9][12] + xor_out[49][9][12];
assign sum_out[10][9][12] = xor_out[50][9][12] + xor_out[51][9][12] + xor_out[52][9][12] + xor_out[53][9][12] + xor_out[54][9][12];
assign sum_out[11][9][12] = xor_out[55][9][12] + xor_out[56][9][12] + xor_out[57][9][12] + xor_out[58][9][12] + xor_out[59][9][12];
assign sum_out[12][9][12] = xor_out[60][9][12] + xor_out[61][9][12] + xor_out[62][9][12] + xor_out[63][9][12] + xor_out[64][9][12];
assign sum_out[13][9][12] = xor_out[65][9][12] + xor_out[66][9][12] + xor_out[67][9][12] + xor_out[68][9][12] + xor_out[69][9][12];
assign sum_out[14][9][12] = xor_out[70][9][12] + xor_out[71][9][12] + xor_out[72][9][12] + xor_out[73][9][12] + xor_out[74][9][12];
assign sum_out[15][9][12] = xor_out[75][9][12] + xor_out[76][9][12] + xor_out[77][9][12] + xor_out[78][9][12] + xor_out[79][9][12];
assign sum_out[16][9][12] = xor_out[80][9][12] + xor_out[81][9][12] + xor_out[82][9][12] + xor_out[83][9][12] + xor_out[84][9][12];
assign sum_out[17][9][12] = xor_out[85][9][12] + xor_out[86][9][12] + xor_out[87][9][12] + xor_out[88][9][12] + xor_out[89][9][12];
assign sum_out[18][9][12] = xor_out[90][9][12] + xor_out[91][9][12] + xor_out[92][9][12] + xor_out[93][9][12] + xor_out[94][9][12];
assign sum_out[19][9][12] = xor_out[95][9][12] + xor_out[96][9][12] + xor_out[97][9][12] + xor_out[98][9][12] + xor_out[99][9][12];

assign sum_out[0][9][13] = xor_out[0][9][13] + xor_out[1][9][13] + xor_out[2][9][13] + xor_out[3][9][13] + xor_out[4][9][13];
assign sum_out[1][9][13] = xor_out[5][9][13] + xor_out[6][9][13] + xor_out[7][9][13] + xor_out[8][9][13] + xor_out[9][9][13];
assign sum_out[2][9][13] = xor_out[10][9][13] + xor_out[11][9][13] + xor_out[12][9][13] + xor_out[13][9][13] + xor_out[14][9][13];
assign sum_out[3][9][13] = xor_out[15][9][13] + xor_out[16][9][13] + xor_out[17][9][13] + xor_out[18][9][13] + xor_out[19][9][13];
assign sum_out[4][9][13] = xor_out[20][9][13] + xor_out[21][9][13] + xor_out[22][9][13] + xor_out[23][9][13] + xor_out[24][9][13];
assign sum_out[5][9][13] = xor_out[25][9][13] + xor_out[26][9][13] + xor_out[27][9][13] + xor_out[28][9][13] + xor_out[29][9][13];
assign sum_out[6][9][13] = xor_out[30][9][13] + xor_out[31][9][13] + xor_out[32][9][13] + xor_out[33][9][13] + xor_out[34][9][13];
assign sum_out[7][9][13] = xor_out[35][9][13] + xor_out[36][9][13] + xor_out[37][9][13] + xor_out[38][9][13] + xor_out[39][9][13];
assign sum_out[8][9][13] = xor_out[40][9][13] + xor_out[41][9][13] + xor_out[42][9][13] + xor_out[43][9][13] + xor_out[44][9][13];
assign sum_out[9][9][13] = xor_out[45][9][13] + xor_out[46][9][13] + xor_out[47][9][13] + xor_out[48][9][13] + xor_out[49][9][13];
assign sum_out[10][9][13] = xor_out[50][9][13] + xor_out[51][9][13] + xor_out[52][9][13] + xor_out[53][9][13] + xor_out[54][9][13];
assign sum_out[11][9][13] = xor_out[55][9][13] + xor_out[56][9][13] + xor_out[57][9][13] + xor_out[58][9][13] + xor_out[59][9][13];
assign sum_out[12][9][13] = xor_out[60][9][13] + xor_out[61][9][13] + xor_out[62][9][13] + xor_out[63][9][13] + xor_out[64][9][13];
assign sum_out[13][9][13] = xor_out[65][9][13] + xor_out[66][9][13] + xor_out[67][9][13] + xor_out[68][9][13] + xor_out[69][9][13];
assign sum_out[14][9][13] = xor_out[70][9][13] + xor_out[71][9][13] + xor_out[72][9][13] + xor_out[73][9][13] + xor_out[74][9][13];
assign sum_out[15][9][13] = xor_out[75][9][13] + xor_out[76][9][13] + xor_out[77][9][13] + xor_out[78][9][13] + xor_out[79][9][13];
assign sum_out[16][9][13] = xor_out[80][9][13] + xor_out[81][9][13] + xor_out[82][9][13] + xor_out[83][9][13] + xor_out[84][9][13];
assign sum_out[17][9][13] = xor_out[85][9][13] + xor_out[86][9][13] + xor_out[87][9][13] + xor_out[88][9][13] + xor_out[89][9][13];
assign sum_out[18][9][13] = xor_out[90][9][13] + xor_out[91][9][13] + xor_out[92][9][13] + xor_out[93][9][13] + xor_out[94][9][13];
assign sum_out[19][9][13] = xor_out[95][9][13] + xor_out[96][9][13] + xor_out[97][9][13] + xor_out[98][9][13] + xor_out[99][9][13];

assign sum_out[0][9][14] = xor_out[0][9][14] + xor_out[1][9][14] + xor_out[2][9][14] + xor_out[3][9][14] + xor_out[4][9][14];
assign sum_out[1][9][14] = xor_out[5][9][14] + xor_out[6][9][14] + xor_out[7][9][14] + xor_out[8][9][14] + xor_out[9][9][14];
assign sum_out[2][9][14] = xor_out[10][9][14] + xor_out[11][9][14] + xor_out[12][9][14] + xor_out[13][9][14] + xor_out[14][9][14];
assign sum_out[3][9][14] = xor_out[15][9][14] + xor_out[16][9][14] + xor_out[17][9][14] + xor_out[18][9][14] + xor_out[19][9][14];
assign sum_out[4][9][14] = xor_out[20][9][14] + xor_out[21][9][14] + xor_out[22][9][14] + xor_out[23][9][14] + xor_out[24][9][14];
assign sum_out[5][9][14] = xor_out[25][9][14] + xor_out[26][9][14] + xor_out[27][9][14] + xor_out[28][9][14] + xor_out[29][9][14];
assign sum_out[6][9][14] = xor_out[30][9][14] + xor_out[31][9][14] + xor_out[32][9][14] + xor_out[33][9][14] + xor_out[34][9][14];
assign sum_out[7][9][14] = xor_out[35][9][14] + xor_out[36][9][14] + xor_out[37][9][14] + xor_out[38][9][14] + xor_out[39][9][14];
assign sum_out[8][9][14] = xor_out[40][9][14] + xor_out[41][9][14] + xor_out[42][9][14] + xor_out[43][9][14] + xor_out[44][9][14];
assign sum_out[9][9][14] = xor_out[45][9][14] + xor_out[46][9][14] + xor_out[47][9][14] + xor_out[48][9][14] + xor_out[49][9][14];
assign sum_out[10][9][14] = xor_out[50][9][14] + xor_out[51][9][14] + xor_out[52][9][14] + xor_out[53][9][14] + xor_out[54][9][14];
assign sum_out[11][9][14] = xor_out[55][9][14] + xor_out[56][9][14] + xor_out[57][9][14] + xor_out[58][9][14] + xor_out[59][9][14];
assign sum_out[12][9][14] = xor_out[60][9][14] + xor_out[61][9][14] + xor_out[62][9][14] + xor_out[63][9][14] + xor_out[64][9][14];
assign sum_out[13][9][14] = xor_out[65][9][14] + xor_out[66][9][14] + xor_out[67][9][14] + xor_out[68][9][14] + xor_out[69][9][14];
assign sum_out[14][9][14] = xor_out[70][9][14] + xor_out[71][9][14] + xor_out[72][9][14] + xor_out[73][9][14] + xor_out[74][9][14];
assign sum_out[15][9][14] = xor_out[75][9][14] + xor_out[76][9][14] + xor_out[77][9][14] + xor_out[78][9][14] + xor_out[79][9][14];
assign sum_out[16][9][14] = xor_out[80][9][14] + xor_out[81][9][14] + xor_out[82][9][14] + xor_out[83][9][14] + xor_out[84][9][14];
assign sum_out[17][9][14] = xor_out[85][9][14] + xor_out[86][9][14] + xor_out[87][9][14] + xor_out[88][9][14] + xor_out[89][9][14];
assign sum_out[18][9][14] = xor_out[90][9][14] + xor_out[91][9][14] + xor_out[92][9][14] + xor_out[93][9][14] + xor_out[94][9][14];
assign sum_out[19][9][14] = xor_out[95][9][14] + xor_out[96][9][14] + xor_out[97][9][14] + xor_out[98][9][14] + xor_out[99][9][14];

assign sum_out[0][9][15] = xor_out[0][9][15] + xor_out[1][9][15] + xor_out[2][9][15] + xor_out[3][9][15] + xor_out[4][9][15];
assign sum_out[1][9][15] = xor_out[5][9][15] + xor_out[6][9][15] + xor_out[7][9][15] + xor_out[8][9][15] + xor_out[9][9][15];
assign sum_out[2][9][15] = xor_out[10][9][15] + xor_out[11][9][15] + xor_out[12][9][15] + xor_out[13][9][15] + xor_out[14][9][15];
assign sum_out[3][9][15] = xor_out[15][9][15] + xor_out[16][9][15] + xor_out[17][9][15] + xor_out[18][9][15] + xor_out[19][9][15];
assign sum_out[4][9][15] = xor_out[20][9][15] + xor_out[21][9][15] + xor_out[22][9][15] + xor_out[23][9][15] + xor_out[24][9][15];
assign sum_out[5][9][15] = xor_out[25][9][15] + xor_out[26][9][15] + xor_out[27][9][15] + xor_out[28][9][15] + xor_out[29][9][15];
assign sum_out[6][9][15] = xor_out[30][9][15] + xor_out[31][9][15] + xor_out[32][9][15] + xor_out[33][9][15] + xor_out[34][9][15];
assign sum_out[7][9][15] = xor_out[35][9][15] + xor_out[36][9][15] + xor_out[37][9][15] + xor_out[38][9][15] + xor_out[39][9][15];
assign sum_out[8][9][15] = xor_out[40][9][15] + xor_out[41][9][15] + xor_out[42][9][15] + xor_out[43][9][15] + xor_out[44][9][15];
assign sum_out[9][9][15] = xor_out[45][9][15] + xor_out[46][9][15] + xor_out[47][9][15] + xor_out[48][9][15] + xor_out[49][9][15];
assign sum_out[10][9][15] = xor_out[50][9][15] + xor_out[51][9][15] + xor_out[52][9][15] + xor_out[53][9][15] + xor_out[54][9][15];
assign sum_out[11][9][15] = xor_out[55][9][15] + xor_out[56][9][15] + xor_out[57][9][15] + xor_out[58][9][15] + xor_out[59][9][15];
assign sum_out[12][9][15] = xor_out[60][9][15] + xor_out[61][9][15] + xor_out[62][9][15] + xor_out[63][9][15] + xor_out[64][9][15];
assign sum_out[13][9][15] = xor_out[65][9][15] + xor_out[66][9][15] + xor_out[67][9][15] + xor_out[68][9][15] + xor_out[69][9][15];
assign sum_out[14][9][15] = xor_out[70][9][15] + xor_out[71][9][15] + xor_out[72][9][15] + xor_out[73][9][15] + xor_out[74][9][15];
assign sum_out[15][9][15] = xor_out[75][9][15] + xor_out[76][9][15] + xor_out[77][9][15] + xor_out[78][9][15] + xor_out[79][9][15];
assign sum_out[16][9][15] = xor_out[80][9][15] + xor_out[81][9][15] + xor_out[82][9][15] + xor_out[83][9][15] + xor_out[84][9][15];
assign sum_out[17][9][15] = xor_out[85][9][15] + xor_out[86][9][15] + xor_out[87][9][15] + xor_out[88][9][15] + xor_out[89][9][15];
assign sum_out[18][9][15] = xor_out[90][9][15] + xor_out[91][9][15] + xor_out[92][9][15] + xor_out[93][9][15] + xor_out[94][9][15];
assign sum_out[19][9][15] = xor_out[95][9][15] + xor_out[96][9][15] + xor_out[97][9][15] + xor_out[98][9][15] + xor_out[99][9][15];

assign sum_out[0][9][16] = xor_out[0][9][16] + xor_out[1][9][16] + xor_out[2][9][16] + xor_out[3][9][16] + xor_out[4][9][16];
assign sum_out[1][9][16] = xor_out[5][9][16] + xor_out[6][9][16] + xor_out[7][9][16] + xor_out[8][9][16] + xor_out[9][9][16];
assign sum_out[2][9][16] = xor_out[10][9][16] + xor_out[11][9][16] + xor_out[12][9][16] + xor_out[13][9][16] + xor_out[14][9][16];
assign sum_out[3][9][16] = xor_out[15][9][16] + xor_out[16][9][16] + xor_out[17][9][16] + xor_out[18][9][16] + xor_out[19][9][16];
assign sum_out[4][9][16] = xor_out[20][9][16] + xor_out[21][9][16] + xor_out[22][9][16] + xor_out[23][9][16] + xor_out[24][9][16];
assign sum_out[5][9][16] = xor_out[25][9][16] + xor_out[26][9][16] + xor_out[27][9][16] + xor_out[28][9][16] + xor_out[29][9][16];
assign sum_out[6][9][16] = xor_out[30][9][16] + xor_out[31][9][16] + xor_out[32][9][16] + xor_out[33][9][16] + xor_out[34][9][16];
assign sum_out[7][9][16] = xor_out[35][9][16] + xor_out[36][9][16] + xor_out[37][9][16] + xor_out[38][9][16] + xor_out[39][9][16];
assign sum_out[8][9][16] = xor_out[40][9][16] + xor_out[41][9][16] + xor_out[42][9][16] + xor_out[43][9][16] + xor_out[44][9][16];
assign sum_out[9][9][16] = xor_out[45][9][16] + xor_out[46][9][16] + xor_out[47][9][16] + xor_out[48][9][16] + xor_out[49][9][16];
assign sum_out[10][9][16] = xor_out[50][9][16] + xor_out[51][9][16] + xor_out[52][9][16] + xor_out[53][9][16] + xor_out[54][9][16];
assign sum_out[11][9][16] = xor_out[55][9][16] + xor_out[56][9][16] + xor_out[57][9][16] + xor_out[58][9][16] + xor_out[59][9][16];
assign sum_out[12][9][16] = xor_out[60][9][16] + xor_out[61][9][16] + xor_out[62][9][16] + xor_out[63][9][16] + xor_out[64][9][16];
assign sum_out[13][9][16] = xor_out[65][9][16] + xor_out[66][9][16] + xor_out[67][9][16] + xor_out[68][9][16] + xor_out[69][9][16];
assign sum_out[14][9][16] = xor_out[70][9][16] + xor_out[71][9][16] + xor_out[72][9][16] + xor_out[73][9][16] + xor_out[74][9][16];
assign sum_out[15][9][16] = xor_out[75][9][16] + xor_out[76][9][16] + xor_out[77][9][16] + xor_out[78][9][16] + xor_out[79][9][16];
assign sum_out[16][9][16] = xor_out[80][9][16] + xor_out[81][9][16] + xor_out[82][9][16] + xor_out[83][9][16] + xor_out[84][9][16];
assign sum_out[17][9][16] = xor_out[85][9][16] + xor_out[86][9][16] + xor_out[87][9][16] + xor_out[88][9][16] + xor_out[89][9][16];
assign sum_out[18][9][16] = xor_out[90][9][16] + xor_out[91][9][16] + xor_out[92][9][16] + xor_out[93][9][16] + xor_out[94][9][16];
assign sum_out[19][9][16] = xor_out[95][9][16] + xor_out[96][9][16] + xor_out[97][9][16] + xor_out[98][9][16] + xor_out[99][9][16];

assign sum_out[0][9][17] = xor_out[0][9][17] + xor_out[1][9][17] + xor_out[2][9][17] + xor_out[3][9][17] + xor_out[4][9][17];
assign sum_out[1][9][17] = xor_out[5][9][17] + xor_out[6][9][17] + xor_out[7][9][17] + xor_out[8][9][17] + xor_out[9][9][17];
assign sum_out[2][9][17] = xor_out[10][9][17] + xor_out[11][9][17] + xor_out[12][9][17] + xor_out[13][9][17] + xor_out[14][9][17];
assign sum_out[3][9][17] = xor_out[15][9][17] + xor_out[16][9][17] + xor_out[17][9][17] + xor_out[18][9][17] + xor_out[19][9][17];
assign sum_out[4][9][17] = xor_out[20][9][17] + xor_out[21][9][17] + xor_out[22][9][17] + xor_out[23][9][17] + xor_out[24][9][17];
assign sum_out[5][9][17] = xor_out[25][9][17] + xor_out[26][9][17] + xor_out[27][9][17] + xor_out[28][9][17] + xor_out[29][9][17];
assign sum_out[6][9][17] = xor_out[30][9][17] + xor_out[31][9][17] + xor_out[32][9][17] + xor_out[33][9][17] + xor_out[34][9][17];
assign sum_out[7][9][17] = xor_out[35][9][17] + xor_out[36][9][17] + xor_out[37][9][17] + xor_out[38][9][17] + xor_out[39][9][17];
assign sum_out[8][9][17] = xor_out[40][9][17] + xor_out[41][9][17] + xor_out[42][9][17] + xor_out[43][9][17] + xor_out[44][9][17];
assign sum_out[9][9][17] = xor_out[45][9][17] + xor_out[46][9][17] + xor_out[47][9][17] + xor_out[48][9][17] + xor_out[49][9][17];
assign sum_out[10][9][17] = xor_out[50][9][17] + xor_out[51][9][17] + xor_out[52][9][17] + xor_out[53][9][17] + xor_out[54][9][17];
assign sum_out[11][9][17] = xor_out[55][9][17] + xor_out[56][9][17] + xor_out[57][9][17] + xor_out[58][9][17] + xor_out[59][9][17];
assign sum_out[12][9][17] = xor_out[60][9][17] + xor_out[61][9][17] + xor_out[62][9][17] + xor_out[63][9][17] + xor_out[64][9][17];
assign sum_out[13][9][17] = xor_out[65][9][17] + xor_out[66][9][17] + xor_out[67][9][17] + xor_out[68][9][17] + xor_out[69][9][17];
assign sum_out[14][9][17] = xor_out[70][9][17] + xor_out[71][9][17] + xor_out[72][9][17] + xor_out[73][9][17] + xor_out[74][9][17];
assign sum_out[15][9][17] = xor_out[75][9][17] + xor_out[76][9][17] + xor_out[77][9][17] + xor_out[78][9][17] + xor_out[79][9][17];
assign sum_out[16][9][17] = xor_out[80][9][17] + xor_out[81][9][17] + xor_out[82][9][17] + xor_out[83][9][17] + xor_out[84][9][17];
assign sum_out[17][9][17] = xor_out[85][9][17] + xor_out[86][9][17] + xor_out[87][9][17] + xor_out[88][9][17] + xor_out[89][9][17];
assign sum_out[18][9][17] = xor_out[90][9][17] + xor_out[91][9][17] + xor_out[92][9][17] + xor_out[93][9][17] + xor_out[94][9][17];
assign sum_out[19][9][17] = xor_out[95][9][17] + xor_out[96][9][17] + xor_out[97][9][17] + xor_out[98][9][17] + xor_out[99][9][17];

assign sum_out[0][9][18] = xor_out[0][9][18] + xor_out[1][9][18] + xor_out[2][9][18] + xor_out[3][9][18] + xor_out[4][9][18];
assign sum_out[1][9][18] = xor_out[5][9][18] + xor_out[6][9][18] + xor_out[7][9][18] + xor_out[8][9][18] + xor_out[9][9][18];
assign sum_out[2][9][18] = xor_out[10][9][18] + xor_out[11][9][18] + xor_out[12][9][18] + xor_out[13][9][18] + xor_out[14][9][18];
assign sum_out[3][9][18] = xor_out[15][9][18] + xor_out[16][9][18] + xor_out[17][9][18] + xor_out[18][9][18] + xor_out[19][9][18];
assign sum_out[4][9][18] = xor_out[20][9][18] + xor_out[21][9][18] + xor_out[22][9][18] + xor_out[23][9][18] + xor_out[24][9][18];
assign sum_out[5][9][18] = xor_out[25][9][18] + xor_out[26][9][18] + xor_out[27][9][18] + xor_out[28][9][18] + xor_out[29][9][18];
assign sum_out[6][9][18] = xor_out[30][9][18] + xor_out[31][9][18] + xor_out[32][9][18] + xor_out[33][9][18] + xor_out[34][9][18];
assign sum_out[7][9][18] = xor_out[35][9][18] + xor_out[36][9][18] + xor_out[37][9][18] + xor_out[38][9][18] + xor_out[39][9][18];
assign sum_out[8][9][18] = xor_out[40][9][18] + xor_out[41][9][18] + xor_out[42][9][18] + xor_out[43][9][18] + xor_out[44][9][18];
assign sum_out[9][9][18] = xor_out[45][9][18] + xor_out[46][9][18] + xor_out[47][9][18] + xor_out[48][9][18] + xor_out[49][9][18];
assign sum_out[10][9][18] = xor_out[50][9][18] + xor_out[51][9][18] + xor_out[52][9][18] + xor_out[53][9][18] + xor_out[54][9][18];
assign sum_out[11][9][18] = xor_out[55][9][18] + xor_out[56][9][18] + xor_out[57][9][18] + xor_out[58][9][18] + xor_out[59][9][18];
assign sum_out[12][9][18] = xor_out[60][9][18] + xor_out[61][9][18] + xor_out[62][9][18] + xor_out[63][9][18] + xor_out[64][9][18];
assign sum_out[13][9][18] = xor_out[65][9][18] + xor_out[66][9][18] + xor_out[67][9][18] + xor_out[68][9][18] + xor_out[69][9][18];
assign sum_out[14][9][18] = xor_out[70][9][18] + xor_out[71][9][18] + xor_out[72][9][18] + xor_out[73][9][18] + xor_out[74][9][18];
assign sum_out[15][9][18] = xor_out[75][9][18] + xor_out[76][9][18] + xor_out[77][9][18] + xor_out[78][9][18] + xor_out[79][9][18];
assign sum_out[16][9][18] = xor_out[80][9][18] + xor_out[81][9][18] + xor_out[82][9][18] + xor_out[83][9][18] + xor_out[84][9][18];
assign sum_out[17][9][18] = xor_out[85][9][18] + xor_out[86][9][18] + xor_out[87][9][18] + xor_out[88][9][18] + xor_out[89][9][18];
assign sum_out[18][9][18] = xor_out[90][9][18] + xor_out[91][9][18] + xor_out[92][9][18] + xor_out[93][9][18] + xor_out[94][9][18];
assign sum_out[19][9][18] = xor_out[95][9][18] + xor_out[96][9][18] + xor_out[97][9][18] + xor_out[98][9][18] + xor_out[99][9][18];

assign sum_out[0][9][19] = xor_out[0][9][19] + xor_out[1][9][19] + xor_out[2][9][19] + xor_out[3][9][19] + xor_out[4][9][19];
assign sum_out[1][9][19] = xor_out[5][9][19] + xor_out[6][9][19] + xor_out[7][9][19] + xor_out[8][9][19] + xor_out[9][9][19];
assign sum_out[2][9][19] = xor_out[10][9][19] + xor_out[11][9][19] + xor_out[12][9][19] + xor_out[13][9][19] + xor_out[14][9][19];
assign sum_out[3][9][19] = xor_out[15][9][19] + xor_out[16][9][19] + xor_out[17][9][19] + xor_out[18][9][19] + xor_out[19][9][19];
assign sum_out[4][9][19] = xor_out[20][9][19] + xor_out[21][9][19] + xor_out[22][9][19] + xor_out[23][9][19] + xor_out[24][9][19];
assign sum_out[5][9][19] = xor_out[25][9][19] + xor_out[26][9][19] + xor_out[27][9][19] + xor_out[28][9][19] + xor_out[29][9][19];
assign sum_out[6][9][19] = xor_out[30][9][19] + xor_out[31][9][19] + xor_out[32][9][19] + xor_out[33][9][19] + xor_out[34][9][19];
assign sum_out[7][9][19] = xor_out[35][9][19] + xor_out[36][9][19] + xor_out[37][9][19] + xor_out[38][9][19] + xor_out[39][9][19];
assign sum_out[8][9][19] = xor_out[40][9][19] + xor_out[41][9][19] + xor_out[42][9][19] + xor_out[43][9][19] + xor_out[44][9][19];
assign sum_out[9][9][19] = xor_out[45][9][19] + xor_out[46][9][19] + xor_out[47][9][19] + xor_out[48][9][19] + xor_out[49][9][19];
assign sum_out[10][9][19] = xor_out[50][9][19] + xor_out[51][9][19] + xor_out[52][9][19] + xor_out[53][9][19] + xor_out[54][9][19];
assign sum_out[11][9][19] = xor_out[55][9][19] + xor_out[56][9][19] + xor_out[57][9][19] + xor_out[58][9][19] + xor_out[59][9][19];
assign sum_out[12][9][19] = xor_out[60][9][19] + xor_out[61][9][19] + xor_out[62][9][19] + xor_out[63][9][19] + xor_out[64][9][19];
assign sum_out[13][9][19] = xor_out[65][9][19] + xor_out[66][9][19] + xor_out[67][9][19] + xor_out[68][9][19] + xor_out[69][9][19];
assign sum_out[14][9][19] = xor_out[70][9][19] + xor_out[71][9][19] + xor_out[72][9][19] + xor_out[73][9][19] + xor_out[74][9][19];
assign sum_out[15][9][19] = xor_out[75][9][19] + xor_out[76][9][19] + xor_out[77][9][19] + xor_out[78][9][19] + xor_out[79][9][19];
assign sum_out[16][9][19] = xor_out[80][9][19] + xor_out[81][9][19] + xor_out[82][9][19] + xor_out[83][9][19] + xor_out[84][9][19];
assign sum_out[17][9][19] = xor_out[85][9][19] + xor_out[86][9][19] + xor_out[87][9][19] + xor_out[88][9][19] + xor_out[89][9][19];
assign sum_out[18][9][19] = xor_out[90][9][19] + xor_out[91][9][19] + xor_out[92][9][19] + xor_out[93][9][19] + xor_out[94][9][19];
assign sum_out[19][9][19] = xor_out[95][9][19] + xor_out[96][9][19] + xor_out[97][9][19] + xor_out[98][9][19] + xor_out[99][9][19];

assign sum_out[0][9][20] = xor_out[0][9][20] + xor_out[1][9][20] + xor_out[2][9][20] + xor_out[3][9][20] + xor_out[4][9][20];
assign sum_out[1][9][20] = xor_out[5][9][20] + xor_out[6][9][20] + xor_out[7][9][20] + xor_out[8][9][20] + xor_out[9][9][20];
assign sum_out[2][9][20] = xor_out[10][9][20] + xor_out[11][9][20] + xor_out[12][9][20] + xor_out[13][9][20] + xor_out[14][9][20];
assign sum_out[3][9][20] = xor_out[15][9][20] + xor_out[16][9][20] + xor_out[17][9][20] + xor_out[18][9][20] + xor_out[19][9][20];
assign sum_out[4][9][20] = xor_out[20][9][20] + xor_out[21][9][20] + xor_out[22][9][20] + xor_out[23][9][20] + xor_out[24][9][20];
assign sum_out[5][9][20] = xor_out[25][9][20] + xor_out[26][9][20] + xor_out[27][9][20] + xor_out[28][9][20] + xor_out[29][9][20];
assign sum_out[6][9][20] = xor_out[30][9][20] + xor_out[31][9][20] + xor_out[32][9][20] + xor_out[33][9][20] + xor_out[34][9][20];
assign sum_out[7][9][20] = xor_out[35][9][20] + xor_out[36][9][20] + xor_out[37][9][20] + xor_out[38][9][20] + xor_out[39][9][20];
assign sum_out[8][9][20] = xor_out[40][9][20] + xor_out[41][9][20] + xor_out[42][9][20] + xor_out[43][9][20] + xor_out[44][9][20];
assign sum_out[9][9][20] = xor_out[45][9][20] + xor_out[46][9][20] + xor_out[47][9][20] + xor_out[48][9][20] + xor_out[49][9][20];
assign sum_out[10][9][20] = xor_out[50][9][20] + xor_out[51][9][20] + xor_out[52][9][20] + xor_out[53][9][20] + xor_out[54][9][20];
assign sum_out[11][9][20] = xor_out[55][9][20] + xor_out[56][9][20] + xor_out[57][9][20] + xor_out[58][9][20] + xor_out[59][9][20];
assign sum_out[12][9][20] = xor_out[60][9][20] + xor_out[61][9][20] + xor_out[62][9][20] + xor_out[63][9][20] + xor_out[64][9][20];
assign sum_out[13][9][20] = xor_out[65][9][20] + xor_out[66][9][20] + xor_out[67][9][20] + xor_out[68][9][20] + xor_out[69][9][20];
assign sum_out[14][9][20] = xor_out[70][9][20] + xor_out[71][9][20] + xor_out[72][9][20] + xor_out[73][9][20] + xor_out[74][9][20];
assign sum_out[15][9][20] = xor_out[75][9][20] + xor_out[76][9][20] + xor_out[77][9][20] + xor_out[78][9][20] + xor_out[79][9][20];
assign sum_out[16][9][20] = xor_out[80][9][20] + xor_out[81][9][20] + xor_out[82][9][20] + xor_out[83][9][20] + xor_out[84][9][20];
assign sum_out[17][9][20] = xor_out[85][9][20] + xor_out[86][9][20] + xor_out[87][9][20] + xor_out[88][9][20] + xor_out[89][9][20];
assign sum_out[18][9][20] = xor_out[90][9][20] + xor_out[91][9][20] + xor_out[92][9][20] + xor_out[93][9][20] + xor_out[94][9][20];
assign sum_out[19][9][20] = xor_out[95][9][20] + xor_out[96][9][20] + xor_out[97][9][20] + xor_out[98][9][20] + xor_out[99][9][20];

assign sum_out[0][9][21] = xor_out[0][9][21] + xor_out[1][9][21] + xor_out[2][9][21] + xor_out[3][9][21] + xor_out[4][9][21];
assign sum_out[1][9][21] = xor_out[5][9][21] + xor_out[6][9][21] + xor_out[7][9][21] + xor_out[8][9][21] + xor_out[9][9][21];
assign sum_out[2][9][21] = xor_out[10][9][21] + xor_out[11][9][21] + xor_out[12][9][21] + xor_out[13][9][21] + xor_out[14][9][21];
assign sum_out[3][9][21] = xor_out[15][9][21] + xor_out[16][9][21] + xor_out[17][9][21] + xor_out[18][9][21] + xor_out[19][9][21];
assign sum_out[4][9][21] = xor_out[20][9][21] + xor_out[21][9][21] + xor_out[22][9][21] + xor_out[23][9][21] + xor_out[24][9][21];
assign sum_out[5][9][21] = xor_out[25][9][21] + xor_out[26][9][21] + xor_out[27][9][21] + xor_out[28][9][21] + xor_out[29][9][21];
assign sum_out[6][9][21] = xor_out[30][9][21] + xor_out[31][9][21] + xor_out[32][9][21] + xor_out[33][9][21] + xor_out[34][9][21];
assign sum_out[7][9][21] = xor_out[35][9][21] + xor_out[36][9][21] + xor_out[37][9][21] + xor_out[38][9][21] + xor_out[39][9][21];
assign sum_out[8][9][21] = xor_out[40][9][21] + xor_out[41][9][21] + xor_out[42][9][21] + xor_out[43][9][21] + xor_out[44][9][21];
assign sum_out[9][9][21] = xor_out[45][9][21] + xor_out[46][9][21] + xor_out[47][9][21] + xor_out[48][9][21] + xor_out[49][9][21];
assign sum_out[10][9][21] = xor_out[50][9][21] + xor_out[51][9][21] + xor_out[52][9][21] + xor_out[53][9][21] + xor_out[54][9][21];
assign sum_out[11][9][21] = xor_out[55][9][21] + xor_out[56][9][21] + xor_out[57][9][21] + xor_out[58][9][21] + xor_out[59][9][21];
assign sum_out[12][9][21] = xor_out[60][9][21] + xor_out[61][9][21] + xor_out[62][9][21] + xor_out[63][9][21] + xor_out[64][9][21];
assign sum_out[13][9][21] = xor_out[65][9][21] + xor_out[66][9][21] + xor_out[67][9][21] + xor_out[68][9][21] + xor_out[69][9][21];
assign sum_out[14][9][21] = xor_out[70][9][21] + xor_out[71][9][21] + xor_out[72][9][21] + xor_out[73][9][21] + xor_out[74][9][21];
assign sum_out[15][9][21] = xor_out[75][9][21] + xor_out[76][9][21] + xor_out[77][9][21] + xor_out[78][9][21] + xor_out[79][9][21];
assign sum_out[16][9][21] = xor_out[80][9][21] + xor_out[81][9][21] + xor_out[82][9][21] + xor_out[83][9][21] + xor_out[84][9][21];
assign sum_out[17][9][21] = xor_out[85][9][21] + xor_out[86][9][21] + xor_out[87][9][21] + xor_out[88][9][21] + xor_out[89][9][21];
assign sum_out[18][9][21] = xor_out[90][9][21] + xor_out[91][9][21] + xor_out[92][9][21] + xor_out[93][9][21] + xor_out[94][9][21];
assign sum_out[19][9][21] = xor_out[95][9][21] + xor_out[96][9][21] + xor_out[97][9][21] + xor_out[98][9][21] + xor_out[99][9][21];

assign sum_out[0][9][22] = xor_out[0][9][22] + xor_out[1][9][22] + xor_out[2][9][22] + xor_out[3][9][22] + xor_out[4][9][22];
assign sum_out[1][9][22] = xor_out[5][9][22] + xor_out[6][9][22] + xor_out[7][9][22] + xor_out[8][9][22] + xor_out[9][9][22];
assign sum_out[2][9][22] = xor_out[10][9][22] + xor_out[11][9][22] + xor_out[12][9][22] + xor_out[13][9][22] + xor_out[14][9][22];
assign sum_out[3][9][22] = xor_out[15][9][22] + xor_out[16][9][22] + xor_out[17][9][22] + xor_out[18][9][22] + xor_out[19][9][22];
assign sum_out[4][9][22] = xor_out[20][9][22] + xor_out[21][9][22] + xor_out[22][9][22] + xor_out[23][9][22] + xor_out[24][9][22];
assign sum_out[5][9][22] = xor_out[25][9][22] + xor_out[26][9][22] + xor_out[27][9][22] + xor_out[28][9][22] + xor_out[29][9][22];
assign sum_out[6][9][22] = xor_out[30][9][22] + xor_out[31][9][22] + xor_out[32][9][22] + xor_out[33][9][22] + xor_out[34][9][22];
assign sum_out[7][9][22] = xor_out[35][9][22] + xor_out[36][9][22] + xor_out[37][9][22] + xor_out[38][9][22] + xor_out[39][9][22];
assign sum_out[8][9][22] = xor_out[40][9][22] + xor_out[41][9][22] + xor_out[42][9][22] + xor_out[43][9][22] + xor_out[44][9][22];
assign sum_out[9][9][22] = xor_out[45][9][22] + xor_out[46][9][22] + xor_out[47][9][22] + xor_out[48][9][22] + xor_out[49][9][22];
assign sum_out[10][9][22] = xor_out[50][9][22] + xor_out[51][9][22] + xor_out[52][9][22] + xor_out[53][9][22] + xor_out[54][9][22];
assign sum_out[11][9][22] = xor_out[55][9][22] + xor_out[56][9][22] + xor_out[57][9][22] + xor_out[58][9][22] + xor_out[59][9][22];
assign sum_out[12][9][22] = xor_out[60][9][22] + xor_out[61][9][22] + xor_out[62][9][22] + xor_out[63][9][22] + xor_out[64][9][22];
assign sum_out[13][9][22] = xor_out[65][9][22] + xor_out[66][9][22] + xor_out[67][9][22] + xor_out[68][9][22] + xor_out[69][9][22];
assign sum_out[14][9][22] = xor_out[70][9][22] + xor_out[71][9][22] + xor_out[72][9][22] + xor_out[73][9][22] + xor_out[74][9][22];
assign sum_out[15][9][22] = xor_out[75][9][22] + xor_out[76][9][22] + xor_out[77][9][22] + xor_out[78][9][22] + xor_out[79][9][22];
assign sum_out[16][9][22] = xor_out[80][9][22] + xor_out[81][9][22] + xor_out[82][9][22] + xor_out[83][9][22] + xor_out[84][9][22];
assign sum_out[17][9][22] = xor_out[85][9][22] + xor_out[86][9][22] + xor_out[87][9][22] + xor_out[88][9][22] + xor_out[89][9][22];
assign sum_out[18][9][22] = xor_out[90][9][22] + xor_out[91][9][22] + xor_out[92][9][22] + xor_out[93][9][22] + xor_out[94][9][22];
assign sum_out[19][9][22] = xor_out[95][9][22] + xor_out[96][9][22] + xor_out[97][9][22] + xor_out[98][9][22] + xor_out[99][9][22];

assign sum_out[0][9][23] = xor_out[0][9][23] + xor_out[1][9][23] + xor_out[2][9][23] + xor_out[3][9][23] + xor_out[4][9][23];
assign sum_out[1][9][23] = xor_out[5][9][23] + xor_out[6][9][23] + xor_out[7][9][23] + xor_out[8][9][23] + xor_out[9][9][23];
assign sum_out[2][9][23] = xor_out[10][9][23] + xor_out[11][9][23] + xor_out[12][9][23] + xor_out[13][9][23] + xor_out[14][9][23];
assign sum_out[3][9][23] = xor_out[15][9][23] + xor_out[16][9][23] + xor_out[17][9][23] + xor_out[18][9][23] + xor_out[19][9][23];
assign sum_out[4][9][23] = xor_out[20][9][23] + xor_out[21][9][23] + xor_out[22][9][23] + xor_out[23][9][23] + xor_out[24][9][23];
assign sum_out[5][9][23] = xor_out[25][9][23] + xor_out[26][9][23] + xor_out[27][9][23] + xor_out[28][9][23] + xor_out[29][9][23];
assign sum_out[6][9][23] = xor_out[30][9][23] + xor_out[31][9][23] + xor_out[32][9][23] + xor_out[33][9][23] + xor_out[34][9][23];
assign sum_out[7][9][23] = xor_out[35][9][23] + xor_out[36][9][23] + xor_out[37][9][23] + xor_out[38][9][23] + xor_out[39][9][23];
assign sum_out[8][9][23] = xor_out[40][9][23] + xor_out[41][9][23] + xor_out[42][9][23] + xor_out[43][9][23] + xor_out[44][9][23];
assign sum_out[9][9][23] = xor_out[45][9][23] + xor_out[46][9][23] + xor_out[47][9][23] + xor_out[48][9][23] + xor_out[49][9][23];
assign sum_out[10][9][23] = xor_out[50][9][23] + xor_out[51][9][23] + xor_out[52][9][23] + xor_out[53][9][23] + xor_out[54][9][23];
assign sum_out[11][9][23] = xor_out[55][9][23] + xor_out[56][9][23] + xor_out[57][9][23] + xor_out[58][9][23] + xor_out[59][9][23];
assign sum_out[12][9][23] = xor_out[60][9][23] + xor_out[61][9][23] + xor_out[62][9][23] + xor_out[63][9][23] + xor_out[64][9][23];
assign sum_out[13][9][23] = xor_out[65][9][23] + xor_out[66][9][23] + xor_out[67][9][23] + xor_out[68][9][23] + xor_out[69][9][23];
assign sum_out[14][9][23] = xor_out[70][9][23] + xor_out[71][9][23] + xor_out[72][9][23] + xor_out[73][9][23] + xor_out[74][9][23];
assign sum_out[15][9][23] = xor_out[75][9][23] + xor_out[76][9][23] + xor_out[77][9][23] + xor_out[78][9][23] + xor_out[79][9][23];
assign sum_out[16][9][23] = xor_out[80][9][23] + xor_out[81][9][23] + xor_out[82][9][23] + xor_out[83][9][23] + xor_out[84][9][23];
assign sum_out[17][9][23] = xor_out[85][9][23] + xor_out[86][9][23] + xor_out[87][9][23] + xor_out[88][9][23] + xor_out[89][9][23];
assign sum_out[18][9][23] = xor_out[90][9][23] + xor_out[91][9][23] + xor_out[92][9][23] + xor_out[93][9][23] + xor_out[94][9][23];
assign sum_out[19][9][23] = xor_out[95][9][23] + xor_out[96][9][23] + xor_out[97][9][23] + xor_out[98][9][23] + xor_out[99][9][23];

assign sum_out[0][10][0] = xor_out[0][10][0] + xor_out[1][10][0] + xor_out[2][10][0] + xor_out[3][10][0] + xor_out[4][10][0];
assign sum_out[1][10][0] = xor_out[5][10][0] + xor_out[6][10][0] + xor_out[7][10][0] + xor_out[8][10][0] + xor_out[9][10][0];
assign sum_out[2][10][0] = xor_out[10][10][0] + xor_out[11][10][0] + xor_out[12][10][0] + xor_out[13][10][0] + xor_out[14][10][0];
assign sum_out[3][10][0] = xor_out[15][10][0] + xor_out[16][10][0] + xor_out[17][10][0] + xor_out[18][10][0] + xor_out[19][10][0];
assign sum_out[4][10][0] = xor_out[20][10][0] + xor_out[21][10][0] + xor_out[22][10][0] + xor_out[23][10][0] + xor_out[24][10][0];
assign sum_out[5][10][0] = xor_out[25][10][0] + xor_out[26][10][0] + xor_out[27][10][0] + xor_out[28][10][0] + xor_out[29][10][0];
assign sum_out[6][10][0] = xor_out[30][10][0] + xor_out[31][10][0] + xor_out[32][10][0] + xor_out[33][10][0] + xor_out[34][10][0];
assign sum_out[7][10][0] = xor_out[35][10][0] + xor_out[36][10][0] + xor_out[37][10][0] + xor_out[38][10][0] + xor_out[39][10][0];
assign sum_out[8][10][0] = xor_out[40][10][0] + xor_out[41][10][0] + xor_out[42][10][0] + xor_out[43][10][0] + xor_out[44][10][0];
assign sum_out[9][10][0] = xor_out[45][10][0] + xor_out[46][10][0] + xor_out[47][10][0] + xor_out[48][10][0] + xor_out[49][10][0];
assign sum_out[10][10][0] = xor_out[50][10][0] + xor_out[51][10][0] + xor_out[52][10][0] + xor_out[53][10][0] + xor_out[54][10][0];
assign sum_out[11][10][0] = xor_out[55][10][0] + xor_out[56][10][0] + xor_out[57][10][0] + xor_out[58][10][0] + xor_out[59][10][0];
assign sum_out[12][10][0] = xor_out[60][10][0] + xor_out[61][10][0] + xor_out[62][10][0] + xor_out[63][10][0] + xor_out[64][10][0];
assign sum_out[13][10][0] = xor_out[65][10][0] + xor_out[66][10][0] + xor_out[67][10][0] + xor_out[68][10][0] + xor_out[69][10][0];
assign sum_out[14][10][0] = xor_out[70][10][0] + xor_out[71][10][0] + xor_out[72][10][0] + xor_out[73][10][0] + xor_out[74][10][0];
assign sum_out[15][10][0] = xor_out[75][10][0] + xor_out[76][10][0] + xor_out[77][10][0] + xor_out[78][10][0] + xor_out[79][10][0];
assign sum_out[16][10][0] = xor_out[80][10][0] + xor_out[81][10][0] + xor_out[82][10][0] + xor_out[83][10][0] + xor_out[84][10][0];
assign sum_out[17][10][0] = xor_out[85][10][0] + xor_out[86][10][0] + xor_out[87][10][0] + xor_out[88][10][0] + xor_out[89][10][0];
assign sum_out[18][10][0] = xor_out[90][10][0] + xor_out[91][10][0] + xor_out[92][10][0] + xor_out[93][10][0] + xor_out[94][10][0];
assign sum_out[19][10][0] = xor_out[95][10][0] + xor_out[96][10][0] + xor_out[97][10][0] + xor_out[98][10][0] + xor_out[99][10][0];

assign sum_out[0][10][1] = xor_out[0][10][1] + xor_out[1][10][1] + xor_out[2][10][1] + xor_out[3][10][1] + xor_out[4][10][1];
assign sum_out[1][10][1] = xor_out[5][10][1] + xor_out[6][10][1] + xor_out[7][10][1] + xor_out[8][10][1] + xor_out[9][10][1];
assign sum_out[2][10][1] = xor_out[10][10][1] + xor_out[11][10][1] + xor_out[12][10][1] + xor_out[13][10][1] + xor_out[14][10][1];
assign sum_out[3][10][1] = xor_out[15][10][1] + xor_out[16][10][1] + xor_out[17][10][1] + xor_out[18][10][1] + xor_out[19][10][1];
assign sum_out[4][10][1] = xor_out[20][10][1] + xor_out[21][10][1] + xor_out[22][10][1] + xor_out[23][10][1] + xor_out[24][10][1];
assign sum_out[5][10][1] = xor_out[25][10][1] + xor_out[26][10][1] + xor_out[27][10][1] + xor_out[28][10][1] + xor_out[29][10][1];
assign sum_out[6][10][1] = xor_out[30][10][1] + xor_out[31][10][1] + xor_out[32][10][1] + xor_out[33][10][1] + xor_out[34][10][1];
assign sum_out[7][10][1] = xor_out[35][10][1] + xor_out[36][10][1] + xor_out[37][10][1] + xor_out[38][10][1] + xor_out[39][10][1];
assign sum_out[8][10][1] = xor_out[40][10][1] + xor_out[41][10][1] + xor_out[42][10][1] + xor_out[43][10][1] + xor_out[44][10][1];
assign sum_out[9][10][1] = xor_out[45][10][1] + xor_out[46][10][1] + xor_out[47][10][1] + xor_out[48][10][1] + xor_out[49][10][1];
assign sum_out[10][10][1] = xor_out[50][10][1] + xor_out[51][10][1] + xor_out[52][10][1] + xor_out[53][10][1] + xor_out[54][10][1];
assign sum_out[11][10][1] = xor_out[55][10][1] + xor_out[56][10][1] + xor_out[57][10][1] + xor_out[58][10][1] + xor_out[59][10][1];
assign sum_out[12][10][1] = xor_out[60][10][1] + xor_out[61][10][1] + xor_out[62][10][1] + xor_out[63][10][1] + xor_out[64][10][1];
assign sum_out[13][10][1] = xor_out[65][10][1] + xor_out[66][10][1] + xor_out[67][10][1] + xor_out[68][10][1] + xor_out[69][10][1];
assign sum_out[14][10][1] = xor_out[70][10][1] + xor_out[71][10][1] + xor_out[72][10][1] + xor_out[73][10][1] + xor_out[74][10][1];
assign sum_out[15][10][1] = xor_out[75][10][1] + xor_out[76][10][1] + xor_out[77][10][1] + xor_out[78][10][1] + xor_out[79][10][1];
assign sum_out[16][10][1] = xor_out[80][10][1] + xor_out[81][10][1] + xor_out[82][10][1] + xor_out[83][10][1] + xor_out[84][10][1];
assign sum_out[17][10][1] = xor_out[85][10][1] + xor_out[86][10][1] + xor_out[87][10][1] + xor_out[88][10][1] + xor_out[89][10][1];
assign sum_out[18][10][1] = xor_out[90][10][1] + xor_out[91][10][1] + xor_out[92][10][1] + xor_out[93][10][1] + xor_out[94][10][1];
assign sum_out[19][10][1] = xor_out[95][10][1] + xor_out[96][10][1] + xor_out[97][10][1] + xor_out[98][10][1] + xor_out[99][10][1];

assign sum_out[0][10][2] = xor_out[0][10][2] + xor_out[1][10][2] + xor_out[2][10][2] + xor_out[3][10][2] + xor_out[4][10][2];
assign sum_out[1][10][2] = xor_out[5][10][2] + xor_out[6][10][2] + xor_out[7][10][2] + xor_out[8][10][2] + xor_out[9][10][2];
assign sum_out[2][10][2] = xor_out[10][10][2] + xor_out[11][10][2] + xor_out[12][10][2] + xor_out[13][10][2] + xor_out[14][10][2];
assign sum_out[3][10][2] = xor_out[15][10][2] + xor_out[16][10][2] + xor_out[17][10][2] + xor_out[18][10][2] + xor_out[19][10][2];
assign sum_out[4][10][2] = xor_out[20][10][2] + xor_out[21][10][2] + xor_out[22][10][2] + xor_out[23][10][2] + xor_out[24][10][2];
assign sum_out[5][10][2] = xor_out[25][10][2] + xor_out[26][10][2] + xor_out[27][10][2] + xor_out[28][10][2] + xor_out[29][10][2];
assign sum_out[6][10][2] = xor_out[30][10][2] + xor_out[31][10][2] + xor_out[32][10][2] + xor_out[33][10][2] + xor_out[34][10][2];
assign sum_out[7][10][2] = xor_out[35][10][2] + xor_out[36][10][2] + xor_out[37][10][2] + xor_out[38][10][2] + xor_out[39][10][2];
assign sum_out[8][10][2] = xor_out[40][10][2] + xor_out[41][10][2] + xor_out[42][10][2] + xor_out[43][10][2] + xor_out[44][10][2];
assign sum_out[9][10][2] = xor_out[45][10][2] + xor_out[46][10][2] + xor_out[47][10][2] + xor_out[48][10][2] + xor_out[49][10][2];
assign sum_out[10][10][2] = xor_out[50][10][2] + xor_out[51][10][2] + xor_out[52][10][2] + xor_out[53][10][2] + xor_out[54][10][2];
assign sum_out[11][10][2] = xor_out[55][10][2] + xor_out[56][10][2] + xor_out[57][10][2] + xor_out[58][10][2] + xor_out[59][10][2];
assign sum_out[12][10][2] = xor_out[60][10][2] + xor_out[61][10][2] + xor_out[62][10][2] + xor_out[63][10][2] + xor_out[64][10][2];
assign sum_out[13][10][2] = xor_out[65][10][2] + xor_out[66][10][2] + xor_out[67][10][2] + xor_out[68][10][2] + xor_out[69][10][2];
assign sum_out[14][10][2] = xor_out[70][10][2] + xor_out[71][10][2] + xor_out[72][10][2] + xor_out[73][10][2] + xor_out[74][10][2];
assign sum_out[15][10][2] = xor_out[75][10][2] + xor_out[76][10][2] + xor_out[77][10][2] + xor_out[78][10][2] + xor_out[79][10][2];
assign sum_out[16][10][2] = xor_out[80][10][2] + xor_out[81][10][2] + xor_out[82][10][2] + xor_out[83][10][2] + xor_out[84][10][2];
assign sum_out[17][10][2] = xor_out[85][10][2] + xor_out[86][10][2] + xor_out[87][10][2] + xor_out[88][10][2] + xor_out[89][10][2];
assign sum_out[18][10][2] = xor_out[90][10][2] + xor_out[91][10][2] + xor_out[92][10][2] + xor_out[93][10][2] + xor_out[94][10][2];
assign sum_out[19][10][2] = xor_out[95][10][2] + xor_out[96][10][2] + xor_out[97][10][2] + xor_out[98][10][2] + xor_out[99][10][2];

assign sum_out[0][10][3] = xor_out[0][10][3] + xor_out[1][10][3] + xor_out[2][10][3] + xor_out[3][10][3] + xor_out[4][10][3];
assign sum_out[1][10][3] = xor_out[5][10][3] + xor_out[6][10][3] + xor_out[7][10][3] + xor_out[8][10][3] + xor_out[9][10][3];
assign sum_out[2][10][3] = xor_out[10][10][3] + xor_out[11][10][3] + xor_out[12][10][3] + xor_out[13][10][3] + xor_out[14][10][3];
assign sum_out[3][10][3] = xor_out[15][10][3] + xor_out[16][10][3] + xor_out[17][10][3] + xor_out[18][10][3] + xor_out[19][10][3];
assign sum_out[4][10][3] = xor_out[20][10][3] + xor_out[21][10][3] + xor_out[22][10][3] + xor_out[23][10][3] + xor_out[24][10][3];
assign sum_out[5][10][3] = xor_out[25][10][3] + xor_out[26][10][3] + xor_out[27][10][3] + xor_out[28][10][3] + xor_out[29][10][3];
assign sum_out[6][10][3] = xor_out[30][10][3] + xor_out[31][10][3] + xor_out[32][10][3] + xor_out[33][10][3] + xor_out[34][10][3];
assign sum_out[7][10][3] = xor_out[35][10][3] + xor_out[36][10][3] + xor_out[37][10][3] + xor_out[38][10][3] + xor_out[39][10][3];
assign sum_out[8][10][3] = xor_out[40][10][3] + xor_out[41][10][3] + xor_out[42][10][3] + xor_out[43][10][3] + xor_out[44][10][3];
assign sum_out[9][10][3] = xor_out[45][10][3] + xor_out[46][10][3] + xor_out[47][10][3] + xor_out[48][10][3] + xor_out[49][10][3];
assign sum_out[10][10][3] = xor_out[50][10][3] + xor_out[51][10][3] + xor_out[52][10][3] + xor_out[53][10][3] + xor_out[54][10][3];
assign sum_out[11][10][3] = xor_out[55][10][3] + xor_out[56][10][3] + xor_out[57][10][3] + xor_out[58][10][3] + xor_out[59][10][3];
assign sum_out[12][10][3] = xor_out[60][10][3] + xor_out[61][10][3] + xor_out[62][10][3] + xor_out[63][10][3] + xor_out[64][10][3];
assign sum_out[13][10][3] = xor_out[65][10][3] + xor_out[66][10][3] + xor_out[67][10][3] + xor_out[68][10][3] + xor_out[69][10][3];
assign sum_out[14][10][3] = xor_out[70][10][3] + xor_out[71][10][3] + xor_out[72][10][3] + xor_out[73][10][3] + xor_out[74][10][3];
assign sum_out[15][10][3] = xor_out[75][10][3] + xor_out[76][10][3] + xor_out[77][10][3] + xor_out[78][10][3] + xor_out[79][10][3];
assign sum_out[16][10][3] = xor_out[80][10][3] + xor_out[81][10][3] + xor_out[82][10][3] + xor_out[83][10][3] + xor_out[84][10][3];
assign sum_out[17][10][3] = xor_out[85][10][3] + xor_out[86][10][3] + xor_out[87][10][3] + xor_out[88][10][3] + xor_out[89][10][3];
assign sum_out[18][10][3] = xor_out[90][10][3] + xor_out[91][10][3] + xor_out[92][10][3] + xor_out[93][10][3] + xor_out[94][10][3];
assign sum_out[19][10][3] = xor_out[95][10][3] + xor_out[96][10][3] + xor_out[97][10][3] + xor_out[98][10][3] + xor_out[99][10][3];

assign sum_out[0][10][4] = xor_out[0][10][4] + xor_out[1][10][4] + xor_out[2][10][4] + xor_out[3][10][4] + xor_out[4][10][4];
assign sum_out[1][10][4] = xor_out[5][10][4] + xor_out[6][10][4] + xor_out[7][10][4] + xor_out[8][10][4] + xor_out[9][10][4];
assign sum_out[2][10][4] = xor_out[10][10][4] + xor_out[11][10][4] + xor_out[12][10][4] + xor_out[13][10][4] + xor_out[14][10][4];
assign sum_out[3][10][4] = xor_out[15][10][4] + xor_out[16][10][4] + xor_out[17][10][4] + xor_out[18][10][4] + xor_out[19][10][4];
assign sum_out[4][10][4] = xor_out[20][10][4] + xor_out[21][10][4] + xor_out[22][10][4] + xor_out[23][10][4] + xor_out[24][10][4];
assign sum_out[5][10][4] = xor_out[25][10][4] + xor_out[26][10][4] + xor_out[27][10][4] + xor_out[28][10][4] + xor_out[29][10][4];
assign sum_out[6][10][4] = xor_out[30][10][4] + xor_out[31][10][4] + xor_out[32][10][4] + xor_out[33][10][4] + xor_out[34][10][4];
assign sum_out[7][10][4] = xor_out[35][10][4] + xor_out[36][10][4] + xor_out[37][10][4] + xor_out[38][10][4] + xor_out[39][10][4];
assign sum_out[8][10][4] = xor_out[40][10][4] + xor_out[41][10][4] + xor_out[42][10][4] + xor_out[43][10][4] + xor_out[44][10][4];
assign sum_out[9][10][4] = xor_out[45][10][4] + xor_out[46][10][4] + xor_out[47][10][4] + xor_out[48][10][4] + xor_out[49][10][4];
assign sum_out[10][10][4] = xor_out[50][10][4] + xor_out[51][10][4] + xor_out[52][10][4] + xor_out[53][10][4] + xor_out[54][10][4];
assign sum_out[11][10][4] = xor_out[55][10][4] + xor_out[56][10][4] + xor_out[57][10][4] + xor_out[58][10][4] + xor_out[59][10][4];
assign sum_out[12][10][4] = xor_out[60][10][4] + xor_out[61][10][4] + xor_out[62][10][4] + xor_out[63][10][4] + xor_out[64][10][4];
assign sum_out[13][10][4] = xor_out[65][10][4] + xor_out[66][10][4] + xor_out[67][10][4] + xor_out[68][10][4] + xor_out[69][10][4];
assign sum_out[14][10][4] = xor_out[70][10][4] + xor_out[71][10][4] + xor_out[72][10][4] + xor_out[73][10][4] + xor_out[74][10][4];
assign sum_out[15][10][4] = xor_out[75][10][4] + xor_out[76][10][4] + xor_out[77][10][4] + xor_out[78][10][4] + xor_out[79][10][4];
assign sum_out[16][10][4] = xor_out[80][10][4] + xor_out[81][10][4] + xor_out[82][10][4] + xor_out[83][10][4] + xor_out[84][10][4];
assign sum_out[17][10][4] = xor_out[85][10][4] + xor_out[86][10][4] + xor_out[87][10][4] + xor_out[88][10][4] + xor_out[89][10][4];
assign sum_out[18][10][4] = xor_out[90][10][4] + xor_out[91][10][4] + xor_out[92][10][4] + xor_out[93][10][4] + xor_out[94][10][4];
assign sum_out[19][10][4] = xor_out[95][10][4] + xor_out[96][10][4] + xor_out[97][10][4] + xor_out[98][10][4] + xor_out[99][10][4];

assign sum_out[0][10][5] = xor_out[0][10][5] + xor_out[1][10][5] + xor_out[2][10][5] + xor_out[3][10][5] + xor_out[4][10][5];
assign sum_out[1][10][5] = xor_out[5][10][5] + xor_out[6][10][5] + xor_out[7][10][5] + xor_out[8][10][5] + xor_out[9][10][5];
assign sum_out[2][10][5] = xor_out[10][10][5] + xor_out[11][10][5] + xor_out[12][10][5] + xor_out[13][10][5] + xor_out[14][10][5];
assign sum_out[3][10][5] = xor_out[15][10][5] + xor_out[16][10][5] + xor_out[17][10][5] + xor_out[18][10][5] + xor_out[19][10][5];
assign sum_out[4][10][5] = xor_out[20][10][5] + xor_out[21][10][5] + xor_out[22][10][5] + xor_out[23][10][5] + xor_out[24][10][5];
assign sum_out[5][10][5] = xor_out[25][10][5] + xor_out[26][10][5] + xor_out[27][10][5] + xor_out[28][10][5] + xor_out[29][10][5];
assign sum_out[6][10][5] = xor_out[30][10][5] + xor_out[31][10][5] + xor_out[32][10][5] + xor_out[33][10][5] + xor_out[34][10][5];
assign sum_out[7][10][5] = xor_out[35][10][5] + xor_out[36][10][5] + xor_out[37][10][5] + xor_out[38][10][5] + xor_out[39][10][5];
assign sum_out[8][10][5] = xor_out[40][10][5] + xor_out[41][10][5] + xor_out[42][10][5] + xor_out[43][10][5] + xor_out[44][10][5];
assign sum_out[9][10][5] = xor_out[45][10][5] + xor_out[46][10][5] + xor_out[47][10][5] + xor_out[48][10][5] + xor_out[49][10][5];
assign sum_out[10][10][5] = xor_out[50][10][5] + xor_out[51][10][5] + xor_out[52][10][5] + xor_out[53][10][5] + xor_out[54][10][5];
assign sum_out[11][10][5] = xor_out[55][10][5] + xor_out[56][10][5] + xor_out[57][10][5] + xor_out[58][10][5] + xor_out[59][10][5];
assign sum_out[12][10][5] = xor_out[60][10][5] + xor_out[61][10][5] + xor_out[62][10][5] + xor_out[63][10][5] + xor_out[64][10][5];
assign sum_out[13][10][5] = xor_out[65][10][5] + xor_out[66][10][5] + xor_out[67][10][5] + xor_out[68][10][5] + xor_out[69][10][5];
assign sum_out[14][10][5] = xor_out[70][10][5] + xor_out[71][10][5] + xor_out[72][10][5] + xor_out[73][10][5] + xor_out[74][10][5];
assign sum_out[15][10][5] = xor_out[75][10][5] + xor_out[76][10][5] + xor_out[77][10][5] + xor_out[78][10][5] + xor_out[79][10][5];
assign sum_out[16][10][5] = xor_out[80][10][5] + xor_out[81][10][5] + xor_out[82][10][5] + xor_out[83][10][5] + xor_out[84][10][5];
assign sum_out[17][10][5] = xor_out[85][10][5] + xor_out[86][10][5] + xor_out[87][10][5] + xor_out[88][10][5] + xor_out[89][10][5];
assign sum_out[18][10][5] = xor_out[90][10][5] + xor_out[91][10][5] + xor_out[92][10][5] + xor_out[93][10][5] + xor_out[94][10][5];
assign sum_out[19][10][5] = xor_out[95][10][5] + xor_out[96][10][5] + xor_out[97][10][5] + xor_out[98][10][5] + xor_out[99][10][5];

assign sum_out[0][10][6] = xor_out[0][10][6] + xor_out[1][10][6] + xor_out[2][10][6] + xor_out[3][10][6] + xor_out[4][10][6];
assign sum_out[1][10][6] = xor_out[5][10][6] + xor_out[6][10][6] + xor_out[7][10][6] + xor_out[8][10][6] + xor_out[9][10][6];
assign sum_out[2][10][6] = xor_out[10][10][6] + xor_out[11][10][6] + xor_out[12][10][6] + xor_out[13][10][6] + xor_out[14][10][6];
assign sum_out[3][10][6] = xor_out[15][10][6] + xor_out[16][10][6] + xor_out[17][10][6] + xor_out[18][10][6] + xor_out[19][10][6];
assign sum_out[4][10][6] = xor_out[20][10][6] + xor_out[21][10][6] + xor_out[22][10][6] + xor_out[23][10][6] + xor_out[24][10][6];
assign sum_out[5][10][6] = xor_out[25][10][6] + xor_out[26][10][6] + xor_out[27][10][6] + xor_out[28][10][6] + xor_out[29][10][6];
assign sum_out[6][10][6] = xor_out[30][10][6] + xor_out[31][10][6] + xor_out[32][10][6] + xor_out[33][10][6] + xor_out[34][10][6];
assign sum_out[7][10][6] = xor_out[35][10][6] + xor_out[36][10][6] + xor_out[37][10][6] + xor_out[38][10][6] + xor_out[39][10][6];
assign sum_out[8][10][6] = xor_out[40][10][6] + xor_out[41][10][6] + xor_out[42][10][6] + xor_out[43][10][6] + xor_out[44][10][6];
assign sum_out[9][10][6] = xor_out[45][10][6] + xor_out[46][10][6] + xor_out[47][10][6] + xor_out[48][10][6] + xor_out[49][10][6];
assign sum_out[10][10][6] = xor_out[50][10][6] + xor_out[51][10][6] + xor_out[52][10][6] + xor_out[53][10][6] + xor_out[54][10][6];
assign sum_out[11][10][6] = xor_out[55][10][6] + xor_out[56][10][6] + xor_out[57][10][6] + xor_out[58][10][6] + xor_out[59][10][6];
assign sum_out[12][10][6] = xor_out[60][10][6] + xor_out[61][10][6] + xor_out[62][10][6] + xor_out[63][10][6] + xor_out[64][10][6];
assign sum_out[13][10][6] = xor_out[65][10][6] + xor_out[66][10][6] + xor_out[67][10][6] + xor_out[68][10][6] + xor_out[69][10][6];
assign sum_out[14][10][6] = xor_out[70][10][6] + xor_out[71][10][6] + xor_out[72][10][6] + xor_out[73][10][6] + xor_out[74][10][6];
assign sum_out[15][10][6] = xor_out[75][10][6] + xor_out[76][10][6] + xor_out[77][10][6] + xor_out[78][10][6] + xor_out[79][10][6];
assign sum_out[16][10][6] = xor_out[80][10][6] + xor_out[81][10][6] + xor_out[82][10][6] + xor_out[83][10][6] + xor_out[84][10][6];
assign sum_out[17][10][6] = xor_out[85][10][6] + xor_out[86][10][6] + xor_out[87][10][6] + xor_out[88][10][6] + xor_out[89][10][6];
assign sum_out[18][10][6] = xor_out[90][10][6] + xor_out[91][10][6] + xor_out[92][10][6] + xor_out[93][10][6] + xor_out[94][10][6];
assign sum_out[19][10][6] = xor_out[95][10][6] + xor_out[96][10][6] + xor_out[97][10][6] + xor_out[98][10][6] + xor_out[99][10][6];

assign sum_out[0][10][7] = xor_out[0][10][7] + xor_out[1][10][7] + xor_out[2][10][7] + xor_out[3][10][7] + xor_out[4][10][7];
assign sum_out[1][10][7] = xor_out[5][10][7] + xor_out[6][10][7] + xor_out[7][10][7] + xor_out[8][10][7] + xor_out[9][10][7];
assign sum_out[2][10][7] = xor_out[10][10][7] + xor_out[11][10][7] + xor_out[12][10][7] + xor_out[13][10][7] + xor_out[14][10][7];
assign sum_out[3][10][7] = xor_out[15][10][7] + xor_out[16][10][7] + xor_out[17][10][7] + xor_out[18][10][7] + xor_out[19][10][7];
assign sum_out[4][10][7] = xor_out[20][10][7] + xor_out[21][10][7] + xor_out[22][10][7] + xor_out[23][10][7] + xor_out[24][10][7];
assign sum_out[5][10][7] = xor_out[25][10][7] + xor_out[26][10][7] + xor_out[27][10][7] + xor_out[28][10][7] + xor_out[29][10][7];
assign sum_out[6][10][7] = xor_out[30][10][7] + xor_out[31][10][7] + xor_out[32][10][7] + xor_out[33][10][7] + xor_out[34][10][7];
assign sum_out[7][10][7] = xor_out[35][10][7] + xor_out[36][10][7] + xor_out[37][10][7] + xor_out[38][10][7] + xor_out[39][10][7];
assign sum_out[8][10][7] = xor_out[40][10][7] + xor_out[41][10][7] + xor_out[42][10][7] + xor_out[43][10][7] + xor_out[44][10][7];
assign sum_out[9][10][7] = xor_out[45][10][7] + xor_out[46][10][7] + xor_out[47][10][7] + xor_out[48][10][7] + xor_out[49][10][7];
assign sum_out[10][10][7] = xor_out[50][10][7] + xor_out[51][10][7] + xor_out[52][10][7] + xor_out[53][10][7] + xor_out[54][10][7];
assign sum_out[11][10][7] = xor_out[55][10][7] + xor_out[56][10][7] + xor_out[57][10][7] + xor_out[58][10][7] + xor_out[59][10][7];
assign sum_out[12][10][7] = xor_out[60][10][7] + xor_out[61][10][7] + xor_out[62][10][7] + xor_out[63][10][7] + xor_out[64][10][7];
assign sum_out[13][10][7] = xor_out[65][10][7] + xor_out[66][10][7] + xor_out[67][10][7] + xor_out[68][10][7] + xor_out[69][10][7];
assign sum_out[14][10][7] = xor_out[70][10][7] + xor_out[71][10][7] + xor_out[72][10][7] + xor_out[73][10][7] + xor_out[74][10][7];
assign sum_out[15][10][7] = xor_out[75][10][7] + xor_out[76][10][7] + xor_out[77][10][7] + xor_out[78][10][7] + xor_out[79][10][7];
assign sum_out[16][10][7] = xor_out[80][10][7] + xor_out[81][10][7] + xor_out[82][10][7] + xor_out[83][10][7] + xor_out[84][10][7];
assign sum_out[17][10][7] = xor_out[85][10][7] + xor_out[86][10][7] + xor_out[87][10][7] + xor_out[88][10][7] + xor_out[89][10][7];
assign sum_out[18][10][7] = xor_out[90][10][7] + xor_out[91][10][7] + xor_out[92][10][7] + xor_out[93][10][7] + xor_out[94][10][7];
assign sum_out[19][10][7] = xor_out[95][10][7] + xor_out[96][10][7] + xor_out[97][10][7] + xor_out[98][10][7] + xor_out[99][10][7];

assign sum_out[0][10][8] = xor_out[0][10][8] + xor_out[1][10][8] + xor_out[2][10][8] + xor_out[3][10][8] + xor_out[4][10][8];
assign sum_out[1][10][8] = xor_out[5][10][8] + xor_out[6][10][8] + xor_out[7][10][8] + xor_out[8][10][8] + xor_out[9][10][8];
assign sum_out[2][10][8] = xor_out[10][10][8] + xor_out[11][10][8] + xor_out[12][10][8] + xor_out[13][10][8] + xor_out[14][10][8];
assign sum_out[3][10][8] = xor_out[15][10][8] + xor_out[16][10][8] + xor_out[17][10][8] + xor_out[18][10][8] + xor_out[19][10][8];
assign sum_out[4][10][8] = xor_out[20][10][8] + xor_out[21][10][8] + xor_out[22][10][8] + xor_out[23][10][8] + xor_out[24][10][8];
assign sum_out[5][10][8] = xor_out[25][10][8] + xor_out[26][10][8] + xor_out[27][10][8] + xor_out[28][10][8] + xor_out[29][10][8];
assign sum_out[6][10][8] = xor_out[30][10][8] + xor_out[31][10][8] + xor_out[32][10][8] + xor_out[33][10][8] + xor_out[34][10][8];
assign sum_out[7][10][8] = xor_out[35][10][8] + xor_out[36][10][8] + xor_out[37][10][8] + xor_out[38][10][8] + xor_out[39][10][8];
assign sum_out[8][10][8] = xor_out[40][10][8] + xor_out[41][10][8] + xor_out[42][10][8] + xor_out[43][10][8] + xor_out[44][10][8];
assign sum_out[9][10][8] = xor_out[45][10][8] + xor_out[46][10][8] + xor_out[47][10][8] + xor_out[48][10][8] + xor_out[49][10][8];
assign sum_out[10][10][8] = xor_out[50][10][8] + xor_out[51][10][8] + xor_out[52][10][8] + xor_out[53][10][8] + xor_out[54][10][8];
assign sum_out[11][10][8] = xor_out[55][10][8] + xor_out[56][10][8] + xor_out[57][10][8] + xor_out[58][10][8] + xor_out[59][10][8];
assign sum_out[12][10][8] = xor_out[60][10][8] + xor_out[61][10][8] + xor_out[62][10][8] + xor_out[63][10][8] + xor_out[64][10][8];
assign sum_out[13][10][8] = xor_out[65][10][8] + xor_out[66][10][8] + xor_out[67][10][8] + xor_out[68][10][8] + xor_out[69][10][8];
assign sum_out[14][10][8] = xor_out[70][10][8] + xor_out[71][10][8] + xor_out[72][10][8] + xor_out[73][10][8] + xor_out[74][10][8];
assign sum_out[15][10][8] = xor_out[75][10][8] + xor_out[76][10][8] + xor_out[77][10][8] + xor_out[78][10][8] + xor_out[79][10][8];
assign sum_out[16][10][8] = xor_out[80][10][8] + xor_out[81][10][8] + xor_out[82][10][8] + xor_out[83][10][8] + xor_out[84][10][8];
assign sum_out[17][10][8] = xor_out[85][10][8] + xor_out[86][10][8] + xor_out[87][10][8] + xor_out[88][10][8] + xor_out[89][10][8];
assign sum_out[18][10][8] = xor_out[90][10][8] + xor_out[91][10][8] + xor_out[92][10][8] + xor_out[93][10][8] + xor_out[94][10][8];
assign sum_out[19][10][8] = xor_out[95][10][8] + xor_out[96][10][8] + xor_out[97][10][8] + xor_out[98][10][8] + xor_out[99][10][8];

assign sum_out[0][10][9] = xor_out[0][10][9] + xor_out[1][10][9] + xor_out[2][10][9] + xor_out[3][10][9] + xor_out[4][10][9];
assign sum_out[1][10][9] = xor_out[5][10][9] + xor_out[6][10][9] + xor_out[7][10][9] + xor_out[8][10][9] + xor_out[9][10][9];
assign sum_out[2][10][9] = xor_out[10][10][9] + xor_out[11][10][9] + xor_out[12][10][9] + xor_out[13][10][9] + xor_out[14][10][9];
assign sum_out[3][10][9] = xor_out[15][10][9] + xor_out[16][10][9] + xor_out[17][10][9] + xor_out[18][10][9] + xor_out[19][10][9];
assign sum_out[4][10][9] = xor_out[20][10][9] + xor_out[21][10][9] + xor_out[22][10][9] + xor_out[23][10][9] + xor_out[24][10][9];
assign sum_out[5][10][9] = xor_out[25][10][9] + xor_out[26][10][9] + xor_out[27][10][9] + xor_out[28][10][9] + xor_out[29][10][9];
assign sum_out[6][10][9] = xor_out[30][10][9] + xor_out[31][10][9] + xor_out[32][10][9] + xor_out[33][10][9] + xor_out[34][10][9];
assign sum_out[7][10][9] = xor_out[35][10][9] + xor_out[36][10][9] + xor_out[37][10][9] + xor_out[38][10][9] + xor_out[39][10][9];
assign sum_out[8][10][9] = xor_out[40][10][9] + xor_out[41][10][9] + xor_out[42][10][9] + xor_out[43][10][9] + xor_out[44][10][9];
assign sum_out[9][10][9] = xor_out[45][10][9] + xor_out[46][10][9] + xor_out[47][10][9] + xor_out[48][10][9] + xor_out[49][10][9];
assign sum_out[10][10][9] = xor_out[50][10][9] + xor_out[51][10][9] + xor_out[52][10][9] + xor_out[53][10][9] + xor_out[54][10][9];
assign sum_out[11][10][9] = xor_out[55][10][9] + xor_out[56][10][9] + xor_out[57][10][9] + xor_out[58][10][9] + xor_out[59][10][9];
assign sum_out[12][10][9] = xor_out[60][10][9] + xor_out[61][10][9] + xor_out[62][10][9] + xor_out[63][10][9] + xor_out[64][10][9];
assign sum_out[13][10][9] = xor_out[65][10][9] + xor_out[66][10][9] + xor_out[67][10][9] + xor_out[68][10][9] + xor_out[69][10][9];
assign sum_out[14][10][9] = xor_out[70][10][9] + xor_out[71][10][9] + xor_out[72][10][9] + xor_out[73][10][9] + xor_out[74][10][9];
assign sum_out[15][10][9] = xor_out[75][10][9] + xor_out[76][10][9] + xor_out[77][10][9] + xor_out[78][10][9] + xor_out[79][10][9];
assign sum_out[16][10][9] = xor_out[80][10][9] + xor_out[81][10][9] + xor_out[82][10][9] + xor_out[83][10][9] + xor_out[84][10][9];
assign sum_out[17][10][9] = xor_out[85][10][9] + xor_out[86][10][9] + xor_out[87][10][9] + xor_out[88][10][9] + xor_out[89][10][9];
assign sum_out[18][10][9] = xor_out[90][10][9] + xor_out[91][10][9] + xor_out[92][10][9] + xor_out[93][10][9] + xor_out[94][10][9];
assign sum_out[19][10][9] = xor_out[95][10][9] + xor_out[96][10][9] + xor_out[97][10][9] + xor_out[98][10][9] + xor_out[99][10][9];

assign sum_out[0][10][10] = xor_out[0][10][10] + xor_out[1][10][10] + xor_out[2][10][10] + xor_out[3][10][10] + xor_out[4][10][10];
assign sum_out[1][10][10] = xor_out[5][10][10] + xor_out[6][10][10] + xor_out[7][10][10] + xor_out[8][10][10] + xor_out[9][10][10];
assign sum_out[2][10][10] = xor_out[10][10][10] + xor_out[11][10][10] + xor_out[12][10][10] + xor_out[13][10][10] + xor_out[14][10][10];
assign sum_out[3][10][10] = xor_out[15][10][10] + xor_out[16][10][10] + xor_out[17][10][10] + xor_out[18][10][10] + xor_out[19][10][10];
assign sum_out[4][10][10] = xor_out[20][10][10] + xor_out[21][10][10] + xor_out[22][10][10] + xor_out[23][10][10] + xor_out[24][10][10];
assign sum_out[5][10][10] = xor_out[25][10][10] + xor_out[26][10][10] + xor_out[27][10][10] + xor_out[28][10][10] + xor_out[29][10][10];
assign sum_out[6][10][10] = xor_out[30][10][10] + xor_out[31][10][10] + xor_out[32][10][10] + xor_out[33][10][10] + xor_out[34][10][10];
assign sum_out[7][10][10] = xor_out[35][10][10] + xor_out[36][10][10] + xor_out[37][10][10] + xor_out[38][10][10] + xor_out[39][10][10];
assign sum_out[8][10][10] = xor_out[40][10][10] + xor_out[41][10][10] + xor_out[42][10][10] + xor_out[43][10][10] + xor_out[44][10][10];
assign sum_out[9][10][10] = xor_out[45][10][10] + xor_out[46][10][10] + xor_out[47][10][10] + xor_out[48][10][10] + xor_out[49][10][10];
assign sum_out[10][10][10] = xor_out[50][10][10] + xor_out[51][10][10] + xor_out[52][10][10] + xor_out[53][10][10] + xor_out[54][10][10];
assign sum_out[11][10][10] = xor_out[55][10][10] + xor_out[56][10][10] + xor_out[57][10][10] + xor_out[58][10][10] + xor_out[59][10][10];
assign sum_out[12][10][10] = xor_out[60][10][10] + xor_out[61][10][10] + xor_out[62][10][10] + xor_out[63][10][10] + xor_out[64][10][10];
assign sum_out[13][10][10] = xor_out[65][10][10] + xor_out[66][10][10] + xor_out[67][10][10] + xor_out[68][10][10] + xor_out[69][10][10];
assign sum_out[14][10][10] = xor_out[70][10][10] + xor_out[71][10][10] + xor_out[72][10][10] + xor_out[73][10][10] + xor_out[74][10][10];
assign sum_out[15][10][10] = xor_out[75][10][10] + xor_out[76][10][10] + xor_out[77][10][10] + xor_out[78][10][10] + xor_out[79][10][10];
assign sum_out[16][10][10] = xor_out[80][10][10] + xor_out[81][10][10] + xor_out[82][10][10] + xor_out[83][10][10] + xor_out[84][10][10];
assign sum_out[17][10][10] = xor_out[85][10][10] + xor_out[86][10][10] + xor_out[87][10][10] + xor_out[88][10][10] + xor_out[89][10][10];
assign sum_out[18][10][10] = xor_out[90][10][10] + xor_out[91][10][10] + xor_out[92][10][10] + xor_out[93][10][10] + xor_out[94][10][10];
assign sum_out[19][10][10] = xor_out[95][10][10] + xor_out[96][10][10] + xor_out[97][10][10] + xor_out[98][10][10] + xor_out[99][10][10];

assign sum_out[0][10][11] = xor_out[0][10][11] + xor_out[1][10][11] + xor_out[2][10][11] + xor_out[3][10][11] + xor_out[4][10][11];
assign sum_out[1][10][11] = xor_out[5][10][11] + xor_out[6][10][11] + xor_out[7][10][11] + xor_out[8][10][11] + xor_out[9][10][11];
assign sum_out[2][10][11] = xor_out[10][10][11] + xor_out[11][10][11] + xor_out[12][10][11] + xor_out[13][10][11] + xor_out[14][10][11];
assign sum_out[3][10][11] = xor_out[15][10][11] + xor_out[16][10][11] + xor_out[17][10][11] + xor_out[18][10][11] + xor_out[19][10][11];
assign sum_out[4][10][11] = xor_out[20][10][11] + xor_out[21][10][11] + xor_out[22][10][11] + xor_out[23][10][11] + xor_out[24][10][11];
assign sum_out[5][10][11] = xor_out[25][10][11] + xor_out[26][10][11] + xor_out[27][10][11] + xor_out[28][10][11] + xor_out[29][10][11];
assign sum_out[6][10][11] = xor_out[30][10][11] + xor_out[31][10][11] + xor_out[32][10][11] + xor_out[33][10][11] + xor_out[34][10][11];
assign sum_out[7][10][11] = xor_out[35][10][11] + xor_out[36][10][11] + xor_out[37][10][11] + xor_out[38][10][11] + xor_out[39][10][11];
assign sum_out[8][10][11] = xor_out[40][10][11] + xor_out[41][10][11] + xor_out[42][10][11] + xor_out[43][10][11] + xor_out[44][10][11];
assign sum_out[9][10][11] = xor_out[45][10][11] + xor_out[46][10][11] + xor_out[47][10][11] + xor_out[48][10][11] + xor_out[49][10][11];
assign sum_out[10][10][11] = xor_out[50][10][11] + xor_out[51][10][11] + xor_out[52][10][11] + xor_out[53][10][11] + xor_out[54][10][11];
assign sum_out[11][10][11] = xor_out[55][10][11] + xor_out[56][10][11] + xor_out[57][10][11] + xor_out[58][10][11] + xor_out[59][10][11];
assign sum_out[12][10][11] = xor_out[60][10][11] + xor_out[61][10][11] + xor_out[62][10][11] + xor_out[63][10][11] + xor_out[64][10][11];
assign sum_out[13][10][11] = xor_out[65][10][11] + xor_out[66][10][11] + xor_out[67][10][11] + xor_out[68][10][11] + xor_out[69][10][11];
assign sum_out[14][10][11] = xor_out[70][10][11] + xor_out[71][10][11] + xor_out[72][10][11] + xor_out[73][10][11] + xor_out[74][10][11];
assign sum_out[15][10][11] = xor_out[75][10][11] + xor_out[76][10][11] + xor_out[77][10][11] + xor_out[78][10][11] + xor_out[79][10][11];
assign sum_out[16][10][11] = xor_out[80][10][11] + xor_out[81][10][11] + xor_out[82][10][11] + xor_out[83][10][11] + xor_out[84][10][11];
assign sum_out[17][10][11] = xor_out[85][10][11] + xor_out[86][10][11] + xor_out[87][10][11] + xor_out[88][10][11] + xor_out[89][10][11];
assign sum_out[18][10][11] = xor_out[90][10][11] + xor_out[91][10][11] + xor_out[92][10][11] + xor_out[93][10][11] + xor_out[94][10][11];
assign sum_out[19][10][11] = xor_out[95][10][11] + xor_out[96][10][11] + xor_out[97][10][11] + xor_out[98][10][11] + xor_out[99][10][11];

assign sum_out[0][10][12] = xor_out[0][10][12] + xor_out[1][10][12] + xor_out[2][10][12] + xor_out[3][10][12] + xor_out[4][10][12];
assign sum_out[1][10][12] = xor_out[5][10][12] + xor_out[6][10][12] + xor_out[7][10][12] + xor_out[8][10][12] + xor_out[9][10][12];
assign sum_out[2][10][12] = xor_out[10][10][12] + xor_out[11][10][12] + xor_out[12][10][12] + xor_out[13][10][12] + xor_out[14][10][12];
assign sum_out[3][10][12] = xor_out[15][10][12] + xor_out[16][10][12] + xor_out[17][10][12] + xor_out[18][10][12] + xor_out[19][10][12];
assign sum_out[4][10][12] = xor_out[20][10][12] + xor_out[21][10][12] + xor_out[22][10][12] + xor_out[23][10][12] + xor_out[24][10][12];
assign sum_out[5][10][12] = xor_out[25][10][12] + xor_out[26][10][12] + xor_out[27][10][12] + xor_out[28][10][12] + xor_out[29][10][12];
assign sum_out[6][10][12] = xor_out[30][10][12] + xor_out[31][10][12] + xor_out[32][10][12] + xor_out[33][10][12] + xor_out[34][10][12];
assign sum_out[7][10][12] = xor_out[35][10][12] + xor_out[36][10][12] + xor_out[37][10][12] + xor_out[38][10][12] + xor_out[39][10][12];
assign sum_out[8][10][12] = xor_out[40][10][12] + xor_out[41][10][12] + xor_out[42][10][12] + xor_out[43][10][12] + xor_out[44][10][12];
assign sum_out[9][10][12] = xor_out[45][10][12] + xor_out[46][10][12] + xor_out[47][10][12] + xor_out[48][10][12] + xor_out[49][10][12];
assign sum_out[10][10][12] = xor_out[50][10][12] + xor_out[51][10][12] + xor_out[52][10][12] + xor_out[53][10][12] + xor_out[54][10][12];
assign sum_out[11][10][12] = xor_out[55][10][12] + xor_out[56][10][12] + xor_out[57][10][12] + xor_out[58][10][12] + xor_out[59][10][12];
assign sum_out[12][10][12] = xor_out[60][10][12] + xor_out[61][10][12] + xor_out[62][10][12] + xor_out[63][10][12] + xor_out[64][10][12];
assign sum_out[13][10][12] = xor_out[65][10][12] + xor_out[66][10][12] + xor_out[67][10][12] + xor_out[68][10][12] + xor_out[69][10][12];
assign sum_out[14][10][12] = xor_out[70][10][12] + xor_out[71][10][12] + xor_out[72][10][12] + xor_out[73][10][12] + xor_out[74][10][12];
assign sum_out[15][10][12] = xor_out[75][10][12] + xor_out[76][10][12] + xor_out[77][10][12] + xor_out[78][10][12] + xor_out[79][10][12];
assign sum_out[16][10][12] = xor_out[80][10][12] + xor_out[81][10][12] + xor_out[82][10][12] + xor_out[83][10][12] + xor_out[84][10][12];
assign sum_out[17][10][12] = xor_out[85][10][12] + xor_out[86][10][12] + xor_out[87][10][12] + xor_out[88][10][12] + xor_out[89][10][12];
assign sum_out[18][10][12] = xor_out[90][10][12] + xor_out[91][10][12] + xor_out[92][10][12] + xor_out[93][10][12] + xor_out[94][10][12];
assign sum_out[19][10][12] = xor_out[95][10][12] + xor_out[96][10][12] + xor_out[97][10][12] + xor_out[98][10][12] + xor_out[99][10][12];

assign sum_out[0][10][13] = xor_out[0][10][13] + xor_out[1][10][13] + xor_out[2][10][13] + xor_out[3][10][13] + xor_out[4][10][13];
assign sum_out[1][10][13] = xor_out[5][10][13] + xor_out[6][10][13] + xor_out[7][10][13] + xor_out[8][10][13] + xor_out[9][10][13];
assign sum_out[2][10][13] = xor_out[10][10][13] + xor_out[11][10][13] + xor_out[12][10][13] + xor_out[13][10][13] + xor_out[14][10][13];
assign sum_out[3][10][13] = xor_out[15][10][13] + xor_out[16][10][13] + xor_out[17][10][13] + xor_out[18][10][13] + xor_out[19][10][13];
assign sum_out[4][10][13] = xor_out[20][10][13] + xor_out[21][10][13] + xor_out[22][10][13] + xor_out[23][10][13] + xor_out[24][10][13];
assign sum_out[5][10][13] = xor_out[25][10][13] + xor_out[26][10][13] + xor_out[27][10][13] + xor_out[28][10][13] + xor_out[29][10][13];
assign sum_out[6][10][13] = xor_out[30][10][13] + xor_out[31][10][13] + xor_out[32][10][13] + xor_out[33][10][13] + xor_out[34][10][13];
assign sum_out[7][10][13] = xor_out[35][10][13] + xor_out[36][10][13] + xor_out[37][10][13] + xor_out[38][10][13] + xor_out[39][10][13];
assign sum_out[8][10][13] = xor_out[40][10][13] + xor_out[41][10][13] + xor_out[42][10][13] + xor_out[43][10][13] + xor_out[44][10][13];
assign sum_out[9][10][13] = xor_out[45][10][13] + xor_out[46][10][13] + xor_out[47][10][13] + xor_out[48][10][13] + xor_out[49][10][13];
assign sum_out[10][10][13] = xor_out[50][10][13] + xor_out[51][10][13] + xor_out[52][10][13] + xor_out[53][10][13] + xor_out[54][10][13];
assign sum_out[11][10][13] = xor_out[55][10][13] + xor_out[56][10][13] + xor_out[57][10][13] + xor_out[58][10][13] + xor_out[59][10][13];
assign sum_out[12][10][13] = xor_out[60][10][13] + xor_out[61][10][13] + xor_out[62][10][13] + xor_out[63][10][13] + xor_out[64][10][13];
assign sum_out[13][10][13] = xor_out[65][10][13] + xor_out[66][10][13] + xor_out[67][10][13] + xor_out[68][10][13] + xor_out[69][10][13];
assign sum_out[14][10][13] = xor_out[70][10][13] + xor_out[71][10][13] + xor_out[72][10][13] + xor_out[73][10][13] + xor_out[74][10][13];
assign sum_out[15][10][13] = xor_out[75][10][13] + xor_out[76][10][13] + xor_out[77][10][13] + xor_out[78][10][13] + xor_out[79][10][13];
assign sum_out[16][10][13] = xor_out[80][10][13] + xor_out[81][10][13] + xor_out[82][10][13] + xor_out[83][10][13] + xor_out[84][10][13];
assign sum_out[17][10][13] = xor_out[85][10][13] + xor_out[86][10][13] + xor_out[87][10][13] + xor_out[88][10][13] + xor_out[89][10][13];
assign sum_out[18][10][13] = xor_out[90][10][13] + xor_out[91][10][13] + xor_out[92][10][13] + xor_out[93][10][13] + xor_out[94][10][13];
assign sum_out[19][10][13] = xor_out[95][10][13] + xor_out[96][10][13] + xor_out[97][10][13] + xor_out[98][10][13] + xor_out[99][10][13];

assign sum_out[0][10][14] = xor_out[0][10][14] + xor_out[1][10][14] + xor_out[2][10][14] + xor_out[3][10][14] + xor_out[4][10][14];
assign sum_out[1][10][14] = xor_out[5][10][14] + xor_out[6][10][14] + xor_out[7][10][14] + xor_out[8][10][14] + xor_out[9][10][14];
assign sum_out[2][10][14] = xor_out[10][10][14] + xor_out[11][10][14] + xor_out[12][10][14] + xor_out[13][10][14] + xor_out[14][10][14];
assign sum_out[3][10][14] = xor_out[15][10][14] + xor_out[16][10][14] + xor_out[17][10][14] + xor_out[18][10][14] + xor_out[19][10][14];
assign sum_out[4][10][14] = xor_out[20][10][14] + xor_out[21][10][14] + xor_out[22][10][14] + xor_out[23][10][14] + xor_out[24][10][14];
assign sum_out[5][10][14] = xor_out[25][10][14] + xor_out[26][10][14] + xor_out[27][10][14] + xor_out[28][10][14] + xor_out[29][10][14];
assign sum_out[6][10][14] = xor_out[30][10][14] + xor_out[31][10][14] + xor_out[32][10][14] + xor_out[33][10][14] + xor_out[34][10][14];
assign sum_out[7][10][14] = xor_out[35][10][14] + xor_out[36][10][14] + xor_out[37][10][14] + xor_out[38][10][14] + xor_out[39][10][14];
assign sum_out[8][10][14] = xor_out[40][10][14] + xor_out[41][10][14] + xor_out[42][10][14] + xor_out[43][10][14] + xor_out[44][10][14];
assign sum_out[9][10][14] = xor_out[45][10][14] + xor_out[46][10][14] + xor_out[47][10][14] + xor_out[48][10][14] + xor_out[49][10][14];
assign sum_out[10][10][14] = xor_out[50][10][14] + xor_out[51][10][14] + xor_out[52][10][14] + xor_out[53][10][14] + xor_out[54][10][14];
assign sum_out[11][10][14] = xor_out[55][10][14] + xor_out[56][10][14] + xor_out[57][10][14] + xor_out[58][10][14] + xor_out[59][10][14];
assign sum_out[12][10][14] = xor_out[60][10][14] + xor_out[61][10][14] + xor_out[62][10][14] + xor_out[63][10][14] + xor_out[64][10][14];
assign sum_out[13][10][14] = xor_out[65][10][14] + xor_out[66][10][14] + xor_out[67][10][14] + xor_out[68][10][14] + xor_out[69][10][14];
assign sum_out[14][10][14] = xor_out[70][10][14] + xor_out[71][10][14] + xor_out[72][10][14] + xor_out[73][10][14] + xor_out[74][10][14];
assign sum_out[15][10][14] = xor_out[75][10][14] + xor_out[76][10][14] + xor_out[77][10][14] + xor_out[78][10][14] + xor_out[79][10][14];
assign sum_out[16][10][14] = xor_out[80][10][14] + xor_out[81][10][14] + xor_out[82][10][14] + xor_out[83][10][14] + xor_out[84][10][14];
assign sum_out[17][10][14] = xor_out[85][10][14] + xor_out[86][10][14] + xor_out[87][10][14] + xor_out[88][10][14] + xor_out[89][10][14];
assign sum_out[18][10][14] = xor_out[90][10][14] + xor_out[91][10][14] + xor_out[92][10][14] + xor_out[93][10][14] + xor_out[94][10][14];
assign sum_out[19][10][14] = xor_out[95][10][14] + xor_out[96][10][14] + xor_out[97][10][14] + xor_out[98][10][14] + xor_out[99][10][14];

assign sum_out[0][10][15] = xor_out[0][10][15] + xor_out[1][10][15] + xor_out[2][10][15] + xor_out[3][10][15] + xor_out[4][10][15];
assign sum_out[1][10][15] = xor_out[5][10][15] + xor_out[6][10][15] + xor_out[7][10][15] + xor_out[8][10][15] + xor_out[9][10][15];
assign sum_out[2][10][15] = xor_out[10][10][15] + xor_out[11][10][15] + xor_out[12][10][15] + xor_out[13][10][15] + xor_out[14][10][15];
assign sum_out[3][10][15] = xor_out[15][10][15] + xor_out[16][10][15] + xor_out[17][10][15] + xor_out[18][10][15] + xor_out[19][10][15];
assign sum_out[4][10][15] = xor_out[20][10][15] + xor_out[21][10][15] + xor_out[22][10][15] + xor_out[23][10][15] + xor_out[24][10][15];
assign sum_out[5][10][15] = xor_out[25][10][15] + xor_out[26][10][15] + xor_out[27][10][15] + xor_out[28][10][15] + xor_out[29][10][15];
assign sum_out[6][10][15] = xor_out[30][10][15] + xor_out[31][10][15] + xor_out[32][10][15] + xor_out[33][10][15] + xor_out[34][10][15];
assign sum_out[7][10][15] = xor_out[35][10][15] + xor_out[36][10][15] + xor_out[37][10][15] + xor_out[38][10][15] + xor_out[39][10][15];
assign sum_out[8][10][15] = xor_out[40][10][15] + xor_out[41][10][15] + xor_out[42][10][15] + xor_out[43][10][15] + xor_out[44][10][15];
assign sum_out[9][10][15] = xor_out[45][10][15] + xor_out[46][10][15] + xor_out[47][10][15] + xor_out[48][10][15] + xor_out[49][10][15];
assign sum_out[10][10][15] = xor_out[50][10][15] + xor_out[51][10][15] + xor_out[52][10][15] + xor_out[53][10][15] + xor_out[54][10][15];
assign sum_out[11][10][15] = xor_out[55][10][15] + xor_out[56][10][15] + xor_out[57][10][15] + xor_out[58][10][15] + xor_out[59][10][15];
assign sum_out[12][10][15] = xor_out[60][10][15] + xor_out[61][10][15] + xor_out[62][10][15] + xor_out[63][10][15] + xor_out[64][10][15];
assign sum_out[13][10][15] = xor_out[65][10][15] + xor_out[66][10][15] + xor_out[67][10][15] + xor_out[68][10][15] + xor_out[69][10][15];
assign sum_out[14][10][15] = xor_out[70][10][15] + xor_out[71][10][15] + xor_out[72][10][15] + xor_out[73][10][15] + xor_out[74][10][15];
assign sum_out[15][10][15] = xor_out[75][10][15] + xor_out[76][10][15] + xor_out[77][10][15] + xor_out[78][10][15] + xor_out[79][10][15];
assign sum_out[16][10][15] = xor_out[80][10][15] + xor_out[81][10][15] + xor_out[82][10][15] + xor_out[83][10][15] + xor_out[84][10][15];
assign sum_out[17][10][15] = xor_out[85][10][15] + xor_out[86][10][15] + xor_out[87][10][15] + xor_out[88][10][15] + xor_out[89][10][15];
assign sum_out[18][10][15] = xor_out[90][10][15] + xor_out[91][10][15] + xor_out[92][10][15] + xor_out[93][10][15] + xor_out[94][10][15];
assign sum_out[19][10][15] = xor_out[95][10][15] + xor_out[96][10][15] + xor_out[97][10][15] + xor_out[98][10][15] + xor_out[99][10][15];

assign sum_out[0][10][16] = xor_out[0][10][16] + xor_out[1][10][16] + xor_out[2][10][16] + xor_out[3][10][16] + xor_out[4][10][16];
assign sum_out[1][10][16] = xor_out[5][10][16] + xor_out[6][10][16] + xor_out[7][10][16] + xor_out[8][10][16] + xor_out[9][10][16];
assign sum_out[2][10][16] = xor_out[10][10][16] + xor_out[11][10][16] + xor_out[12][10][16] + xor_out[13][10][16] + xor_out[14][10][16];
assign sum_out[3][10][16] = xor_out[15][10][16] + xor_out[16][10][16] + xor_out[17][10][16] + xor_out[18][10][16] + xor_out[19][10][16];
assign sum_out[4][10][16] = xor_out[20][10][16] + xor_out[21][10][16] + xor_out[22][10][16] + xor_out[23][10][16] + xor_out[24][10][16];
assign sum_out[5][10][16] = xor_out[25][10][16] + xor_out[26][10][16] + xor_out[27][10][16] + xor_out[28][10][16] + xor_out[29][10][16];
assign sum_out[6][10][16] = xor_out[30][10][16] + xor_out[31][10][16] + xor_out[32][10][16] + xor_out[33][10][16] + xor_out[34][10][16];
assign sum_out[7][10][16] = xor_out[35][10][16] + xor_out[36][10][16] + xor_out[37][10][16] + xor_out[38][10][16] + xor_out[39][10][16];
assign sum_out[8][10][16] = xor_out[40][10][16] + xor_out[41][10][16] + xor_out[42][10][16] + xor_out[43][10][16] + xor_out[44][10][16];
assign sum_out[9][10][16] = xor_out[45][10][16] + xor_out[46][10][16] + xor_out[47][10][16] + xor_out[48][10][16] + xor_out[49][10][16];
assign sum_out[10][10][16] = xor_out[50][10][16] + xor_out[51][10][16] + xor_out[52][10][16] + xor_out[53][10][16] + xor_out[54][10][16];
assign sum_out[11][10][16] = xor_out[55][10][16] + xor_out[56][10][16] + xor_out[57][10][16] + xor_out[58][10][16] + xor_out[59][10][16];
assign sum_out[12][10][16] = xor_out[60][10][16] + xor_out[61][10][16] + xor_out[62][10][16] + xor_out[63][10][16] + xor_out[64][10][16];
assign sum_out[13][10][16] = xor_out[65][10][16] + xor_out[66][10][16] + xor_out[67][10][16] + xor_out[68][10][16] + xor_out[69][10][16];
assign sum_out[14][10][16] = xor_out[70][10][16] + xor_out[71][10][16] + xor_out[72][10][16] + xor_out[73][10][16] + xor_out[74][10][16];
assign sum_out[15][10][16] = xor_out[75][10][16] + xor_out[76][10][16] + xor_out[77][10][16] + xor_out[78][10][16] + xor_out[79][10][16];
assign sum_out[16][10][16] = xor_out[80][10][16] + xor_out[81][10][16] + xor_out[82][10][16] + xor_out[83][10][16] + xor_out[84][10][16];
assign sum_out[17][10][16] = xor_out[85][10][16] + xor_out[86][10][16] + xor_out[87][10][16] + xor_out[88][10][16] + xor_out[89][10][16];
assign sum_out[18][10][16] = xor_out[90][10][16] + xor_out[91][10][16] + xor_out[92][10][16] + xor_out[93][10][16] + xor_out[94][10][16];
assign sum_out[19][10][16] = xor_out[95][10][16] + xor_out[96][10][16] + xor_out[97][10][16] + xor_out[98][10][16] + xor_out[99][10][16];

assign sum_out[0][10][17] = xor_out[0][10][17] + xor_out[1][10][17] + xor_out[2][10][17] + xor_out[3][10][17] + xor_out[4][10][17];
assign sum_out[1][10][17] = xor_out[5][10][17] + xor_out[6][10][17] + xor_out[7][10][17] + xor_out[8][10][17] + xor_out[9][10][17];
assign sum_out[2][10][17] = xor_out[10][10][17] + xor_out[11][10][17] + xor_out[12][10][17] + xor_out[13][10][17] + xor_out[14][10][17];
assign sum_out[3][10][17] = xor_out[15][10][17] + xor_out[16][10][17] + xor_out[17][10][17] + xor_out[18][10][17] + xor_out[19][10][17];
assign sum_out[4][10][17] = xor_out[20][10][17] + xor_out[21][10][17] + xor_out[22][10][17] + xor_out[23][10][17] + xor_out[24][10][17];
assign sum_out[5][10][17] = xor_out[25][10][17] + xor_out[26][10][17] + xor_out[27][10][17] + xor_out[28][10][17] + xor_out[29][10][17];
assign sum_out[6][10][17] = xor_out[30][10][17] + xor_out[31][10][17] + xor_out[32][10][17] + xor_out[33][10][17] + xor_out[34][10][17];
assign sum_out[7][10][17] = xor_out[35][10][17] + xor_out[36][10][17] + xor_out[37][10][17] + xor_out[38][10][17] + xor_out[39][10][17];
assign sum_out[8][10][17] = xor_out[40][10][17] + xor_out[41][10][17] + xor_out[42][10][17] + xor_out[43][10][17] + xor_out[44][10][17];
assign sum_out[9][10][17] = xor_out[45][10][17] + xor_out[46][10][17] + xor_out[47][10][17] + xor_out[48][10][17] + xor_out[49][10][17];
assign sum_out[10][10][17] = xor_out[50][10][17] + xor_out[51][10][17] + xor_out[52][10][17] + xor_out[53][10][17] + xor_out[54][10][17];
assign sum_out[11][10][17] = xor_out[55][10][17] + xor_out[56][10][17] + xor_out[57][10][17] + xor_out[58][10][17] + xor_out[59][10][17];
assign sum_out[12][10][17] = xor_out[60][10][17] + xor_out[61][10][17] + xor_out[62][10][17] + xor_out[63][10][17] + xor_out[64][10][17];
assign sum_out[13][10][17] = xor_out[65][10][17] + xor_out[66][10][17] + xor_out[67][10][17] + xor_out[68][10][17] + xor_out[69][10][17];
assign sum_out[14][10][17] = xor_out[70][10][17] + xor_out[71][10][17] + xor_out[72][10][17] + xor_out[73][10][17] + xor_out[74][10][17];
assign sum_out[15][10][17] = xor_out[75][10][17] + xor_out[76][10][17] + xor_out[77][10][17] + xor_out[78][10][17] + xor_out[79][10][17];
assign sum_out[16][10][17] = xor_out[80][10][17] + xor_out[81][10][17] + xor_out[82][10][17] + xor_out[83][10][17] + xor_out[84][10][17];
assign sum_out[17][10][17] = xor_out[85][10][17] + xor_out[86][10][17] + xor_out[87][10][17] + xor_out[88][10][17] + xor_out[89][10][17];
assign sum_out[18][10][17] = xor_out[90][10][17] + xor_out[91][10][17] + xor_out[92][10][17] + xor_out[93][10][17] + xor_out[94][10][17];
assign sum_out[19][10][17] = xor_out[95][10][17] + xor_out[96][10][17] + xor_out[97][10][17] + xor_out[98][10][17] + xor_out[99][10][17];

assign sum_out[0][10][18] = xor_out[0][10][18] + xor_out[1][10][18] + xor_out[2][10][18] + xor_out[3][10][18] + xor_out[4][10][18];
assign sum_out[1][10][18] = xor_out[5][10][18] + xor_out[6][10][18] + xor_out[7][10][18] + xor_out[8][10][18] + xor_out[9][10][18];
assign sum_out[2][10][18] = xor_out[10][10][18] + xor_out[11][10][18] + xor_out[12][10][18] + xor_out[13][10][18] + xor_out[14][10][18];
assign sum_out[3][10][18] = xor_out[15][10][18] + xor_out[16][10][18] + xor_out[17][10][18] + xor_out[18][10][18] + xor_out[19][10][18];
assign sum_out[4][10][18] = xor_out[20][10][18] + xor_out[21][10][18] + xor_out[22][10][18] + xor_out[23][10][18] + xor_out[24][10][18];
assign sum_out[5][10][18] = xor_out[25][10][18] + xor_out[26][10][18] + xor_out[27][10][18] + xor_out[28][10][18] + xor_out[29][10][18];
assign sum_out[6][10][18] = xor_out[30][10][18] + xor_out[31][10][18] + xor_out[32][10][18] + xor_out[33][10][18] + xor_out[34][10][18];
assign sum_out[7][10][18] = xor_out[35][10][18] + xor_out[36][10][18] + xor_out[37][10][18] + xor_out[38][10][18] + xor_out[39][10][18];
assign sum_out[8][10][18] = xor_out[40][10][18] + xor_out[41][10][18] + xor_out[42][10][18] + xor_out[43][10][18] + xor_out[44][10][18];
assign sum_out[9][10][18] = xor_out[45][10][18] + xor_out[46][10][18] + xor_out[47][10][18] + xor_out[48][10][18] + xor_out[49][10][18];
assign sum_out[10][10][18] = xor_out[50][10][18] + xor_out[51][10][18] + xor_out[52][10][18] + xor_out[53][10][18] + xor_out[54][10][18];
assign sum_out[11][10][18] = xor_out[55][10][18] + xor_out[56][10][18] + xor_out[57][10][18] + xor_out[58][10][18] + xor_out[59][10][18];
assign sum_out[12][10][18] = xor_out[60][10][18] + xor_out[61][10][18] + xor_out[62][10][18] + xor_out[63][10][18] + xor_out[64][10][18];
assign sum_out[13][10][18] = xor_out[65][10][18] + xor_out[66][10][18] + xor_out[67][10][18] + xor_out[68][10][18] + xor_out[69][10][18];
assign sum_out[14][10][18] = xor_out[70][10][18] + xor_out[71][10][18] + xor_out[72][10][18] + xor_out[73][10][18] + xor_out[74][10][18];
assign sum_out[15][10][18] = xor_out[75][10][18] + xor_out[76][10][18] + xor_out[77][10][18] + xor_out[78][10][18] + xor_out[79][10][18];
assign sum_out[16][10][18] = xor_out[80][10][18] + xor_out[81][10][18] + xor_out[82][10][18] + xor_out[83][10][18] + xor_out[84][10][18];
assign sum_out[17][10][18] = xor_out[85][10][18] + xor_out[86][10][18] + xor_out[87][10][18] + xor_out[88][10][18] + xor_out[89][10][18];
assign sum_out[18][10][18] = xor_out[90][10][18] + xor_out[91][10][18] + xor_out[92][10][18] + xor_out[93][10][18] + xor_out[94][10][18];
assign sum_out[19][10][18] = xor_out[95][10][18] + xor_out[96][10][18] + xor_out[97][10][18] + xor_out[98][10][18] + xor_out[99][10][18];

assign sum_out[0][10][19] = xor_out[0][10][19] + xor_out[1][10][19] + xor_out[2][10][19] + xor_out[3][10][19] + xor_out[4][10][19];
assign sum_out[1][10][19] = xor_out[5][10][19] + xor_out[6][10][19] + xor_out[7][10][19] + xor_out[8][10][19] + xor_out[9][10][19];
assign sum_out[2][10][19] = xor_out[10][10][19] + xor_out[11][10][19] + xor_out[12][10][19] + xor_out[13][10][19] + xor_out[14][10][19];
assign sum_out[3][10][19] = xor_out[15][10][19] + xor_out[16][10][19] + xor_out[17][10][19] + xor_out[18][10][19] + xor_out[19][10][19];
assign sum_out[4][10][19] = xor_out[20][10][19] + xor_out[21][10][19] + xor_out[22][10][19] + xor_out[23][10][19] + xor_out[24][10][19];
assign sum_out[5][10][19] = xor_out[25][10][19] + xor_out[26][10][19] + xor_out[27][10][19] + xor_out[28][10][19] + xor_out[29][10][19];
assign sum_out[6][10][19] = xor_out[30][10][19] + xor_out[31][10][19] + xor_out[32][10][19] + xor_out[33][10][19] + xor_out[34][10][19];
assign sum_out[7][10][19] = xor_out[35][10][19] + xor_out[36][10][19] + xor_out[37][10][19] + xor_out[38][10][19] + xor_out[39][10][19];
assign sum_out[8][10][19] = xor_out[40][10][19] + xor_out[41][10][19] + xor_out[42][10][19] + xor_out[43][10][19] + xor_out[44][10][19];
assign sum_out[9][10][19] = xor_out[45][10][19] + xor_out[46][10][19] + xor_out[47][10][19] + xor_out[48][10][19] + xor_out[49][10][19];
assign sum_out[10][10][19] = xor_out[50][10][19] + xor_out[51][10][19] + xor_out[52][10][19] + xor_out[53][10][19] + xor_out[54][10][19];
assign sum_out[11][10][19] = xor_out[55][10][19] + xor_out[56][10][19] + xor_out[57][10][19] + xor_out[58][10][19] + xor_out[59][10][19];
assign sum_out[12][10][19] = xor_out[60][10][19] + xor_out[61][10][19] + xor_out[62][10][19] + xor_out[63][10][19] + xor_out[64][10][19];
assign sum_out[13][10][19] = xor_out[65][10][19] + xor_out[66][10][19] + xor_out[67][10][19] + xor_out[68][10][19] + xor_out[69][10][19];
assign sum_out[14][10][19] = xor_out[70][10][19] + xor_out[71][10][19] + xor_out[72][10][19] + xor_out[73][10][19] + xor_out[74][10][19];
assign sum_out[15][10][19] = xor_out[75][10][19] + xor_out[76][10][19] + xor_out[77][10][19] + xor_out[78][10][19] + xor_out[79][10][19];
assign sum_out[16][10][19] = xor_out[80][10][19] + xor_out[81][10][19] + xor_out[82][10][19] + xor_out[83][10][19] + xor_out[84][10][19];
assign sum_out[17][10][19] = xor_out[85][10][19] + xor_out[86][10][19] + xor_out[87][10][19] + xor_out[88][10][19] + xor_out[89][10][19];
assign sum_out[18][10][19] = xor_out[90][10][19] + xor_out[91][10][19] + xor_out[92][10][19] + xor_out[93][10][19] + xor_out[94][10][19];
assign sum_out[19][10][19] = xor_out[95][10][19] + xor_out[96][10][19] + xor_out[97][10][19] + xor_out[98][10][19] + xor_out[99][10][19];

assign sum_out[0][10][20] = xor_out[0][10][20] + xor_out[1][10][20] + xor_out[2][10][20] + xor_out[3][10][20] + xor_out[4][10][20];
assign sum_out[1][10][20] = xor_out[5][10][20] + xor_out[6][10][20] + xor_out[7][10][20] + xor_out[8][10][20] + xor_out[9][10][20];
assign sum_out[2][10][20] = xor_out[10][10][20] + xor_out[11][10][20] + xor_out[12][10][20] + xor_out[13][10][20] + xor_out[14][10][20];
assign sum_out[3][10][20] = xor_out[15][10][20] + xor_out[16][10][20] + xor_out[17][10][20] + xor_out[18][10][20] + xor_out[19][10][20];
assign sum_out[4][10][20] = xor_out[20][10][20] + xor_out[21][10][20] + xor_out[22][10][20] + xor_out[23][10][20] + xor_out[24][10][20];
assign sum_out[5][10][20] = xor_out[25][10][20] + xor_out[26][10][20] + xor_out[27][10][20] + xor_out[28][10][20] + xor_out[29][10][20];
assign sum_out[6][10][20] = xor_out[30][10][20] + xor_out[31][10][20] + xor_out[32][10][20] + xor_out[33][10][20] + xor_out[34][10][20];
assign sum_out[7][10][20] = xor_out[35][10][20] + xor_out[36][10][20] + xor_out[37][10][20] + xor_out[38][10][20] + xor_out[39][10][20];
assign sum_out[8][10][20] = xor_out[40][10][20] + xor_out[41][10][20] + xor_out[42][10][20] + xor_out[43][10][20] + xor_out[44][10][20];
assign sum_out[9][10][20] = xor_out[45][10][20] + xor_out[46][10][20] + xor_out[47][10][20] + xor_out[48][10][20] + xor_out[49][10][20];
assign sum_out[10][10][20] = xor_out[50][10][20] + xor_out[51][10][20] + xor_out[52][10][20] + xor_out[53][10][20] + xor_out[54][10][20];
assign sum_out[11][10][20] = xor_out[55][10][20] + xor_out[56][10][20] + xor_out[57][10][20] + xor_out[58][10][20] + xor_out[59][10][20];
assign sum_out[12][10][20] = xor_out[60][10][20] + xor_out[61][10][20] + xor_out[62][10][20] + xor_out[63][10][20] + xor_out[64][10][20];
assign sum_out[13][10][20] = xor_out[65][10][20] + xor_out[66][10][20] + xor_out[67][10][20] + xor_out[68][10][20] + xor_out[69][10][20];
assign sum_out[14][10][20] = xor_out[70][10][20] + xor_out[71][10][20] + xor_out[72][10][20] + xor_out[73][10][20] + xor_out[74][10][20];
assign sum_out[15][10][20] = xor_out[75][10][20] + xor_out[76][10][20] + xor_out[77][10][20] + xor_out[78][10][20] + xor_out[79][10][20];
assign sum_out[16][10][20] = xor_out[80][10][20] + xor_out[81][10][20] + xor_out[82][10][20] + xor_out[83][10][20] + xor_out[84][10][20];
assign sum_out[17][10][20] = xor_out[85][10][20] + xor_out[86][10][20] + xor_out[87][10][20] + xor_out[88][10][20] + xor_out[89][10][20];
assign sum_out[18][10][20] = xor_out[90][10][20] + xor_out[91][10][20] + xor_out[92][10][20] + xor_out[93][10][20] + xor_out[94][10][20];
assign sum_out[19][10][20] = xor_out[95][10][20] + xor_out[96][10][20] + xor_out[97][10][20] + xor_out[98][10][20] + xor_out[99][10][20];

assign sum_out[0][10][21] = xor_out[0][10][21] + xor_out[1][10][21] + xor_out[2][10][21] + xor_out[3][10][21] + xor_out[4][10][21];
assign sum_out[1][10][21] = xor_out[5][10][21] + xor_out[6][10][21] + xor_out[7][10][21] + xor_out[8][10][21] + xor_out[9][10][21];
assign sum_out[2][10][21] = xor_out[10][10][21] + xor_out[11][10][21] + xor_out[12][10][21] + xor_out[13][10][21] + xor_out[14][10][21];
assign sum_out[3][10][21] = xor_out[15][10][21] + xor_out[16][10][21] + xor_out[17][10][21] + xor_out[18][10][21] + xor_out[19][10][21];
assign sum_out[4][10][21] = xor_out[20][10][21] + xor_out[21][10][21] + xor_out[22][10][21] + xor_out[23][10][21] + xor_out[24][10][21];
assign sum_out[5][10][21] = xor_out[25][10][21] + xor_out[26][10][21] + xor_out[27][10][21] + xor_out[28][10][21] + xor_out[29][10][21];
assign sum_out[6][10][21] = xor_out[30][10][21] + xor_out[31][10][21] + xor_out[32][10][21] + xor_out[33][10][21] + xor_out[34][10][21];
assign sum_out[7][10][21] = xor_out[35][10][21] + xor_out[36][10][21] + xor_out[37][10][21] + xor_out[38][10][21] + xor_out[39][10][21];
assign sum_out[8][10][21] = xor_out[40][10][21] + xor_out[41][10][21] + xor_out[42][10][21] + xor_out[43][10][21] + xor_out[44][10][21];
assign sum_out[9][10][21] = xor_out[45][10][21] + xor_out[46][10][21] + xor_out[47][10][21] + xor_out[48][10][21] + xor_out[49][10][21];
assign sum_out[10][10][21] = xor_out[50][10][21] + xor_out[51][10][21] + xor_out[52][10][21] + xor_out[53][10][21] + xor_out[54][10][21];
assign sum_out[11][10][21] = xor_out[55][10][21] + xor_out[56][10][21] + xor_out[57][10][21] + xor_out[58][10][21] + xor_out[59][10][21];
assign sum_out[12][10][21] = xor_out[60][10][21] + xor_out[61][10][21] + xor_out[62][10][21] + xor_out[63][10][21] + xor_out[64][10][21];
assign sum_out[13][10][21] = xor_out[65][10][21] + xor_out[66][10][21] + xor_out[67][10][21] + xor_out[68][10][21] + xor_out[69][10][21];
assign sum_out[14][10][21] = xor_out[70][10][21] + xor_out[71][10][21] + xor_out[72][10][21] + xor_out[73][10][21] + xor_out[74][10][21];
assign sum_out[15][10][21] = xor_out[75][10][21] + xor_out[76][10][21] + xor_out[77][10][21] + xor_out[78][10][21] + xor_out[79][10][21];
assign sum_out[16][10][21] = xor_out[80][10][21] + xor_out[81][10][21] + xor_out[82][10][21] + xor_out[83][10][21] + xor_out[84][10][21];
assign sum_out[17][10][21] = xor_out[85][10][21] + xor_out[86][10][21] + xor_out[87][10][21] + xor_out[88][10][21] + xor_out[89][10][21];
assign sum_out[18][10][21] = xor_out[90][10][21] + xor_out[91][10][21] + xor_out[92][10][21] + xor_out[93][10][21] + xor_out[94][10][21];
assign sum_out[19][10][21] = xor_out[95][10][21] + xor_out[96][10][21] + xor_out[97][10][21] + xor_out[98][10][21] + xor_out[99][10][21];

assign sum_out[0][10][22] = xor_out[0][10][22] + xor_out[1][10][22] + xor_out[2][10][22] + xor_out[3][10][22] + xor_out[4][10][22];
assign sum_out[1][10][22] = xor_out[5][10][22] + xor_out[6][10][22] + xor_out[7][10][22] + xor_out[8][10][22] + xor_out[9][10][22];
assign sum_out[2][10][22] = xor_out[10][10][22] + xor_out[11][10][22] + xor_out[12][10][22] + xor_out[13][10][22] + xor_out[14][10][22];
assign sum_out[3][10][22] = xor_out[15][10][22] + xor_out[16][10][22] + xor_out[17][10][22] + xor_out[18][10][22] + xor_out[19][10][22];
assign sum_out[4][10][22] = xor_out[20][10][22] + xor_out[21][10][22] + xor_out[22][10][22] + xor_out[23][10][22] + xor_out[24][10][22];
assign sum_out[5][10][22] = xor_out[25][10][22] + xor_out[26][10][22] + xor_out[27][10][22] + xor_out[28][10][22] + xor_out[29][10][22];
assign sum_out[6][10][22] = xor_out[30][10][22] + xor_out[31][10][22] + xor_out[32][10][22] + xor_out[33][10][22] + xor_out[34][10][22];
assign sum_out[7][10][22] = xor_out[35][10][22] + xor_out[36][10][22] + xor_out[37][10][22] + xor_out[38][10][22] + xor_out[39][10][22];
assign sum_out[8][10][22] = xor_out[40][10][22] + xor_out[41][10][22] + xor_out[42][10][22] + xor_out[43][10][22] + xor_out[44][10][22];
assign sum_out[9][10][22] = xor_out[45][10][22] + xor_out[46][10][22] + xor_out[47][10][22] + xor_out[48][10][22] + xor_out[49][10][22];
assign sum_out[10][10][22] = xor_out[50][10][22] + xor_out[51][10][22] + xor_out[52][10][22] + xor_out[53][10][22] + xor_out[54][10][22];
assign sum_out[11][10][22] = xor_out[55][10][22] + xor_out[56][10][22] + xor_out[57][10][22] + xor_out[58][10][22] + xor_out[59][10][22];
assign sum_out[12][10][22] = xor_out[60][10][22] + xor_out[61][10][22] + xor_out[62][10][22] + xor_out[63][10][22] + xor_out[64][10][22];
assign sum_out[13][10][22] = xor_out[65][10][22] + xor_out[66][10][22] + xor_out[67][10][22] + xor_out[68][10][22] + xor_out[69][10][22];
assign sum_out[14][10][22] = xor_out[70][10][22] + xor_out[71][10][22] + xor_out[72][10][22] + xor_out[73][10][22] + xor_out[74][10][22];
assign sum_out[15][10][22] = xor_out[75][10][22] + xor_out[76][10][22] + xor_out[77][10][22] + xor_out[78][10][22] + xor_out[79][10][22];
assign sum_out[16][10][22] = xor_out[80][10][22] + xor_out[81][10][22] + xor_out[82][10][22] + xor_out[83][10][22] + xor_out[84][10][22];
assign sum_out[17][10][22] = xor_out[85][10][22] + xor_out[86][10][22] + xor_out[87][10][22] + xor_out[88][10][22] + xor_out[89][10][22];
assign sum_out[18][10][22] = xor_out[90][10][22] + xor_out[91][10][22] + xor_out[92][10][22] + xor_out[93][10][22] + xor_out[94][10][22];
assign sum_out[19][10][22] = xor_out[95][10][22] + xor_out[96][10][22] + xor_out[97][10][22] + xor_out[98][10][22] + xor_out[99][10][22];

assign sum_out[0][10][23] = xor_out[0][10][23] + xor_out[1][10][23] + xor_out[2][10][23] + xor_out[3][10][23] + xor_out[4][10][23];
assign sum_out[1][10][23] = xor_out[5][10][23] + xor_out[6][10][23] + xor_out[7][10][23] + xor_out[8][10][23] + xor_out[9][10][23];
assign sum_out[2][10][23] = xor_out[10][10][23] + xor_out[11][10][23] + xor_out[12][10][23] + xor_out[13][10][23] + xor_out[14][10][23];
assign sum_out[3][10][23] = xor_out[15][10][23] + xor_out[16][10][23] + xor_out[17][10][23] + xor_out[18][10][23] + xor_out[19][10][23];
assign sum_out[4][10][23] = xor_out[20][10][23] + xor_out[21][10][23] + xor_out[22][10][23] + xor_out[23][10][23] + xor_out[24][10][23];
assign sum_out[5][10][23] = xor_out[25][10][23] + xor_out[26][10][23] + xor_out[27][10][23] + xor_out[28][10][23] + xor_out[29][10][23];
assign sum_out[6][10][23] = xor_out[30][10][23] + xor_out[31][10][23] + xor_out[32][10][23] + xor_out[33][10][23] + xor_out[34][10][23];
assign sum_out[7][10][23] = xor_out[35][10][23] + xor_out[36][10][23] + xor_out[37][10][23] + xor_out[38][10][23] + xor_out[39][10][23];
assign sum_out[8][10][23] = xor_out[40][10][23] + xor_out[41][10][23] + xor_out[42][10][23] + xor_out[43][10][23] + xor_out[44][10][23];
assign sum_out[9][10][23] = xor_out[45][10][23] + xor_out[46][10][23] + xor_out[47][10][23] + xor_out[48][10][23] + xor_out[49][10][23];
assign sum_out[10][10][23] = xor_out[50][10][23] + xor_out[51][10][23] + xor_out[52][10][23] + xor_out[53][10][23] + xor_out[54][10][23];
assign sum_out[11][10][23] = xor_out[55][10][23] + xor_out[56][10][23] + xor_out[57][10][23] + xor_out[58][10][23] + xor_out[59][10][23];
assign sum_out[12][10][23] = xor_out[60][10][23] + xor_out[61][10][23] + xor_out[62][10][23] + xor_out[63][10][23] + xor_out[64][10][23];
assign sum_out[13][10][23] = xor_out[65][10][23] + xor_out[66][10][23] + xor_out[67][10][23] + xor_out[68][10][23] + xor_out[69][10][23];
assign sum_out[14][10][23] = xor_out[70][10][23] + xor_out[71][10][23] + xor_out[72][10][23] + xor_out[73][10][23] + xor_out[74][10][23];
assign sum_out[15][10][23] = xor_out[75][10][23] + xor_out[76][10][23] + xor_out[77][10][23] + xor_out[78][10][23] + xor_out[79][10][23];
assign sum_out[16][10][23] = xor_out[80][10][23] + xor_out[81][10][23] + xor_out[82][10][23] + xor_out[83][10][23] + xor_out[84][10][23];
assign sum_out[17][10][23] = xor_out[85][10][23] + xor_out[86][10][23] + xor_out[87][10][23] + xor_out[88][10][23] + xor_out[89][10][23];
assign sum_out[18][10][23] = xor_out[90][10][23] + xor_out[91][10][23] + xor_out[92][10][23] + xor_out[93][10][23] + xor_out[94][10][23];
assign sum_out[19][10][23] = xor_out[95][10][23] + xor_out[96][10][23] + xor_out[97][10][23] + xor_out[98][10][23] + xor_out[99][10][23];

assign sum_out[0][11][0] = xor_out[0][11][0] + xor_out[1][11][0] + xor_out[2][11][0] + xor_out[3][11][0] + xor_out[4][11][0];
assign sum_out[1][11][0] = xor_out[5][11][0] + xor_out[6][11][0] + xor_out[7][11][0] + xor_out[8][11][0] + xor_out[9][11][0];
assign sum_out[2][11][0] = xor_out[10][11][0] + xor_out[11][11][0] + xor_out[12][11][0] + xor_out[13][11][0] + xor_out[14][11][0];
assign sum_out[3][11][0] = xor_out[15][11][0] + xor_out[16][11][0] + xor_out[17][11][0] + xor_out[18][11][0] + xor_out[19][11][0];
assign sum_out[4][11][0] = xor_out[20][11][0] + xor_out[21][11][0] + xor_out[22][11][0] + xor_out[23][11][0] + xor_out[24][11][0];
assign sum_out[5][11][0] = xor_out[25][11][0] + xor_out[26][11][0] + xor_out[27][11][0] + xor_out[28][11][0] + xor_out[29][11][0];
assign sum_out[6][11][0] = xor_out[30][11][0] + xor_out[31][11][0] + xor_out[32][11][0] + xor_out[33][11][0] + xor_out[34][11][0];
assign sum_out[7][11][0] = xor_out[35][11][0] + xor_out[36][11][0] + xor_out[37][11][0] + xor_out[38][11][0] + xor_out[39][11][0];
assign sum_out[8][11][0] = xor_out[40][11][0] + xor_out[41][11][0] + xor_out[42][11][0] + xor_out[43][11][0] + xor_out[44][11][0];
assign sum_out[9][11][0] = xor_out[45][11][0] + xor_out[46][11][0] + xor_out[47][11][0] + xor_out[48][11][0] + xor_out[49][11][0];
assign sum_out[10][11][0] = xor_out[50][11][0] + xor_out[51][11][0] + xor_out[52][11][0] + xor_out[53][11][0] + xor_out[54][11][0];
assign sum_out[11][11][0] = xor_out[55][11][0] + xor_out[56][11][0] + xor_out[57][11][0] + xor_out[58][11][0] + xor_out[59][11][0];
assign sum_out[12][11][0] = xor_out[60][11][0] + xor_out[61][11][0] + xor_out[62][11][0] + xor_out[63][11][0] + xor_out[64][11][0];
assign sum_out[13][11][0] = xor_out[65][11][0] + xor_out[66][11][0] + xor_out[67][11][0] + xor_out[68][11][0] + xor_out[69][11][0];
assign sum_out[14][11][0] = xor_out[70][11][0] + xor_out[71][11][0] + xor_out[72][11][0] + xor_out[73][11][0] + xor_out[74][11][0];
assign sum_out[15][11][0] = xor_out[75][11][0] + xor_out[76][11][0] + xor_out[77][11][0] + xor_out[78][11][0] + xor_out[79][11][0];
assign sum_out[16][11][0] = xor_out[80][11][0] + xor_out[81][11][0] + xor_out[82][11][0] + xor_out[83][11][0] + xor_out[84][11][0];
assign sum_out[17][11][0] = xor_out[85][11][0] + xor_out[86][11][0] + xor_out[87][11][0] + xor_out[88][11][0] + xor_out[89][11][0];
assign sum_out[18][11][0] = xor_out[90][11][0] + xor_out[91][11][0] + xor_out[92][11][0] + xor_out[93][11][0] + xor_out[94][11][0];
assign sum_out[19][11][0] = xor_out[95][11][0] + xor_out[96][11][0] + xor_out[97][11][0] + xor_out[98][11][0] + xor_out[99][11][0];

assign sum_out[0][11][1] = xor_out[0][11][1] + xor_out[1][11][1] + xor_out[2][11][1] + xor_out[3][11][1] + xor_out[4][11][1];
assign sum_out[1][11][1] = xor_out[5][11][1] + xor_out[6][11][1] + xor_out[7][11][1] + xor_out[8][11][1] + xor_out[9][11][1];
assign sum_out[2][11][1] = xor_out[10][11][1] + xor_out[11][11][1] + xor_out[12][11][1] + xor_out[13][11][1] + xor_out[14][11][1];
assign sum_out[3][11][1] = xor_out[15][11][1] + xor_out[16][11][1] + xor_out[17][11][1] + xor_out[18][11][1] + xor_out[19][11][1];
assign sum_out[4][11][1] = xor_out[20][11][1] + xor_out[21][11][1] + xor_out[22][11][1] + xor_out[23][11][1] + xor_out[24][11][1];
assign sum_out[5][11][1] = xor_out[25][11][1] + xor_out[26][11][1] + xor_out[27][11][1] + xor_out[28][11][1] + xor_out[29][11][1];
assign sum_out[6][11][1] = xor_out[30][11][1] + xor_out[31][11][1] + xor_out[32][11][1] + xor_out[33][11][1] + xor_out[34][11][1];
assign sum_out[7][11][1] = xor_out[35][11][1] + xor_out[36][11][1] + xor_out[37][11][1] + xor_out[38][11][1] + xor_out[39][11][1];
assign sum_out[8][11][1] = xor_out[40][11][1] + xor_out[41][11][1] + xor_out[42][11][1] + xor_out[43][11][1] + xor_out[44][11][1];
assign sum_out[9][11][1] = xor_out[45][11][1] + xor_out[46][11][1] + xor_out[47][11][1] + xor_out[48][11][1] + xor_out[49][11][1];
assign sum_out[10][11][1] = xor_out[50][11][1] + xor_out[51][11][1] + xor_out[52][11][1] + xor_out[53][11][1] + xor_out[54][11][1];
assign sum_out[11][11][1] = xor_out[55][11][1] + xor_out[56][11][1] + xor_out[57][11][1] + xor_out[58][11][1] + xor_out[59][11][1];
assign sum_out[12][11][1] = xor_out[60][11][1] + xor_out[61][11][1] + xor_out[62][11][1] + xor_out[63][11][1] + xor_out[64][11][1];
assign sum_out[13][11][1] = xor_out[65][11][1] + xor_out[66][11][1] + xor_out[67][11][1] + xor_out[68][11][1] + xor_out[69][11][1];
assign sum_out[14][11][1] = xor_out[70][11][1] + xor_out[71][11][1] + xor_out[72][11][1] + xor_out[73][11][1] + xor_out[74][11][1];
assign sum_out[15][11][1] = xor_out[75][11][1] + xor_out[76][11][1] + xor_out[77][11][1] + xor_out[78][11][1] + xor_out[79][11][1];
assign sum_out[16][11][1] = xor_out[80][11][1] + xor_out[81][11][1] + xor_out[82][11][1] + xor_out[83][11][1] + xor_out[84][11][1];
assign sum_out[17][11][1] = xor_out[85][11][1] + xor_out[86][11][1] + xor_out[87][11][1] + xor_out[88][11][1] + xor_out[89][11][1];
assign sum_out[18][11][1] = xor_out[90][11][1] + xor_out[91][11][1] + xor_out[92][11][1] + xor_out[93][11][1] + xor_out[94][11][1];
assign sum_out[19][11][1] = xor_out[95][11][1] + xor_out[96][11][1] + xor_out[97][11][1] + xor_out[98][11][1] + xor_out[99][11][1];

assign sum_out[0][11][2] = xor_out[0][11][2] + xor_out[1][11][2] + xor_out[2][11][2] + xor_out[3][11][2] + xor_out[4][11][2];
assign sum_out[1][11][2] = xor_out[5][11][2] + xor_out[6][11][2] + xor_out[7][11][2] + xor_out[8][11][2] + xor_out[9][11][2];
assign sum_out[2][11][2] = xor_out[10][11][2] + xor_out[11][11][2] + xor_out[12][11][2] + xor_out[13][11][2] + xor_out[14][11][2];
assign sum_out[3][11][2] = xor_out[15][11][2] + xor_out[16][11][2] + xor_out[17][11][2] + xor_out[18][11][2] + xor_out[19][11][2];
assign sum_out[4][11][2] = xor_out[20][11][2] + xor_out[21][11][2] + xor_out[22][11][2] + xor_out[23][11][2] + xor_out[24][11][2];
assign sum_out[5][11][2] = xor_out[25][11][2] + xor_out[26][11][2] + xor_out[27][11][2] + xor_out[28][11][2] + xor_out[29][11][2];
assign sum_out[6][11][2] = xor_out[30][11][2] + xor_out[31][11][2] + xor_out[32][11][2] + xor_out[33][11][2] + xor_out[34][11][2];
assign sum_out[7][11][2] = xor_out[35][11][2] + xor_out[36][11][2] + xor_out[37][11][2] + xor_out[38][11][2] + xor_out[39][11][2];
assign sum_out[8][11][2] = xor_out[40][11][2] + xor_out[41][11][2] + xor_out[42][11][2] + xor_out[43][11][2] + xor_out[44][11][2];
assign sum_out[9][11][2] = xor_out[45][11][2] + xor_out[46][11][2] + xor_out[47][11][2] + xor_out[48][11][2] + xor_out[49][11][2];
assign sum_out[10][11][2] = xor_out[50][11][2] + xor_out[51][11][2] + xor_out[52][11][2] + xor_out[53][11][2] + xor_out[54][11][2];
assign sum_out[11][11][2] = xor_out[55][11][2] + xor_out[56][11][2] + xor_out[57][11][2] + xor_out[58][11][2] + xor_out[59][11][2];
assign sum_out[12][11][2] = xor_out[60][11][2] + xor_out[61][11][2] + xor_out[62][11][2] + xor_out[63][11][2] + xor_out[64][11][2];
assign sum_out[13][11][2] = xor_out[65][11][2] + xor_out[66][11][2] + xor_out[67][11][2] + xor_out[68][11][2] + xor_out[69][11][2];
assign sum_out[14][11][2] = xor_out[70][11][2] + xor_out[71][11][2] + xor_out[72][11][2] + xor_out[73][11][2] + xor_out[74][11][2];
assign sum_out[15][11][2] = xor_out[75][11][2] + xor_out[76][11][2] + xor_out[77][11][2] + xor_out[78][11][2] + xor_out[79][11][2];
assign sum_out[16][11][2] = xor_out[80][11][2] + xor_out[81][11][2] + xor_out[82][11][2] + xor_out[83][11][2] + xor_out[84][11][2];
assign sum_out[17][11][2] = xor_out[85][11][2] + xor_out[86][11][2] + xor_out[87][11][2] + xor_out[88][11][2] + xor_out[89][11][2];
assign sum_out[18][11][2] = xor_out[90][11][2] + xor_out[91][11][2] + xor_out[92][11][2] + xor_out[93][11][2] + xor_out[94][11][2];
assign sum_out[19][11][2] = xor_out[95][11][2] + xor_out[96][11][2] + xor_out[97][11][2] + xor_out[98][11][2] + xor_out[99][11][2];

assign sum_out[0][11][3] = xor_out[0][11][3] + xor_out[1][11][3] + xor_out[2][11][3] + xor_out[3][11][3] + xor_out[4][11][3];
assign sum_out[1][11][3] = xor_out[5][11][3] + xor_out[6][11][3] + xor_out[7][11][3] + xor_out[8][11][3] + xor_out[9][11][3];
assign sum_out[2][11][3] = xor_out[10][11][3] + xor_out[11][11][3] + xor_out[12][11][3] + xor_out[13][11][3] + xor_out[14][11][3];
assign sum_out[3][11][3] = xor_out[15][11][3] + xor_out[16][11][3] + xor_out[17][11][3] + xor_out[18][11][3] + xor_out[19][11][3];
assign sum_out[4][11][3] = xor_out[20][11][3] + xor_out[21][11][3] + xor_out[22][11][3] + xor_out[23][11][3] + xor_out[24][11][3];
assign sum_out[5][11][3] = xor_out[25][11][3] + xor_out[26][11][3] + xor_out[27][11][3] + xor_out[28][11][3] + xor_out[29][11][3];
assign sum_out[6][11][3] = xor_out[30][11][3] + xor_out[31][11][3] + xor_out[32][11][3] + xor_out[33][11][3] + xor_out[34][11][3];
assign sum_out[7][11][3] = xor_out[35][11][3] + xor_out[36][11][3] + xor_out[37][11][3] + xor_out[38][11][3] + xor_out[39][11][3];
assign sum_out[8][11][3] = xor_out[40][11][3] + xor_out[41][11][3] + xor_out[42][11][3] + xor_out[43][11][3] + xor_out[44][11][3];
assign sum_out[9][11][3] = xor_out[45][11][3] + xor_out[46][11][3] + xor_out[47][11][3] + xor_out[48][11][3] + xor_out[49][11][3];
assign sum_out[10][11][3] = xor_out[50][11][3] + xor_out[51][11][3] + xor_out[52][11][3] + xor_out[53][11][3] + xor_out[54][11][3];
assign sum_out[11][11][3] = xor_out[55][11][3] + xor_out[56][11][3] + xor_out[57][11][3] + xor_out[58][11][3] + xor_out[59][11][3];
assign sum_out[12][11][3] = xor_out[60][11][3] + xor_out[61][11][3] + xor_out[62][11][3] + xor_out[63][11][3] + xor_out[64][11][3];
assign sum_out[13][11][3] = xor_out[65][11][3] + xor_out[66][11][3] + xor_out[67][11][3] + xor_out[68][11][3] + xor_out[69][11][3];
assign sum_out[14][11][3] = xor_out[70][11][3] + xor_out[71][11][3] + xor_out[72][11][3] + xor_out[73][11][3] + xor_out[74][11][3];
assign sum_out[15][11][3] = xor_out[75][11][3] + xor_out[76][11][3] + xor_out[77][11][3] + xor_out[78][11][3] + xor_out[79][11][3];
assign sum_out[16][11][3] = xor_out[80][11][3] + xor_out[81][11][3] + xor_out[82][11][3] + xor_out[83][11][3] + xor_out[84][11][3];
assign sum_out[17][11][3] = xor_out[85][11][3] + xor_out[86][11][3] + xor_out[87][11][3] + xor_out[88][11][3] + xor_out[89][11][3];
assign sum_out[18][11][3] = xor_out[90][11][3] + xor_out[91][11][3] + xor_out[92][11][3] + xor_out[93][11][3] + xor_out[94][11][3];
assign sum_out[19][11][3] = xor_out[95][11][3] + xor_out[96][11][3] + xor_out[97][11][3] + xor_out[98][11][3] + xor_out[99][11][3];

assign sum_out[0][11][4] = xor_out[0][11][4] + xor_out[1][11][4] + xor_out[2][11][4] + xor_out[3][11][4] + xor_out[4][11][4];
assign sum_out[1][11][4] = xor_out[5][11][4] + xor_out[6][11][4] + xor_out[7][11][4] + xor_out[8][11][4] + xor_out[9][11][4];
assign sum_out[2][11][4] = xor_out[10][11][4] + xor_out[11][11][4] + xor_out[12][11][4] + xor_out[13][11][4] + xor_out[14][11][4];
assign sum_out[3][11][4] = xor_out[15][11][4] + xor_out[16][11][4] + xor_out[17][11][4] + xor_out[18][11][4] + xor_out[19][11][4];
assign sum_out[4][11][4] = xor_out[20][11][4] + xor_out[21][11][4] + xor_out[22][11][4] + xor_out[23][11][4] + xor_out[24][11][4];
assign sum_out[5][11][4] = xor_out[25][11][4] + xor_out[26][11][4] + xor_out[27][11][4] + xor_out[28][11][4] + xor_out[29][11][4];
assign sum_out[6][11][4] = xor_out[30][11][4] + xor_out[31][11][4] + xor_out[32][11][4] + xor_out[33][11][4] + xor_out[34][11][4];
assign sum_out[7][11][4] = xor_out[35][11][4] + xor_out[36][11][4] + xor_out[37][11][4] + xor_out[38][11][4] + xor_out[39][11][4];
assign sum_out[8][11][4] = xor_out[40][11][4] + xor_out[41][11][4] + xor_out[42][11][4] + xor_out[43][11][4] + xor_out[44][11][4];
assign sum_out[9][11][4] = xor_out[45][11][4] + xor_out[46][11][4] + xor_out[47][11][4] + xor_out[48][11][4] + xor_out[49][11][4];
assign sum_out[10][11][4] = xor_out[50][11][4] + xor_out[51][11][4] + xor_out[52][11][4] + xor_out[53][11][4] + xor_out[54][11][4];
assign sum_out[11][11][4] = xor_out[55][11][4] + xor_out[56][11][4] + xor_out[57][11][4] + xor_out[58][11][4] + xor_out[59][11][4];
assign sum_out[12][11][4] = xor_out[60][11][4] + xor_out[61][11][4] + xor_out[62][11][4] + xor_out[63][11][4] + xor_out[64][11][4];
assign sum_out[13][11][4] = xor_out[65][11][4] + xor_out[66][11][4] + xor_out[67][11][4] + xor_out[68][11][4] + xor_out[69][11][4];
assign sum_out[14][11][4] = xor_out[70][11][4] + xor_out[71][11][4] + xor_out[72][11][4] + xor_out[73][11][4] + xor_out[74][11][4];
assign sum_out[15][11][4] = xor_out[75][11][4] + xor_out[76][11][4] + xor_out[77][11][4] + xor_out[78][11][4] + xor_out[79][11][4];
assign sum_out[16][11][4] = xor_out[80][11][4] + xor_out[81][11][4] + xor_out[82][11][4] + xor_out[83][11][4] + xor_out[84][11][4];
assign sum_out[17][11][4] = xor_out[85][11][4] + xor_out[86][11][4] + xor_out[87][11][4] + xor_out[88][11][4] + xor_out[89][11][4];
assign sum_out[18][11][4] = xor_out[90][11][4] + xor_out[91][11][4] + xor_out[92][11][4] + xor_out[93][11][4] + xor_out[94][11][4];
assign sum_out[19][11][4] = xor_out[95][11][4] + xor_out[96][11][4] + xor_out[97][11][4] + xor_out[98][11][4] + xor_out[99][11][4];

assign sum_out[0][11][5] = xor_out[0][11][5] + xor_out[1][11][5] + xor_out[2][11][5] + xor_out[3][11][5] + xor_out[4][11][5];
assign sum_out[1][11][5] = xor_out[5][11][5] + xor_out[6][11][5] + xor_out[7][11][5] + xor_out[8][11][5] + xor_out[9][11][5];
assign sum_out[2][11][5] = xor_out[10][11][5] + xor_out[11][11][5] + xor_out[12][11][5] + xor_out[13][11][5] + xor_out[14][11][5];
assign sum_out[3][11][5] = xor_out[15][11][5] + xor_out[16][11][5] + xor_out[17][11][5] + xor_out[18][11][5] + xor_out[19][11][5];
assign sum_out[4][11][5] = xor_out[20][11][5] + xor_out[21][11][5] + xor_out[22][11][5] + xor_out[23][11][5] + xor_out[24][11][5];
assign sum_out[5][11][5] = xor_out[25][11][5] + xor_out[26][11][5] + xor_out[27][11][5] + xor_out[28][11][5] + xor_out[29][11][5];
assign sum_out[6][11][5] = xor_out[30][11][5] + xor_out[31][11][5] + xor_out[32][11][5] + xor_out[33][11][5] + xor_out[34][11][5];
assign sum_out[7][11][5] = xor_out[35][11][5] + xor_out[36][11][5] + xor_out[37][11][5] + xor_out[38][11][5] + xor_out[39][11][5];
assign sum_out[8][11][5] = xor_out[40][11][5] + xor_out[41][11][5] + xor_out[42][11][5] + xor_out[43][11][5] + xor_out[44][11][5];
assign sum_out[9][11][5] = xor_out[45][11][5] + xor_out[46][11][5] + xor_out[47][11][5] + xor_out[48][11][5] + xor_out[49][11][5];
assign sum_out[10][11][5] = xor_out[50][11][5] + xor_out[51][11][5] + xor_out[52][11][5] + xor_out[53][11][5] + xor_out[54][11][5];
assign sum_out[11][11][5] = xor_out[55][11][5] + xor_out[56][11][5] + xor_out[57][11][5] + xor_out[58][11][5] + xor_out[59][11][5];
assign sum_out[12][11][5] = xor_out[60][11][5] + xor_out[61][11][5] + xor_out[62][11][5] + xor_out[63][11][5] + xor_out[64][11][5];
assign sum_out[13][11][5] = xor_out[65][11][5] + xor_out[66][11][5] + xor_out[67][11][5] + xor_out[68][11][5] + xor_out[69][11][5];
assign sum_out[14][11][5] = xor_out[70][11][5] + xor_out[71][11][5] + xor_out[72][11][5] + xor_out[73][11][5] + xor_out[74][11][5];
assign sum_out[15][11][5] = xor_out[75][11][5] + xor_out[76][11][5] + xor_out[77][11][5] + xor_out[78][11][5] + xor_out[79][11][5];
assign sum_out[16][11][5] = xor_out[80][11][5] + xor_out[81][11][5] + xor_out[82][11][5] + xor_out[83][11][5] + xor_out[84][11][5];
assign sum_out[17][11][5] = xor_out[85][11][5] + xor_out[86][11][5] + xor_out[87][11][5] + xor_out[88][11][5] + xor_out[89][11][5];
assign sum_out[18][11][5] = xor_out[90][11][5] + xor_out[91][11][5] + xor_out[92][11][5] + xor_out[93][11][5] + xor_out[94][11][5];
assign sum_out[19][11][5] = xor_out[95][11][5] + xor_out[96][11][5] + xor_out[97][11][5] + xor_out[98][11][5] + xor_out[99][11][5];

assign sum_out[0][11][6] = xor_out[0][11][6] + xor_out[1][11][6] + xor_out[2][11][6] + xor_out[3][11][6] + xor_out[4][11][6];
assign sum_out[1][11][6] = xor_out[5][11][6] + xor_out[6][11][6] + xor_out[7][11][6] + xor_out[8][11][6] + xor_out[9][11][6];
assign sum_out[2][11][6] = xor_out[10][11][6] + xor_out[11][11][6] + xor_out[12][11][6] + xor_out[13][11][6] + xor_out[14][11][6];
assign sum_out[3][11][6] = xor_out[15][11][6] + xor_out[16][11][6] + xor_out[17][11][6] + xor_out[18][11][6] + xor_out[19][11][6];
assign sum_out[4][11][6] = xor_out[20][11][6] + xor_out[21][11][6] + xor_out[22][11][6] + xor_out[23][11][6] + xor_out[24][11][6];
assign sum_out[5][11][6] = xor_out[25][11][6] + xor_out[26][11][6] + xor_out[27][11][6] + xor_out[28][11][6] + xor_out[29][11][6];
assign sum_out[6][11][6] = xor_out[30][11][6] + xor_out[31][11][6] + xor_out[32][11][6] + xor_out[33][11][6] + xor_out[34][11][6];
assign sum_out[7][11][6] = xor_out[35][11][6] + xor_out[36][11][6] + xor_out[37][11][6] + xor_out[38][11][6] + xor_out[39][11][6];
assign sum_out[8][11][6] = xor_out[40][11][6] + xor_out[41][11][6] + xor_out[42][11][6] + xor_out[43][11][6] + xor_out[44][11][6];
assign sum_out[9][11][6] = xor_out[45][11][6] + xor_out[46][11][6] + xor_out[47][11][6] + xor_out[48][11][6] + xor_out[49][11][6];
assign sum_out[10][11][6] = xor_out[50][11][6] + xor_out[51][11][6] + xor_out[52][11][6] + xor_out[53][11][6] + xor_out[54][11][6];
assign sum_out[11][11][6] = xor_out[55][11][6] + xor_out[56][11][6] + xor_out[57][11][6] + xor_out[58][11][6] + xor_out[59][11][6];
assign sum_out[12][11][6] = xor_out[60][11][6] + xor_out[61][11][6] + xor_out[62][11][6] + xor_out[63][11][6] + xor_out[64][11][6];
assign sum_out[13][11][6] = xor_out[65][11][6] + xor_out[66][11][6] + xor_out[67][11][6] + xor_out[68][11][6] + xor_out[69][11][6];
assign sum_out[14][11][6] = xor_out[70][11][6] + xor_out[71][11][6] + xor_out[72][11][6] + xor_out[73][11][6] + xor_out[74][11][6];
assign sum_out[15][11][6] = xor_out[75][11][6] + xor_out[76][11][6] + xor_out[77][11][6] + xor_out[78][11][6] + xor_out[79][11][6];
assign sum_out[16][11][6] = xor_out[80][11][6] + xor_out[81][11][6] + xor_out[82][11][6] + xor_out[83][11][6] + xor_out[84][11][6];
assign sum_out[17][11][6] = xor_out[85][11][6] + xor_out[86][11][6] + xor_out[87][11][6] + xor_out[88][11][6] + xor_out[89][11][6];
assign sum_out[18][11][6] = xor_out[90][11][6] + xor_out[91][11][6] + xor_out[92][11][6] + xor_out[93][11][6] + xor_out[94][11][6];
assign sum_out[19][11][6] = xor_out[95][11][6] + xor_out[96][11][6] + xor_out[97][11][6] + xor_out[98][11][6] + xor_out[99][11][6];

assign sum_out[0][11][7] = xor_out[0][11][7] + xor_out[1][11][7] + xor_out[2][11][7] + xor_out[3][11][7] + xor_out[4][11][7];
assign sum_out[1][11][7] = xor_out[5][11][7] + xor_out[6][11][7] + xor_out[7][11][7] + xor_out[8][11][7] + xor_out[9][11][7];
assign sum_out[2][11][7] = xor_out[10][11][7] + xor_out[11][11][7] + xor_out[12][11][7] + xor_out[13][11][7] + xor_out[14][11][7];
assign sum_out[3][11][7] = xor_out[15][11][7] + xor_out[16][11][7] + xor_out[17][11][7] + xor_out[18][11][7] + xor_out[19][11][7];
assign sum_out[4][11][7] = xor_out[20][11][7] + xor_out[21][11][7] + xor_out[22][11][7] + xor_out[23][11][7] + xor_out[24][11][7];
assign sum_out[5][11][7] = xor_out[25][11][7] + xor_out[26][11][7] + xor_out[27][11][7] + xor_out[28][11][7] + xor_out[29][11][7];
assign sum_out[6][11][7] = xor_out[30][11][7] + xor_out[31][11][7] + xor_out[32][11][7] + xor_out[33][11][7] + xor_out[34][11][7];
assign sum_out[7][11][7] = xor_out[35][11][7] + xor_out[36][11][7] + xor_out[37][11][7] + xor_out[38][11][7] + xor_out[39][11][7];
assign sum_out[8][11][7] = xor_out[40][11][7] + xor_out[41][11][7] + xor_out[42][11][7] + xor_out[43][11][7] + xor_out[44][11][7];
assign sum_out[9][11][7] = xor_out[45][11][7] + xor_out[46][11][7] + xor_out[47][11][7] + xor_out[48][11][7] + xor_out[49][11][7];
assign sum_out[10][11][7] = xor_out[50][11][7] + xor_out[51][11][7] + xor_out[52][11][7] + xor_out[53][11][7] + xor_out[54][11][7];
assign sum_out[11][11][7] = xor_out[55][11][7] + xor_out[56][11][7] + xor_out[57][11][7] + xor_out[58][11][7] + xor_out[59][11][7];
assign sum_out[12][11][7] = xor_out[60][11][7] + xor_out[61][11][7] + xor_out[62][11][7] + xor_out[63][11][7] + xor_out[64][11][7];
assign sum_out[13][11][7] = xor_out[65][11][7] + xor_out[66][11][7] + xor_out[67][11][7] + xor_out[68][11][7] + xor_out[69][11][7];
assign sum_out[14][11][7] = xor_out[70][11][7] + xor_out[71][11][7] + xor_out[72][11][7] + xor_out[73][11][7] + xor_out[74][11][7];
assign sum_out[15][11][7] = xor_out[75][11][7] + xor_out[76][11][7] + xor_out[77][11][7] + xor_out[78][11][7] + xor_out[79][11][7];
assign sum_out[16][11][7] = xor_out[80][11][7] + xor_out[81][11][7] + xor_out[82][11][7] + xor_out[83][11][7] + xor_out[84][11][7];
assign sum_out[17][11][7] = xor_out[85][11][7] + xor_out[86][11][7] + xor_out[87][11][7] + xor_out[88][11][7] + xor_out[89][11][7];
assign sum_out[18][11][7] = xor_out[90][11][7] + xor_out[91][11][7] + xor_out[92][11][7] + xor_out[93][11][7] + xor_out[94][11][7];
assign sum_out[19][11][7] = xor_out[95][11][7] + xor_out[96][11][7] + xor_out[97][11][7] + xor_out[98][11][7] + xor_out[99][11][7];

assign sum_out[0][11][8] = xor_out[0][11][8] + xor_out[1][11][8] + xor_out[2][11][8] + xor_out[3][11][8] + xor_out[4][11][8];
assign sum_out[1][11][8] = xor_out[5][11][8] + xor_out[6][11][8] + xor_out[7][11][8] + xor_out[8][11][8] + xor_out[9][11][8];
assign sum_out[2][11][8] = xor_out[10][11][8] + xor_out[11][11][8] + xor_out[12][11][8] + xor_out[13][11][8] + xor_out[14][11][8];
assign sum_out[3][11][8] = xor_out[15][11][8] + xor_out[16][11][8] + xor_out[17][11][8] + xor_out[18][11][8] + xor_out[19][11][8];
assign sum_out[4][11][8] = xor_out[20][11][8] + xor_out[21][11][8] + xor_out[22][11][8] + xor_out[23][11][8] + xor_out[24][11][8];
assign sum_out[5][11][8] = xor_out[25][11][8] + xor_out[26][11][8] + xor_out[27][11][8] + xor_out[28][11][8] + xor_out[29][11][8];
assign sum_out[6][11][8] = xor_out[30][11][8] + xor_out[31][11][8] + xor_out[32][11][8] + xor_out[33][11][8] + xor_out[34][11][8];
assign sum_out[7][11][8] = xor_out[35][11][8] + xor_out[36][11][8] + xor_out[37][11][8] + xor_out[38][11][8] + xor_out[39][11][8];
assign sum_out[8][11][8] = xor_out[40][11][8] + xor_out[41][11][8] + xor_out[42][11][8] + xor_out[43][11][8] + xor_out[44][11][8];
assign sum_out[9][11][8] = xor_out[45][11][8] + xor_out[46][11][8] + xor_out[47][11][8] + xor_out[48][11][8] + xor_out[49][11][8];
assign sum_out[10][11][8] = xor_out[50][11][8] + xor_out[51][11][8] + xor_out[52][11][8] + xor_out[53][11][8] + xor_out[54][11][8];
assign sum_out[11][11][8] = xor_out[55][11][8] + xor_out[56][11][8] + xor_out[57][11][8] + xor_out[58][11][8] + xor_out[59][11][8];
assign sum_out[12][11][8] = xor_out[60][11][8] + xor_out[61][11][8] + xor_out[62][11][8] + xor_out[63][11][8] + xor_out[64][11][8];
assign sum_out[13][11][8] = xor_out[65][11][8] + xor_out[66][11][8] + xor_out[67][11][8] + xor_out[68][11][8] + xor_out[69][11][8];
assign sum_out[14][11][8] = xor_out[70][11][8] + xor_out[71][11][8] + xor_out[72][11][8] + xor_out[73][11][8] + xor_out[74][11][8];
assign sum_out[15][11][8] = xor_out[75][11][8] + xor_out[76][11][8] + xor_out[77][11][8] + xor_out[78][11][8] + xor_out[79][11][8];
assign sum_out[16][11][8] = xor_out[80][11][8] + xor_out[81][11][8] + xor_out[82][11][8] + xor_out[83][11][8] + xor_out[84][11][8];
assign sum_out[17][11][8] = xor_out[85][11][8] + xor_out[86][11][8] + xor_out[87][11][8] + xor_out[88][11][8] + xor_out[89][11][8];
assign sum_out[18][11][8] = xor_out[90][11][8] + xor_out[91][11][8] + xor_out[92][11][8] + xor_out[93][11][8] + xor_out[94][11][8];
assign sum_out[19][11][8] = xor_out[95][11][8] + xor_out[96][11][8] + xor_out[97][11][8] + xor_out[98][11][8] + xor_out[99][11][8];

assign sum_out[0][11][9] = xor_out[0][11][9] + xor_out[1][11][9] + xor_out[2][11][9] + xor_out[3][11][9] + xor_out[4][11][9];
assign sum_out[1][11][9] = xor_out[5][11][9] + xor_out[6][11][9] + xor_out[7][11][9] + xor_out[8][11][9] + xor_out[9][11][9];
assign sum_out[2][11][9] = xor_out[10][11][9] + xor_out[11][11][9] + xor_out[12][11][9] + xor_out[13][11][9] + xor_out[14][11][9];
assign sum_out[3][11][9] = xor_out[15][11][9] + xor_out[16][11][9] + xor_out[17][11][9] + xor_out[18][11][9] + xor_out[19][11][9];
assign sum_out[4][11][9] = xor_out[20][11][9] + xor_out[21][11][9] + xor_out[22][11][9] + xor_out[23][11][9] + xor_out[24][11][9];
assign sum_out[5][11][9] = xor_out[25][11][9] + xor_out[26][11][9] + xor_out[27][11][9] + xor_out[28][11][9] + xor_out[29][11][9];
assign sum_out[6][11][9] = xor_out[30][11][9] + xor_out[31][11][9] + xor_out[32][11][9] + xor_out[33][11][9] + xor_out[34][11][9];
assign sum_out[7][11][9] = xor_out[35][11][9] + xor_out[36][11][9] + xor_out[37][11][9] + xor_out[38][11][9] + xor_out[39][11][9];
assign sum_out[8][11][9] = xor_out[40][11][9] + xor_out[41][11][9] + xor_out[42][11][9] + xor_out[43][11][9] + xor_out[44][11][9];
assign sum_out[9][11][9] = xor_out[45][11][9] + xor_out[46][11][9] + xor_out[47][11][9] + xor_out[48][11][9] + xor_out[49][11][9];
assign sum_out[10][11][9] = xor_out[50][11][9] + xor_out[51][11][9] + xor_out[52][11][9] + xor_out[53][11][9] + xor_out[54][11][9];
assign sum_out[11][11][9] = xor_out[55][11][9] + xor_out[56][11][9] + xor_out[57][11][9] + xor_out[58][11][9] + xor_out[59][11][9];
assign sum_out[12][11][9] = xor_out[60][11][9] + xor_out[61][11][9] + xor_out[62][11][9] + xor_out[63][11][9] + xor_out[64][11][9];
assign sum_out[13][11][9] = xor_out[65][11][9] + xor_out[66][11][9] + xor_out[67][11][9] + xor_out[68][11][9] + xor_out[69][11][9];
assign sum_out[14][11][9] = xor_out[70][11][9] + xor_out[71][11][9] + xor_out[72][11][9] + xor_out[73][11][9] + xor_out[74][11][9];
assign sum_out[15][11][9] = xor_out[75][11][9] + xor_out[76][11][9] + xor_out[77][11][9] + xor_out[78][11][9] + xor_out[79][11][9];
assign sum_out[16][11][9] = xor_out[80][11][9] + xor_out[81][11][9] + xor_out[82][11][9] + xor_out[83][11][9] + xor_out[84][11][9];
assign sum_out[17][11][9] = xor_out[85][11][9] + xor_out[86][11][9] + xor_out[87][11][9] + xor_out[88][11][9] + xor_out[89][11][9];
assign sum_out[18][11][9] = xor_out[90][11][9] + xor_out[91][11][9] + xor_out[92][11][9] + xor_out[93][11][9] + xor_out[94][11][9];
assign sum_out[19][11][9] = xor_out[95][11][9] + xor_out[96][11][9] + xor_out[97][11][9] + xor_out[98][11][9] + xor_out[99][11][9];

assign sum_out[0][11][10] = xor_out[0][11][10] + xor_out[1][11][10] + xor_out[2][11][10] + xor_out[3][11][10] + xor_out[4][11][10];
assign sum_out[1][11][10] = xor_out[5][11][10] + xor_out[6][11][10] + xor_out[7][11][10] + xor_out[8][11][10] + xor_out[9][11][10];
assign sum_out[2][11][10] = xor_out[10][11][10] + xor_out[11][11][10] + xor_out[12][11][10] + xor_out[13][11][10] + xor_out[14][11][10];
assign sum_out[3][11][10] = xor_out[15][11][10] + xor_out[16][11][10] + xor_out[17][11][10] + xor_out[18][11][10] + xor_out[19][11][10];
assign sum_out[4][11][10] = xor_out[20][11][10] + xor_out[21][11][10] + xor_out[22][11][10] + xor_out[23][11][10] + xor_out[24][11][10];
assign sum_out[5][11][10] = xor_out[25][11][10] + xor_out[26][11][10] + xor_out[27][11][10] + xor_out[28][11][10] + xor_out[29][11][10];
assign sum_out[6][11][10] = xor_out[30][11][10] + xor_out[31][11][10] + xor_out[32][11][10] + xor_out[33][11][10] + xor_out[34][11][10];
assign sum_out[7][11][10] = xor_out[35][11][10] + xor_out[36][11][10] + xor_out[37][11][10] + xor_out[38][11][10] + xor_out[39][11][10];
assign sum_out[8][11][10] = xor_out[40][11][10] + xor_out[41][11][10] + xor_out[42][11][10] + xor_out[43][11][10] + xor_out[44][11][10];
assign sum_out[9][11][10] = xor_out[45][11][10] + xor_out[46][11][10] + xor_out[47][11][10] + xor_out[48][11][10] + xor_out[49][11][10];
assign sum_out[10][11][10] = xor_out[50][11][10] + xor_out[51][11][10] + xor_out[52][11][10] + xor_out[53][11][10] + xor_out[54][11][10];
assign sum_out[11][11][10] = xor_out[55][11][10] + xor_out[56][11][10] + xor_out[57][11][10] + xor_out[58][11][10] + xor_out[59][11][10];
assign sum_out[12][11][10] = xor_out[60][11][10] + xor_out[61][11][10] + xor_out[62][11][10] + xor_out[63][11][10] + xor_out[64][11][10];
assign sum_out[13][11][10] = xor_out[65][11][10] + xor_out[66][11][10] + xor_out[67][11][10] + xor_out[68][11][10] + xor_out[69][11][10];
assign sum_out[14][11][10] = xor_out[70][11][10] + xor_out[71][11][10] + xor_out[72][11][10] + xor_out[73][11][10] + xor_out[74][11][10];
assign sum_out[15][11][10] = xor_out[75][11][10] + xor_out[76][11][10] + xor_out[77][11][10] + xor_out[78][11][10] + xor_out[79][11][10];
assign sum_out[16][11][10] = xor_out[80][11][10] + xor_out[81][11][10] + xor_out[82][11][10] + xor_out[83][11][10] + xor_out[84][11][10];
assign sum_out[17][11][10] = xor_out[85][11][10] + xor_out[86][11][10] + xor_out[87][11][10] + xor_out[88][11][10] + xor_out[89][11][10];
assign sum_out[18][11][10] = xor_out[90][11][10] + xor_out[91][11][10] + xor_out[92][11][10] + xor_out[93][11][10] + xor_out[94][11][10];
assign sum_out[19][11][10] = xor_out[95][11][10] + xor_out[96][11][10] + xor_out[97][11][10] + xor_out[98][11][10] + xor_out[99][11][10];

assign sum_out[0][11][11] = xor_out[0][11][11] + xor_out[1][11][11] + xor_out[2][11][11] + xor_out[3][11][11] + xor_out[4][11][11];
assign sum_out[1][11][11] = xor_out[5][11][11] + xor_out[6][11][11] + xor_out[7][11][11] + xor_out[8][11][11] + xor_out[9][11][11];
assign sum_out[2][11][11] = xor_out[10][11][11] + xor_out[11][11][11] + xor_out[12][11][11] + xor_out[13][11][11] + xor_out[14][11][11];
assign sum_out[3][11][11] = xor_out[15][11][11] + xor_out[16][11][11] + xor_out[17][11][11] + xor_out[18][11][11] + xor_out[19][11][11];
assign sum_out[4][11][11] = xor_out[20][11][11] + xor_out[21][11][11] + xor_out[22][11][11] + xor_out[23][11][11] + xor_out[24][11][11];
assign sum_out[5][11][11] = xor_out[25][11][11] + xor_out[26][11][11] + xor_out[27][11][11] + xor_out[28][11][11] + xor_out[29][11][11];
assign sum_out[6][11][11] = xor_out[30][11][11] + xor_out[31][11][11] + xor_out[32][11][11] + xor_out[33][11][11] + xor_out[34][11][11];
assign sum_out[7][11][11] = xor_out[35][11][11] + xor_out[36][11][11] + xor_out[37][11][11] + xor_out[38][11][11] + xor_out[39][11][11];
assign sum_out[8][11][11] = xor_out[40][11][11] + xor_out[41][11][11] + xor_out[42][11][11] + xor_out[43][11][11] + xor_out[44][11][11];
assign sum_out[9][11][11] = xor_out[45][11][11] + xor_out[46][11][11] + xor_out[47][11][11] + xor_out[48][11][11] + xor_out[49][11][11];
assign sum_out[10][11][11] = xor_out[50][11][11] + xor_out[51][11][11] + xor_out[52][11][11] + xor_out[53][11][11] + xor_out[54][11][11];
assign sum_out[11][11][11] = xor_out[55][11][11] + xor_out[56][11][11] + xor_out[57][11][11] + xor_out[58][11][11] + xor_out[59][11][11];
assign sum_out[12][11][11] = xor_out[60][11][11] + xor_out[61][11][11] + xor_out[62][11][11] + xor_out[63][11][11] + xor_out[64][11][11];
assign sum_out[13][11][11] = xor_out[65][11][11] + xor_out[66][11][11] + xor_out[67][11][11] + xor_out[68][11][11] + xor_out[69][11][11];
assign sum_out[14][11][11] = xor_out[70][11][11] + xor_out[71][11][11] + xor_out[72][11][11] + xor_out[73][11][11] + xor_out[74][11][11];
assign sum_out[15][11][11] = xor_out[75][11][11] + xor_out[76][11][11] + xor_out[77][11][11] + xor_out[78][11][11] + xor_out[79][11][11];
assign sum_out[16][11][11] = xor_out[80][11][11] + xor_out[81][11][11] + xor_out[82][11][11] + xor_out[83][11][11] + xor_out[84][11][11];
assign sum_out[17][11][11] = xor_out[85][11][11] + xor_out[86][11][11] + xor_out[87][11][11] + xor_out[88][11][11] + xor_out[89][11][11];
assign sum_out[18][11][11] = xor_out[90][11][11] + xor_out[91][11][11] + xor_out[92][11][11] + xor_out[93][11][11] + xor_out[94][11][11];
assign sum_out[19][11][11] = xor_out[95][11][11] + xor_out[96][11][11] + xor_out[97][11][11] + xor_out[98][11][11] + xor_out[99][11][11];

assign sum_out[0][11][12] = xor_out[0][11][12] + xor_out[1][11][12] + xor_out[2][11][12] + xor_out[3][11][12] + xor_out[4][11][12];
assign sum_out[1][11][12] = xor_out[5][11][12] + xor_out[6][11][12] + xor_out[7][11][12] + xor_out[8][11][12] + xor_out[9][11][12];
assign sum_out[2][11][12] = xor_out[10][11][12] + xor_out[11][11][12] + xor_out[12][11][12] + xor_out[13][11][12] + xor_out[14][11][12];
assign sum_out[3][11][12] = xor_out[15][11][12] + xor_out[16][11][12] + xor_out[17][11][12] + xor_out[18][11][12] + xor_out[19][11][12];
assign sum_out[4][11][12] = xor_out[20][11][12] + xor_out[21][11][12] + xor_out[22][11][12] + xor_out[23][11][12] + xor_out[24][11][12];
assign sum_out[5][11][12] = xor_out[25][11][12] + xor_out[26][11][12] + xor_out[27][11][12] + xor_out[28][11][12] + xor_out[29][11][12];
assign sum_out[6][11][12] = xor_out[30][11][12] + xor_out[31][11][12] + xor_out[32][11][12] + xor_out[33][11][12] + xor_out[34][11][12];
assign sum_out[7][11][12] = xor_out[35][11][12] + xor_out[36][11][12] + xor_out[37][11][12] + xor_out[38][11][12] + xor_out[39][11][12];
assign sum_out[8][11][12] = xor_out[40][11][12] + xor_out[41][11][12] + xor_out[42][11][12] + xor_out[43][11][12] + xor_out[44][11][12];
assign sum_out[9][11][12] = xor_out[45][11][12] + xor_out[46][11][12] + xor_out[47][11][12] + xor_out[48][11][12] + xor_out[49][11][12];
assign sum_out[10][11][12] = xor_out[50][11][12] + xor_out[51][11][12] + xor_out[52][11][12] + xor_out[53][11][12] + xor_out[54][11][12];
assign sum_out[11][11][12] = xor_out[55][11][12] + xor_out[56][11][12] + xor_out[57][11][12] + xor_out[58][11][12] + xor_out[59][11][12];
assign sum_out[12][11][12] = xor_out[60][11][12] + xor_out[61][11][12] + xor_out[62][11][12] + xor_out[63][11][12] + xor_out[64][11][12];
assign sum_out[13][11][12] = xor_out[65][11][12] + xor_out[66][11][12] + xor_out[67][11][12] + xor_out[68][11][12] + xor_out[69][11][12];
assign sum_out[14][11][12] = xor_out[70][11][12] + xor_out[71][11][12] + xor_out[72][11][12] + xor_out[73][11][12] + xor_out[74][11][12];
assign sum_out[15][11][12] = xor_out[75][11][12] + xor_out[76][11][12] + xor_out[77][11][12] + xor_out[78][11][12] + xor_out[79][11][12];
assign sum_out[16][11][12] = xor_out[80][11][12] + xor_out[81][11][12] + xor_out[82][11][12] + xor_out[83][11][12] + xor_out[84][11][12];
assign sum_out[17][11][12] = xor_out[85][11][12] + xor_out[86][11][12] + xor_out[87][11][12] + xor_out[88][11][12] + xor_out[89][11][12];
assign sum_out[18][11][12] = xor_out[90][11][12] + xor_out[91][11][12] + xor_out[92][11][12] + xor_out[93][11][12] + xor_out[94][11][12];
assign sum_out[19][11][12] = xor_out[95][11][12] + xor_out[96][11][12] + xor_out[97][11][12] + xor_out[98][11][12] + xor_out[99][11][12];

assign sum_out[0][11][13] = xor_out[0][11][13] + xor_out[1][11][13] + xor_out[2][11][13] + xor_out[3][11][13] + xor_out[4][11][13];
assign sum_out[1][11][13] = xor_out[5][11][13] + xor_out[6][11][13] + xor_out[7][11][13] + xor_out[8][11][13] + xor_out[9][11][13];
assign sum_out[2][11][13] = xor_out[10][11][13] + xor_out[11][11][13] + xor_out[12][11][13] + xor_out[13][11][13] + xor_out[14][11][13];
assign sum_out[3][11][13] = xor_out[15][11][13] + xor_out[16][11][13] + xor_out[17][11][13] + xor_out[18][11][13] + xor_out[19][11][13];
assign sum_out[4][11][13] = xor_out[20][11][13] + xor_out[21][11][13] + xor_out[22][11][13] + xor_out[23][11][13] + xor_out[24][11][13];
assign sum_out[5][11][13] = xor_out[25][11][13] + xor_out[26][11][13] + xor_out[27][11][13] + xor_out[28][11][13] + xor_out[29][11][13];
assign sum_out[6][11][13] = xor_out[30][11][13] + xor_out[31][11][13] + xor_out[32][11][13] + xor_out[33][11][13] + xor_out[34][11][13];
assign sum_out[7][11][13] = xor_out[35][11][13] + xor_out[36][11][13] + xor_out[37][11][13] + xor_out[38][11][13] + xor_out[39][11][13];
assign sum_out[8][11][13] = xor_out[40][11][13] + xor_out[41][11][13] + xor_out[42][11][13] + xor_out[43][11][13] + xor_out[44][11][13];
assign sum_out[9][11][13] = xor_out[45][11][13] + xor_out[46][11][13] + xor_out[47][11][13] + xor_out[48][11][13] + xor_out[49][11][13];
assign sum_out[10][11][13] = xor_out[50][11][13] + xor_out[51][11][13] + xor_out[52][11][13] + xor_out[53][11][13] + xor_out[54][11][13];
assign sum_out[11][11][13] = xor_out[55][11][13] + xor_out[56][11][13] + xor_out[57][11][13] + xor_out[58][11][13] + xor_out[59][11][13];
assign sum_out[12][11][13] = xor_out[60][11][13] + xor_out[61][11][13] + xor_out[62][11][13] + xor_out[63][11][13] + xor_out[64][11][13];
assign sum_out[13][11][13] = xor_out[65][11][13] + xor_out[66][11][13] + xor_out[67][11][13] + xor_out[68][11][13] + xor_out[69][11][13];
assign sum_out[14][11][13] = xor_out[70][11][13] + xor_out[71][11][13] + xor_out[72][11][13] + xor_out[73][11][13] + xor_out[74][11][13];
assign sum_out[15][11][13] = xor_out[75][11][13] + xor_out[76][11][13] + xor_out[77][11][13] + xor_out[78][11][13] + xor_out[79][11][13];
assign sum_out[16][11][13] = xor_out[80][11][13] + xor_out[81][11][13] + xor_out[82][11][13] + xor_out[83][11][13] + xor_out[84][11][13];
assign sum_out[17][11][13] = xor_out[85][11][13] + xor_out[86][11][13] + xor_out[87][11][13] + xor_out[88][11][13] + xor_out[89][11][13];
assign sum_out[18][11][13] = xor_out[90][11][13] + xor_out[91][11][13] + xor_out[92][11][13] + xor_out[93][11][13] + xor_out[94][11][13];
assign sum_out[19][11][13] = xor_out[95][11][13] + xor_out[96][11][13] + xor_out[97][11][13] + xor_out[98][11][13] + xor_out[99][11][13];

assign sum_out[0][11][14] = xor_out[0][11][14] + xor_out[1][11][14] + xor_out[2][11][14] + xor_out[3][11][14] + xor_out[4][11][14];
assign sum_out[1][11][14] = xor_out[5][11][14] + xor_out[6][11][14] + xor_out[7][11][14] + xor_out[8][11][14] + xor_out[9][11][14];
assign sum_out[2][11][14] = xor_out[10][11][14] + xor_out[11][11][14] + xor_out[12][11][14] + xor_out[13][11][14] + xor_out[14][11][14];
assign sum_out[3][11][14] = xor_out[15][11][14] + xor_out[16][11][14] + xor_out[17][11][14] + xor_out[18][11][14] + xor_out[19][11][14];
assign sum_out[4][11][14] = xor_out[20][11][14] + xor_out[21][11][14] + xor_out[22][11][14] + xor_out[23][11][14] + xor_out[24][11][14];
assign sum_out[5][11][14] = xor_out[25][11][14] + xor_out[26][11][14] + xor_out[27][11][14] + xor_out[28][11][14] + xor_out[29][11][14];
assign sum_out[6][11][14] = xor_out[30][11][14] + xor_out[31][11][14] + xor_out[32][11][14] + xor_out[33][11][14] + xor_out[34][11][14];
assign sum_out[7][11][14] = xor_out[35][11][14] + xor_out[36][11][14] + xor_out[37][11][14] + xor_out[38][11][14] + xor_out[39][11][14];
assign sum_out[8][11][14] = xor_out[40][11][14] + xor_out[41][11][14] + xor_out[42][11][14] + xor_out[43][11][14] + xor_out[44][11][14];
assign sum_out[9][11][14] = xor_out[45][11][14] + xor_out[46][11][14] + xor_out[47][11][14] + xor_out[48][11][14] + xor_out[49][11][14];
assign sum_out[10][11][14] = xor_out[50][11][14] + xor_out[51][11][14] + xor_out[52][11][14] + xor_out[53][11][14] + xor_out[54][11][14];
assign sum_out[11][11][14] = xor_out[55][11][14] + xor_out[56][11][14] + xor_out[57][11][14] + xor_out[58][11][14] + xor_out[59][11][14];
assign sum_out[12][11][14] = xor_out[60][11][14] + xor_out[61][11][14] + xor_out[62][11][14] + xor_out[63][11][14] + xor_out[64][11][14];
assign sum_out[13][11][14] = xor_out[65][11][14] + xor_out[66][11][14] + xor_out[67][11][14] + xor_out[68][11][14] + xor_out[69][11][14];
assign sum_out[14][11][14] = xor_out[70][11][14] + xor_out[71][11][14] + xor_out[72][11][14] + xor_out[73][11][14] + xor_out[74][11][14];
assign sum_out[15][11][14] = xor_out[75][11][14] + xor_out[76][11][14] + xor_out[77][11][14] + xor_out[78][11][14] + xor_out[79][11][14];
assign sum_out[16][11][14] = xor_out[80][11][14] + xor_out[81][11][14] + xor_out[82][11][14] + xor_out[83][11][14] + xor_out[84][11][14];
assign sum_out[17][11][14] = xor_out[85][11][14] + xor_out[86][11][14] + xor_out[87][11][14] + xor_out[88][11][14] + xor_out[89][11][14];
assign sum_out[18][11][14] = xor_out[90][11][14] + xor_out[91][11][14] + xor_out[92][11][14] + xor_out[93][11][14] + xor_out[94][11][14];
assign sum_out[19][11][14] = xor_out[95][11][14] + xor_out[96][11][14] + xor_out[97][11][14] + xor_out[98][11][14] + xor_out[99][11][14];

assign sum_out[0][11][15] = xor_out[0][11][15] + xor_out[1][11][15] + xor_out[2][11][15] + xor_out[3][11][15] + xor_out[4][11][15];
assign sum_out[1][11][15] = xor_out[5][11][15] + xor_out[6][11][15] + xor_out[7][11][15] + xor_out[8][11][15] + xor_out[9][11][15];
assign sum_out[2][11][15] = xor_out[10][11][15] + xor_out[11][11][15] + xor_out[12][11][15] + xor_out[13][11][15] + xor_out[14][11][15];
assign sum_out[3][11][15] = xor_out[15][11][15] + xor_out[16][11][15] + xor_out[17][11][15] + xor_out[18][11][15] + xor_out[19][11][15];
assign sum_out[4][11][15] = xor_out[20][11][15] + xor_out[21][11][15] + xor_out[22][11][15] + xor_out[23][11][15] + xor_out[24][11][15];
assign sum_out[5][11][15] = xor_out[25][11][15] + xor_out[26][11][15] + xor_out[27][11][15] + xor_out[28][11][15] + xor_out[29][11][15];
assign sum_out[6][11][15] = xor_out[30][11][15] + xor_out[31][11][15] + xor_out[32][11][15] + xor_out[33][11][15] + xor_out[34][11][15];
assign sum_out[7][11][15] = xor_out[35][11][15] + xor_out[36][11][15] + xor_out[37][11][15] + xor_out[38][11][15] + xor_out[39][11][15];
assign sum_out[8][11][15] = xor_out[40][11][15] + xor_out[41][11][15] + xor_out[42][11][15] + xor_out[43][11][15] + xor_out[44][11][15];
assign sum_out[9][11][15] = xor_out[45][11][15] + xor_out[46][11][15] + xor_out[47][11][15] + xor_out[48][11][15] + xor_out[49][11][15];
assign sum_out[10][11][15] = xor_out[50][11][15] + xor_out[51][11][15] + xor_out[52][11][15] + xor_out[53][11][15] + xor_out[54][11][15];
assign sum_out[11][11][15] = xor_out[55][11][15] + xor_out[56][11][15] + xor_out[57][11][15] + xor_out[58][11][15] + xor_out[59][11][15];
assign sum_out[12][11][15] = xor_out[60][11][15] + xor_out[61][11][15] + xor_out[62][11][15] + xor_out[63][11][15] + xor_out[64][11][15];
assign sum_out[13][11][15] = xor_out[65][11][15] + xor_out[66][11][15] + xor_out[67][11][15] + xor_out[68][11][15] + xor_out[69][11][15];
assign sum_out[14][11][15] = xor_out[70][11][15] + xor_out[71][11][15] + xor_out[72][11][15] + xor_out[73][11][15] + xor_out[74][11][15];
assign sum_out[15][11][15] = xor_out[75][11][15] + xor_out[76][11][15] + xor_out[77][11][15] + xor_out[78][11][15] + xor_out[79][11][15];
assign sum_out[16][11][15] = xor_out[80][11][15] + xor_out[81][11][15] + xor_out[82][11][15] + xor_out[83][11][15] + xor_out[84][11][15];
assign sum_out[17][11][15] = xor_out[85][11][15] + xor_out[86][11][15] + xor_out[87][11][15] + xor_out[88][11][15] + xor_out[89][11][15];
assign sum_out[18][11][15] = xor_out[90][11][15] + xor_out[91][11][15] + xor_out[92][11][15] + xor_out[93][11][15] + xor_out[94][11][15];
assign sum_out[19][11][15] = xor_out[95][11][15] + xor_out[96][11][15] + xor_out[97][11][15] + xor_out[98][11][15] + xor_out[99][11][15];

assign sum_out[0][11][16] = xor_out[0][11][16] + xor_out[1][11][16] + xor_out[2][11][16] + xor_out[3][11][16] + xor_out[4][11][16];
assign sum_out[1][11][16] = xor_out[5][11][16] + xor_out[6][11][16] + xor_out[7][11][16] + xor_out[8][11][16] + xor_out[9][11][16];
assign sum_out[2][11][16] = xor_out[10][11][16] + xor_out[11][11][16] + xor_out[12][11][16] + xor_out[13][11][16] + xor_out[14][11][16];
assign sum_out[3][11][16] = xor_out[15][11][16] + xor_out[16][11][16] + xor_out[17][11][16] + xor_out[18][11][16] + xor_out[19][11][16];
assign sum_out[4][11][16] = xor_out[20][11][16] + xor_out[21][11][16] + xor_out[22][11][16] + xor_out[23][11][16] + xor_out[24][11][16];
assign sum_out[5][11][16] = xor_out[25][11][16] + xor_out[26][11][16] + xor_out[27][11][16] + xor_out[28][11][16] + xor_out[29][11][16];
assign sum_out[6][11][16] = xor_out[30][11][16] + xor_out[31][11][16] + xor_out[32][11][16] + xor_out[33][11][16] + xor_out[34][11][16];
assign sum_out[7][11][16] = xor_out[35][11][16] + xor_out[36][11][16] + xor_out[37][11][16] + xor_out[38][11][16] + xor_out[39][11][16];
assign sum_out[8][11][16] = xor_out[40][11][16] + xor_out[41][11][16] + xor_out[42][11][16] + xor_out[43][11][16] + xor_out[44][11][16];
assign sum_out[9][11][16] = xor_out[45][11][16] + xor_out[46][11][16] + xor_out[47][11][16] + xor_out[48][11][16] + xor_out[49][11][16];
assign sum_out[10][11][16] = xor_out[50][11][16] + xor_out[51][11][16] + xor_out[52][11][16] + xor_out[53][11][16] + xor_out[54][11][16];
assign sum_out[11][11][16] = xor_out[55][11][16] + xor_out[56][11][16] + xor_out[57][11][16] + xor_out[58][11][16] + xor_out[59][11][16];
assign sum_out[12][11][16] = xor_out[60][11][16] + xor_out[61][11][16] + xor_out[62][11][16] + xor_out[63][11][16] + xor_out[64][11][16];
assign sum_out[13][11][16] = xor_out[65][11][16] + xor_out[66][11][16] + xor_out[67][11][16] + xor_out[68][11][16] + xor_out[69][11][16];
assign sum_out[14][11][16] = xor_out[70][11][16] + xor_out[71][11][16] + xor_out[72][11][16] + xor_out[73][11][16] + xor_out[74][11][16];
assign sum_out[15][11][16] = xor_out[75][11][16] + xor_out[76][11][16] + xor_out[77][11][16] + xor_out[78][11][16] + xor_out[79][11][16];
assign sum_out[16][11][16] = xor_out[80][11][16] + xor_out[81][11][16] + xor_out[82][11][16] + xor_out[83][11][16] + xor_out[84][11][16];
assign sum_out[17][11][16] = xor_out[85][11][16] + xor_out[86][11][16] + xor_out[87][11][16] + xor_out[88][11][16] + xor_out[89][11][16];
assign sum_out[18][11][16] = xor_out[90][11][16] + xor_out[91][11][16] + xor_out[92][11][16] + xor_out[93][11][16] + xor_out[94][11][16];
assign sum_out[19][11][16] = xor_out[95][11][16] + xor_out[96][11][16] + xor_out[97][11][16] + xor_out[98][11][16] + xor_out[99][11][16];

assign sum_out[0][11][17] = xor_out[0][11][17] + xor_out[1][11][17] + xor_out[2][11][17] + xor_out[3][11][17] + xor_out[4][11][17];
assign sum_out[1][11][17] = xor_out[5][11][17] + xor_out[6][11][17] + xor_out[7][11][17] + xor_out[8][11][17] + xor_out[9][11][17];
assign sum_out[2][11][17] = xor_out[10][11][17] + xor_out[11][11][17] + xor_out[12][11][17] + xor_out[13][11][17] + xor_out[14][11][17];
assign sum_out[3][11][17] = xor_out[15][11][17] + xor_out[16][11][17] + xor_out[17][11][17] + xor_out[18][11][17] + xor_out[19][11][17];
assign sum_out[4][11][17] = xor_out[20][11][17] + xor_out[21][11][17] + xor_out[22][11][17] + xor_out[23][11][17] + xor_out[24][11][17];
assign sum_out[5][11][17] = xor_out[25][11][17] + xor_out[26][11][17] + xor_out[27][11][17] + xor_out[28][11][17] + xor_out[29][11][17];
assign sum_out[6][11][17] = xor_out[30][11][17] + xor_out[31][11][17] + xor_out[32][11][17] + xor_out[33][11][17] + xor_out[34][11][17];
assign sum_out[7][11][17] = xor_out[35][11][17] + xor_out[36][11][17] + xor_out[37][11][17] + xor_out[38][11][17] + xor_out[39][11][17];
assign sum_out[8][11][17] = xor_out[40][11][17] + xor_out[41][11][17] + xor_out[42][11][17] + xor_out[43][11][17] + xor_out[44][11][17];
assign sum_out[9][11][17] = xor_out[45][11][17] + xor_out[46][11][17] + xor_out[47][11][17] + xor_out[48][11][17] + xor_out[49][11][17];
assign sum_out[10][11][17] = xor_out[50][11][17] + xor_out[51][11][17] + xor_out[52][11][17] + xor_out[53][11][17] + xor_out[54][11][17];
assign sum_out[11][11][17] = xor_out[55][11][17] + xor_out[56][11][17] + xor_out[57][11][17] + xor_out[58][11][17] + xor_out[59][11][17];
assign sum_out[12][11][17] = xor_out[60][11][17] + xor_out[61][11][17] + xor_out[62][11][17] + xor_out[63][11][17] + xor_out[64][11][17];
assign sum_out[13][11][17] = xor_out[65][11][17] + xor_out[66][11][17] + xor_out[67][11][17] + xor_out[68][11][17] + xor_out[69][11][17];
assign sum_out[14][11][17] = xor_out[70][11][17] + xor_out[71][11][17] + xor_out[72][11][17] + xor_out[73][11][17] + xor_out[74][11][17];
assign sum_out[15][11][17] = xor_out[75][11][17] + xor_out[76][11][17] + xor_out[77][11][17] + xor_out[78][11][17] + xor_out[79][11][17];
assign sum_out[16][11][17] = xor_out[80][11][17] + xor_out[81][11][17] + xor_out[82][11][17] + xor_out[83][11][17] + xor_out[84][11][17];
assign sum_out[17][11][17] = xor_out[85][11][17] + xor_out[86][11][17] + xor_out[87][11][17] + xor_out[88][11][17] + xor_out[89][11][17];
assign sum_out[18][11][17] = xor_out[90][11][17] + xor_out[91][11][17] + xor_out[92][11][17] + xor_out[93][11][17] + xor_out[94][11][17];
assign sum_out[19][11][17] = xor_out[95][11][17] + xor_out[96][11][17] + xor_out[97][11][17] + xor_out[98][11][17] + xor_out[99][11][17];

assign sum_out[0][11][18] = xor_out[0][11][18] + xor_out[1][11][18] + xor_out[2][11][18] + xor_out[3][11][18] + xor_out[4][11][18];
assign sum_out[1][11][18] = xor_out[5][11][18] + xor_out[6][11][18] + xor_out[7][11][18] + xor_out[8][11][18] + xor_out[9][11][18];
assign sum_out[2][11][18] = xor_out[10][11][18] + xor_out[11][11][18] + xor_out[12][11][18] + xor_out[13][11][18] + xor_out[14][11][18];
assign sum_out[3][11][18] = xor_out[15][11][18] + xor_out[16][11][18] + xor_out[17][11][18] + xor_out[18][11][18] + xor_out[19][11][18];
assign sum_out[4][11][18] = xor_out[20][11][18] + xor_out[21][11][18] + xor_out[22][11][18] + xor_out[23][11][18] + xor_out[24][11][18];
assign sum_out[5][11][18] = xor_out[25][11][18] + xor_out[26][11][18] + xor_out[27][11][18] + xor_out[28][11][18] + xor_out[29][11][18];
assign sum_out[6][11][18] = xor_out[30][11][18] + xor_out[31][11][18] + xor_out[32][11][18] + xor_out[33][11][18] + xor_out[34][11][18];
assign sum_out[7][11][18] = xor_out[35][11][18] + xor_out[36][11][18] + xor_out[37][11][18] + xor_out[38][11][18] + xor_out[39][11][18];
assign sum_out[8][11][18] = xor_out[40][11][18] + xor_out[41][11][18] + xor_out[42][11][18] + xor_out[43][11][18] + xor_out[44][11][18];
assign sum_out[9][11][18] = xor_out[45][11][18] + xor_out[46][11][18] + xor_out[47][11][18] + xor_out[48][11][18] + xor_out[49][11][18];
assign sum_out[10][11][18] = xor_out[50][11][18] + xor_out[51][11][18] + xor_out[52][11][18] + xor_out[53][11][18] + xor_out[54][11][18];
assign sum_out[11][11][18] = xor_out[55][11][18] + xor_out[56][11][18] + xor_out[57][11][18] + xor_out[58][11][18] + xor_out[59][11][18];
assign sum_out[12][11][18] = xor_out[60][11][18] + xor_out[61][11][18] + xor_out[62][11][18] + xor_out[63][11][18] + xor_out[64][11][18];
assign sum_out[13][11][18] = xor_out[65][11][18] + xor_out[66][11][18] + xor_out[67][11][18] + xor_out[68][11][18] + xor_out[69][11][18];
assign sum_out[14][11][18] = xor_out[70][11][18] + xor_out[71][11][18] + xor_out[72][11][18] + xor_out[73][11][18] + xor_out[74][11][18];
assign sum_out[15][11][18] = xor_out[75][11][18] + xor_out[76][11][18] + xor_out[77][11][18] + xor_out[78][11][18] + xor_out[79][11][18];
assign sum_out[16][11][18] = xor_out[80][11][18] + xor_out[81][11][18] + xor_out[82][11][18] + xor_out[83][11][18] + xor_out[84][11][18];
assign sum_out[17][11][18] = xor_out[85][11][18] + xor_out[86][11][18] + xor_out[87][11][18] + xor_out[88][11][18] + xor_out[89][11][18];
assign sum_out[18][11][18] = xor_out[90][11][18] + xor_out[91][11][18] + xor_out[92][11][18] + xor_out[93][11][18] + xor_out[94][11][18];
assign sum_out[19][11][18] = xor_out[95][11][18] + xor_out[96][11][18] + xor_out[97][11][18] + xor_out[98][11][18] + xor_out[99][11][18];

assign sum_out[0][11][19] = xor_out[0][11][19] + xor_out[1][11][19] + xor_out[2][11][19] + xor_out[3][11][19] + xor_out[4][11][19];
assign sum_out[1][11][19] = xor_out[5][11][19] + xor_out[6][11][19] + xor_out[7][11][19] + xor_out[8][11][19] + xor_out[9][11][19];
assign sum_out[2][11][19] = xor_out[10][11][19] + xor_out[11][11][19] + xor_out[12][11][19] + xor_out[13][11][19] + xor_out[14][11][19];
assign sum_out[3][11][19] = xor_out[15][11][19] + xor_out[16][11][19] + xor_out[17][11][19] + xor_out[18][11][19] + xor_out[19][11][19];
assign sum_out[4][11][19] = xor_out[20][11][19] + xor_out[21][11][19] + xor_out[22][11][19] + xor_out[23][11][19] + xor_out[24][11][19];
assign sum_out[5][11][19] = xor_out[25][11][19] + xor_out[26][11][19] + xor_out[27][11][19] + xor_out[28][11][19] + xor_out[29][11][19];
assign sum_out[6][11][19] = xor_out[30][11][19] + xor_out[31][11][19] + xor_out[32][11][19] + xor_out[33][11][19] + xor_out[34][11][19];
assign sum_out[7][11][19] = xor_out[35][11][19] + xor_out[36][11][19] + xor_out[37][11][19] + xor_out[38][11][19] + xor_out[39][11][19];
assign sum_out[8][11][19] = xor_out[40][11][19] + xor_out[41][11][19] + xor_out[42][11][19] + xor_out[43][11][19] + xor_out[44][11][19];
assign sum_out[9][11][19] = xor_out[45][11][19] + xor_out[46][11][19] + xor_out[47][11][19] + xor_out[48][11][19] + xor_out[49][11][19];
assign sum_out[10][11][19] = xor_out[50][11][19] + xor_out[51][11][19] + xor_out[52][11][19] + xor_out[53][11][19] + xor_out[54][11][19];
assign sum_out[11][11][19] = xor_out[55][11][19] + xor_out[56][11][19] + xor_out[57][11][19] + xor_out[58][11][19] + xor_out[59][11][19];
assign sum_out[12][11][19] = xor_out[60][11][19] + xor_out[61][11][19] + xor_out[62][11][19] + xor_out[63][11][19] + xor_out[64][11][19];
assign sum_out[13][11][19] = xor_out[65][11][19] + xor_out[66][11][19] + xor_out[67][11][19] + xor_out[68][11][19] + xor_out[69][11][19];
assign sum_out[14][11][19] = xor_out[70][11][19] + xor_out[71][11][19] + xor_out[72][11][19] + xor_out[73][11][19] + xor_out[74][11][19];
assign sum_out[15][11][19] = xor_out[75][11][19] + xor_out[76][11][19] + xor_out[77][11][19] + xor_out[78][11][19] + xor_out[79][11][19];
assign sum_out[16][11][19] = xor_out[80][11][19] + xor_out[81][11][19] + xor_out[82][11][19] + xor_out[83][11][19] + xor_out[84][11][19];
assign sum_out[17][11][19] = xor_out[85][11][19] + xor_out[86][11][19] + xor_out[87][11][19] + xor_out[88][11][19] + xor_out[89][11][19];
assign sum_out[18][11][19] = xor_out[90][11][19] + xor_out[91][11][19] + xor_out[92][11][19] + xor_out[93][11][19] + xor_out[94][11][19];
assign sum_out[19][11][19] = xor_out[95][11][19] + xor_out[96][11][19] + xor_out[97][11][19] + xor_out[98][11][19] + xor_out[99][11][19];

assign sum_out[0][11][20] = xor_out[0][11][20] + xor_out[1][11][20] + xor_out[2][11][20] + xor_out[3][11][20] + xor_out[4][11][20];
assign sum_out[1][11][20] = xor_out[5][11][20] + xor_out[6][11][20] + xor_out[7][11][20] + xor_out[8][11][20] + xor_out[9][11][20];
assign sum_out[2][11][20] = xor_out[10][11][20] + xor_out[11][11][20] + xor_out[12][11][20] + xor_out[13][11][20] + xor_out[14][11][20];
assign sum_out[3][11][20] = xor_out[15][11][20] + xor_out[16][11][20] + xor_out[17][11][20] + xor_out[18][11][20] + xor_out[19][11][20];
assign sum_out[4][11][20] = xor_out[20][11][20] + xor_out[21][11][20] + xor_out[22][11][20] + xor_out[23][11][20] + xor_out[24][11][20];
assign sum_out[5][11][20] = xor_out[25][11][20] + xor_out[26][11][20] + xor_out[27][11][20] + xor_out[28][11][20] + xor_out[29][11][20];
assign sum_out[6][11][20] = xor_out[30][11][20] + xor_out[31][11][20] + xor_out[32][11][20] + xor_out[33][11][20] + xor_out[34][11][20];
assign sum_out[7][11][20] = xor_out[35][11][20] + xor_out[36][11][20] + xor_out[37][11][20] + xor_out[38][11][20] + xor_out[39][11][20];
assign sum_out[8][11][20] = xor_out[40][11][20] + xor_out[41][11][20] + xor_out[42][11][20] + xor_out[43][11][20] + xor_out[44][11][20];
assign sum_out[9][11][20] = xor_out[45][11][20] + xor_out[46][11][20] + xor_out[47][11][20] + xor_out[48][11][20] + xor_out[49][11][20];
assign sum_out[10][11][20] = xor_out[50][11][20] + xor_out[51][11][20] + xor_out[52][11][20] + xor_out[53][11][20] + xor_out[54][11][20];
assign sum_out[11][11][20] = xor_out[55][11][20] + xor_out[56][11][20] + xor_out[57][11][20] + xor_out[58][11][20] + xor_out[59][11][20];
assign sum_out[12][11][20] = xor_out[60][11][20] + xor_out[61][11][20] + xor_out[62][11][20] + xor_out[63][11][20] + xor_out[64][11][20];
assign sum_out[13][11][20] = xor_out[65][11][20] + xor_out[66][11][20] + xor_out[67][11][20] + xor_out[68][11][20] + xor_out[69][11][20];
assign sum_out[14][11][20] = xor_out[70][11][20] + xor_out[71][11][20] + xor_out[72][11][20] + xor_out[73][11][20] + xor_out[74][11][20];
assign sum_out[15][11][20] = xor_out[75][11][20] + xor_out[76][11][20] + xor_out[77][11][20] + xor_out[78][11][20] + xor_out[79][11][20];
assign sum_out[16][11][20] = xor_out[80][11][20] + xor_out[81][11][20] + xor_out[82][11][20] + xor_out[83][11][20] + xor_out[84][11][20];
assign sum_out[17][11][20] = xor_out[85][11][20] + xor_out[86][11][20] + xor_out[87][11][20] + xor_out[88][11][20] + xor_out[89][11][20];
assign sum_out[18][11][20] = xor_out[90][11][20] + xor_out[91][11][20] + xor_out[92][11][20] + xor_out[93][11][20] + xor_out[94][11][20];
assign sum_out[19][11][20] = xor_out[95][11][20] + xor_out[96][11][20] + xor_out[97][11][20] + xor_out[98][11][20] + xor_out[99][11][20];

assign sum_out[0][11][21] = xor_out[0][11][21] + xor_out[1][11][21] + xor_out[2][11][21] + xor_out[3][11][21] + xor_out[4][11][21];
assign sum_out[1][11][21] = xor_out[5][11][21] + xor_out[6][11][21] + xor_out[7][11][21] + xor_out[8][11][21] + xor_out[9][11][21];
assign sum_out[2][11][21] = xor_out[10][11][21] + xor_out[11][11][21] + xor_out[12][11][21] + xor_out[13][11][21] + xor_out[14][11][21];
assign sum_out[3][11][21] = xor_out[15][11][21] + xor_out[16][11][21] + xor_out[17][11][21] + xor_out[18][11][21] + xor_out[19][11][21];
assign sum_out[4][11][21] = xor_out[20][11][21] + xor_out[21][11][21] + xor_out[22][11][21] + xor_out[23][11][21] + xor_out[24][11][21];
assign sum_out[5][11][21] = xor_out[25][11][21] + xor_out[26][11][21] + xor_out[27][11][21] + xor_out[28][11][21] + xor_out[29][11][21];
assign sum_out[6][11][21] = xor_out[30][11][21] + xor_out[31][11][21] + xor_out[32][11][21] + xor_out[33][11][21] + xor_out[34][11][21];
assign sum_out[7][11][21] = xor_out[35][11][21] + xor_out[36][11][21] + xor_out[37][11][21] + xor_out[38][11][21] + xor_out[39][11][21];
assign sum_out[8][11][21] = xor_out[40][11][21] + xor_out[41][11][21] + xor_out[42][11][21] + xor_out[43][11][21] + xor_out[44][11][21];
assign sum_out[9][11][21] = xor_out[45][11][21] + xor_out[46][11][21] + xor_out[47][11][21] + xor_out[48][11][21] + xor_out[49][11][21];
assign sum_out[10][11][21] = xor_out[50][11][21] + xor_out[51][11][21] + xor_out[52][11][21] + xor_out[53][11][21] + xor_out[54][11][21];
assign sum_out[11][11][21] = xor_out[55][11][21] + xor_out[56][11][21] + xor_out[57][11][21] + xor_out[58][11][21] + xor_out[59][11][21];
assign sum_out[12][11][21] = xor_out[60][11][21] + xor_out[61][11][21] + xor_out[62][11][21] + xor_out[63][11][21] + xor_out[64][11][21];
assign sum_out[13][11][21] = xor_out[65][11][21] + xor_out[66][11][21] + xor_out[67][11][21] + xor_out[68][11][21] + xor_out[69][11][21];
assign sum_out[14][11][21] = xor_out[70][11][21] + xor_out[71][11][21] + xor_out[72][11][21] + xor_out[73][11][21] + xor_out[74][11][21];
assign sum_out[15][11][21] = xor_out[75][11][21] + xor_out[76][11][21] + xor_out[77][11][21] + xor_out[78][11][21] + xor_out[79][11][21];
assign sum_out[16][11][21] = xor_out[80][11][21] + xor_out[81][11][21] + xor_out[82][11][21] + xor_out[83][11][21] + xor_out[84][11][21];
assign sum_out[17][11][21] = xor_out[85][11][21] + xor_out[86][11][21] + xor_out[87][11][21] + xor_out[88][11][21] + xor_out[89][11][21];
assign sum_out[18][11][21] = xor_out[90][11][21] + xor_out[91][11][21] + xor_out[92][11][21] + xor_out[93][11][21] + xor_out[94][11][21];
assign sum_out[19][11][21] = xor_out[95][11][21] + xor_out[96][11][21] + xor_out[97][11][21] + xor_out[98][11][21] + xor_out[99][11][21];

assign sum_out[0][11][22] = xor_out[0][11][22] + xor_out[1][11][22] + xor_out[2][11][22] + xor_out[3][11][22] + xor_out[4][11][22];
assign sum_out[1][11][22] = xor_out[5][11][22] + xor_out[6][11][22] + xor_out[7][11][22] + xor_out[8][11][22] + xor_out[9][11][22];
assign sum_out[2][11][22] = xor_out[10][11][22] + xor_out[11][11][22] + xor_out[12][11][22] + xor_out[13][11][22] + xor_out[14][11][22];
assign sum_out[3][11][22] = xor_out[15][11][22] + xor_out[16][11][22] + xor_out[17][11][22] + xor_out[18][11][22] + xor_out[19][11][22];
assign sum_out[4][11][22] = xor_out[20][11][22] + xor_out[21][11][22] + xor_out[22][11][22] + xor_out[23][11][22] + xor_out[24][11][22];
assign sum_out[5][11][22] = xor_out[25][11][22] + xor_out[26][11][22] + xor_out[27][11][22] + xor_out[28][11][22] + xor_out[29][11][22];
assign sum_out[6][11][22] = xor_out[30][11][22] + xor_out[31][11][22] + xor_out[32][11][22] + xor_out[33][11][22] + xor_out[34][11][22];
assign sum_out[7][11][22] = xor_out[35][11][22] + xor_out[36][11][22] + xor_out[37][11][22] + xor_out[38][11][22] + xor_out[39][11][22];
assign sum_out[8][11][22] = xor_out[40][11][22] + xor_out[41][11][22] + xor_out[42][11][22] + xor_out[43][11][22] + xor_out[44][11][22];
assign sum_out[9][11][22] = xor_out[45][11][22] + xor_out[46][11][22] + xor_out[47][11][22] + xor_out[48][11][22] + xor_out[49][11][22];
assign sum_out[10][11][22] = xor_out[50][11][22] + xor_out[51][11][22] + xor_out[52][11][22] + xor_out[53][11][22] + xor_out[54][11][22];
assign sum_out[11][11][22] = xor_out[55][11][22] + xor_out[56][11][22] + xor_out[57][11][22] + xor_out[58][11][22] + xor_out[59][11][22];
assign sum_out[12][11][22] = xor_out[60][11][22] + xor_out[61][11][22] + xor_out[62][11][22] + xor_out[63][11][22] + xor_out[64][11][22];
assign sum_out[13][11][22] = xor_out[65][11][22] + xor_out[66][11][22] + xor_out[67][11][22] + xor_out[68][11][22] + xor_out[69][11][22];
assign sum_out[14][11][22] = xor_out[70][11][22] + xor_out[71][11][22] + xor_out[72][11][22] + xor_out[73][11][22] + xor_out[74][11][22];
assign sum_out[15][11][22] = xor_out[75][11][22] + xor_out[76][11][22] + xor_out[77][11][22] + xor_out[78][11][22] + xor_out[79][11][22];
assign sum_out[16][11][22] = xor_out[80][11][22] + xor_out[81][11][22] + xor_out[82][11][22] + xor_out[83][11][22] + xor_out[84][11][22];
assign sum_out[17][11][22] = xor_out[85][11][22] + xor_out[86][11][22] + xor_out[87][11][22] + xor_out[88][11][22] + xor_out[89][11][22];
assign sum_out[18][11][22] = xor_out[90][11][22] + xor_out[91][11][22] + xor_out[92][11][22] + xor_out[93][11][22] + xor_out[94][11][22];
assign sum_out[19][11][22] = xor_out[95][11][22] + xor_out[96][11][22] + xor_out[97][11][22] + xor_out[98][11][22] + xor_out[99][11][22];

assign sum_out[0][11][23] = xor_out[0][11][23] + xor_out[1][11][23] + xor_out[2][11][23] + xor_out[3][11][23] + xor_out[4][11][23];
assign sum_out[1][11][23] = xor_out[5][11][23] + xor_out[6][11][23] + xor_out[7][11][23] + xor_out[8][11][23] + xor_out[9][11][23];
assign sum_out[2][11][23] = xor_out[10][11][23] + xor_out[11][11][23] + xor_out[12][11][23] + xor_out[13][11][23] + xor_out[14][11][23];
assign sum_out[3][11][23] = xor_out[15][11][23] + xor_out[16][11][23] + xor_out[17][11][23] + xor_out[18][11][23] + xor_out[19][11][23];
assign sum_out[4][11][23] = xor_out[20][11][23] + xor_out[21][11][23] + xor_out[22][11][23] + xor_out[23][11][23] + xor_out[24][11][23];
assign sum_out[5][11][23] = xor_out[25][11][23] + xor_out[26][11][23] + xor_out[27][11][23] + xor_out[28][11][23] + xor_out[29][11][23];
assign sum_out[6][11][23] = xor_out[30][11][23] + xor_out[31][11][23] + xor_out[32][11][23] + xor_out[33][11][23] + xor_out[34][11][23];
assign sum_out[7][11][23] = xor_out[35][11][23] + xor_out[36][11][23] + xor_out[37][11][23] + xor_out[38][11][23] + xor_out[39][11][23];
assign sum_out[8][11][23] = xor_out[40][11][23] + xor_out[41][11][23] + xor_out[42][11][23] + xor_out[43][11][23] + xor_out[44][11][23];
assign sum_out[9][11][23] = xor_out[45][11][23] + xor_out[46][11][23] + xor_out[47][11][23] + xor_out[48][11][23] + xor_out[49][11][23];
assign sum_out[10][11][23] = xor_out[50][11][23] + xor_out[51][11][23] + xor_out[52][11][23] + xor_out[53][11][23] + xor_out[54][11][23];
assign sum_out[11][11][23] = xor_out[55][11][23] + xor_out[56][11][23] + xor_out[57][11][23] + xor_out[58][11][23] + xor_out[59][11][23];
assign sum_out[12][11][23] = xor_out[60][11][23] + xor_out[61][11][23] + xor_out[62][11][23] + xor_out[63][11][23] + xor_out[64][11][23];
assign sum_out[13][11][23] = xor_out[65][11][23] + xor_out[66][11][23] + xor_out[67][11][23] + xor_out[68][11][23] + xor_out[69][11][23];
assign sum_out[14][11][23] = xor_out[70][11][23] + xor_out[71][11][23] + xor_out[72][11][23] + xor_out[73][11][23] + xor_out[74][11][23];
assign sum_out[15][11][23] = xor_out[75][11][23] + xor_out[76][11][23] + xor_out[77][11][23] + xor_out[78][11][23] + xor_out[79][11][23];
assign sum_out[16][11][23] = xor_out[80][11][23] + xor_out[81][11][23] + xor_out[82][11][23] + xor_out[83][11][23] + xor_out[84][11][23];
assign sum_out[17][11][23] = xor_out[85][11][23] + xor_out[86][11][23] + xor_out[87][11][23] + xor_out[88][11][23] + xor_out[89][11][23];
assign sum_out[18][11][23] = xor_out[90][11][23] + xor_out[91][11][23] + xor_out[92][11][23] + xor_out[93][11][23] + xor_out[94][11][23];
assign sum_out[19][11][23] = xor_out[95][11][23] + xor_out[96][11][23] + xor_out[97][11][23] + xor_out[98][11][23] + xor_out[99][11][23];

assign sum_out[0][12][0] = xor_out[0][12][0] + xor_out[1][12][0] + xor_out[2][12][0] + xor_out[3][12][0] + xor_out[4][12][0];
assign sum_out[1][12][0] = xor_out[5][12][0] + xor_out[6][12][0] + xor_out[7][12][0] + xor_out[8][12][0] + xor_out[9][12][0];
assign sum_out[2][12][0] = xor_out[10][12][0] + xor_out[11][12][0] + xor_out[12][12][0] + xor_out[13][12][0] + xor_out[14][12][0];
assign sum_out[3][12][0] = xor_out[15][12][0] + xor_out[16][12][0] + xor_out[17][12][0] + xor_out[18][12][0] + xor_out[19][12][0];
assign sum_out[4][12][0] = xor_out[20][12][0] + xor_out[21][12][0] + xor_out[22][12][0] + xor_out[23][12][0] + xor_out[24][12][0];
assign sum_out[5][12][0] = xor_out[25][12][0] + xor_out[26][12][0] + xor_out[27][12][0] + xor_out[28][12][0] + xor_out[29][12][0];
assign sum_out[6][12][0] = xor_out[30][12][0] + xor_out[31][12][0] + xor_out[32][12][0] + xor_out[33][12][0] + xor_out[34][12][0];
assign sum_out[7][12][0] = xor_out[35][12][0] + xor_out[36][12][0] + xor_out[37][12][0] + xor_out[38][12][0] + xor_out[39][12][0];
assign sum_out[8][12][0] = xor_out[40][12][0] + xor_out[41][12][0] + xor_out[42][12][0] + xor_out[43][12][0] + xor_out[44][12][0];
assign sum_out[9][12][0] = xor_out[45][12][0] + xor_out[46][12][0] + xor_out[47][12][0] + xor_out[48][12][0] + xor_out[49][12][0];
assign sum_out[10][12][0] = xor_out[50][12][0] + xor_out[51][12][0] + xor_out[52][12][0] + xor_out[53][12][0] + xor_out[54][12][0];
assign sum_out[11][12][0] = xor_out[55][12][0] + xor_out[56][12][0] + xor_out[57][12][0] + xor_out[58][12][0] + xor_out[59][12][0];
assign sum_out[12][12][0] = xor_out[60][12][0] + xor_out[61][12][0] + xor_out[62][12][0] + xor_out[63][12][0] + xor_out[64][12][0];
assign sum_out[13][12][0] = xor_out[65][12][0] + xor_out[66][12][0] + xor_out[67][12][0] + xor_out[68][12][0] + xor_out[69][12][0];
assign sum_out[14][12][0] = xor_out[70][12][0] + xor_out[71][12][0] + xor_out[72][12][0] + xor_out[73][12][0] + xor_out[74][12][0];
assign sum_out[15][12][0] = xor_out[75][12][0] + xor_out[76][12][0] + xor_out[77][12][0] + xor_out[78][12][0] + xor_out[79][12][0];
assign sum_out[16][12][0] = xor_out[80][12][0] + xor_out[81][12][0] + xor_out[82][12][0] + xor_out[83][12][0] + xor_out[84][12][0];
assign sum_out[17][12][0] = xor_out[85][12][0] + xor_out[86][12][0] + xor_out[87][12][0] + xor_out[88][12][0] + xor_out[89][12][0];
assign sum_out[18][12][0] = xor_out[90][12][0] + xor_out[91][12][0] + xor_out[92][12][0] + xor_out[93][12][0] + xor_out[94][12][0];
assign sum_out[19][12][0] = xor_out[95][12][0] + xor_out[96][12][0] + xor_out[97][12][0] + xor_out[98][12][0] + xor_out[99][12][0];

assign sum_out[0][12][1] = xor_out[0][12][1] + xor_out[1][12][1] + xor_out[2][12][1] + xor_out[3][12][1] + xor_out[4][12][1];
assign sum_out[1][12][1] = xor_out[5][12][1] + xor_out[6][12][1] + xor_out[7][12][1] + xor_out[8][12][1] + xor_out[9][12][1];
assign sum_out[2][12][1] = xor_out[10][12][1] + xor_out[11][12][1] + xor_out[12][12][1] + xor_out[13][12][1] + xor_out[14][12][1];
assign sum_out[3][12][1] = xor_out[15][12][1] + xor_out[16][12][1] + xor_out[17][12][1] + xor_out[18][12][1] + xor_out[19][12][1];
assign sum_out[4][12][1] = xor_out[20][12][1] + xor_out[21][12][1] + xor_out[22][12][1] + xor_out[23][12][1] + xor_out[24][12][1];
assign sum_out[5][12][1] = xor_out[25][12][1] + xor_out[26][12][1] + xor_out[27][12][1] + xor_out[28][12][1] + xor_out[29][12][1];
assign sum_out[6][12][1] = xor_out[30][12][1] + xor_out[31][12][1] + xor_out[32][12][1] + xor_out[33][12][1] + xor_out[34][12][1];
assign sum_out[7][12][1] = xor_out[35][12][1] + xor_out[36][12][1] + xor_out[37][12][1] + xor_out[38][12][1] + xor_out[39][12][1];
assign sum_out[8][12][1] = xor_out[40][12][1] + xor_out[41][12][1] + xor_out[42][12][1] + xor_out[43][12][1] + xor_out[44][12][1];
assign sum_out[9][12][1] = xor_out[45][12][1] + xor_out[46][12][1] + xor_out[47][12][1] + xor_out[48][12][1] + xor_out[49][12][1];
assign sum_out[10][12][1] = xor_out[50][12][1] + xor_out[51][12][1] + xor_out[52][12][1] + xor_out[53][12][1] + xor_out[54][12][1];
assign sum_out[11][12][1] = xor_out[55][12][1] + xor_out[56][12][1] + xor_out[57][12][1] + xor_out[58][12][1] + xor_out[59][12][1];
assign sum_out[12][12][1] = xor_out[60][12][1] + xor_out[61][12][1] + xor_out[62][12][1] + xor_out[63][12][1] + xor_out[64][12][1];
assign sum_out[13][12][1] = xor_out[65][12][1] + xor_out[66][12][1] + xor_out[67][12][1] + xor_out[68][12][1] + xor_out[69][12][1];
assign sum_out[14][12][1] = xor_out[70][12][1] + xor_out[71][12][1] + xor_out[72][12][1] + xor_out[73][12][1] + xor_out[74][12][1];
assign sum_out[15][12][1] = xor_out[75][12][1] + xor_out[76][12][1] + xor_out[77][12][1] + xor_out[78][12][1] + xor_out[79][12][1];
assign sum_out[16][12][1] = xor_out[80][12][1] + xor_out[81][12][1] + xor_out[82][12][1] + xor_out[83][12][1] + xor_out[84][12][1];
assign sum_out[17][12][1] = xor_out[85][12][1] + xor_out[86][12][1] + xor_out[87][12][1] + xor_out[88][12][1] + xor_out[89][12][1];
assign sum_out[18][12][1] = xor_out[90][12][1] + xor_out[91][12][1] + xor_out[92][12][1] + xor_out[93][12][1] + xor_out[94][12][1];
assign sum_out[19][12][1] = xor_out[95][12][1] + xor_out[96][12][1] + xor_out[97][12][1] + xor_out[98][12][1] + xor_out[99][12][1];

assign sum_out[0][12][2] = xor_out[0][12][2] + xor_out[1][12][2] + xor_out[2][12][2] + xor_out[3][12][2] + xor_out[4][12][2];
assign sum_out[1][12][2] = xor_out[5][12][2] + xor_out[6][12][2] + xor_out[7][12][2] + xor_out[8][12][2] + xor_out[9][12][2];
assign sum_out[2][12][2] = xor_out[10][12][2] + xor_out[11][12][2] + xor_out[12][12][2] + xor_out[13][12][2] + xor_out[14][12][2];
assign sum_out[3][12][2] = xor_out[15][12][2] + xor_out[16][12][2] + xor_out[17][12][2] + xor_out[18][12][2] + xor_out[19][12][2];
assign sum_out[4][12][2] = xor_out[20][12][2] + xor_out[21][12][2] + xor_out[22][12][2] + xor_out[23][12][2] + xor_out[24][12][2];
assign sum_out[5][12][2] = xor_out[25][12][2] + xor_out[26][12][2] + xor_out[27][12][2] + xor_out[28][12][2] + xor_out[29][12][2];
assign sum_out[6][12][2] = xor_out[30][12][2] + xor_out[31][12][2] + xor_out[32][12][2] + xor_out[33][12][2] + xor_out[34][12][2];
assign sum_out[7][12][2] = xor_out[35][12][2] + xor_out[36][12][2] + xor_out[37][12][2] + xor_out[38][12][2] + xor_out[39][12][2];
assign sum_out[8][12][2] = xor_out[40][12][2] + xor_out[41][12][2] + xor_out[42][12][2] + xor_out[43][12][2] + xor_out[44][12][2];
assign sum_out[9][12][2] = xor_out[45][12][2] + xor_out[46][12][2] + xor_out[47][12][2] + xor_out[48][12][2] + xor_out[49][12][2];
assign sum_out[10][12][2] = xor_out[50][12][2] + xor_out[51][12][2] + xor_out[52][12][2] + xor_out[53][12][2] + xor_out[54][12][2];
assign sum_out[11][12][2] = xor_out[55][12][2] + xor_out[56][12][2] + xor_out[57][12][2] + xor_out[58][12][2] + xor_out[59][12][2];
assign sum_out[12][12][2] = xor_out[60][12][2] + xor_out[61][12][2] + xor_out[62][12][2] + xor_out[63][12][2] + xor_out[64][12][2];
assign sum_out[13][12][2] = xor_out[65][12][2] + xor_out[66][12][2] + xor_out[67][12][2] + xor_out[68][12][2] + xor_out[69][12][2];
assign sum_out[14][12][2] = xor_out[70][12][2] + xor_out[71][12][2] + xor_out[72][12][2] + xor_out[73][12][2] + xor_out[74][12][2];
assign sum_out[15][12][2] = xor_out[75][12][2] + xor_out[76][12][2] + xor_out[77][12][2] + xor_out[78][12][2] + xor_out[79][12][2];
assign sum_out[16][12][2] = xor_out[80][12][2] + xor_out[81][12][2] + xor_out[82][12][2] + xor_out[83][12][2] + xor_out[84][12][2];
assign sum_out[17][12][2] = xor_out[85][12][2] + xor_out[86][12][2] + xor_out[87][12][2] + xor_out[88][12][2] + xor_out[89][12][2];
assign sum_out[18][12][2] = xor_out[90][12][2] + xor_out[91][12][2] + xor_out[92][12][2] + xor_out[93][12][2] + xor_out[94][12][2];
assign sum_out[19][12][2] = xor_out[95][12][2] + xor_out[96][12][2] + xor_out[97][12][2] + xor_out[98][12][2] + xor_out[99][12][2];

assign sum_out[0][12][3] = xor_out[0][12][3] + xor_out[1][12][3] + xor_out[2][12][3] + xor_out[3][12][3] + xor_out[4][12][3];
assign sum_out[1][12][3] = xor_out[5][12][3] + xor_out[6][12][3] + xor_out[7][12][3] + xor_out[8][12][3] + xor_out[9][12][3];
assign sum_out[2][12][3] = xor_out[10][12][3] + xor_out[11][12][3] + xor_out[12][12][3] + xor_out[13][12][3] + xor_out[14][12][3];
assign sum_out[3][12][3] = xor_out[15][12][3] + xor_out[16][12][3] + xor_out[17][12][3] + xor_out[18][12][3] + xor_out[19][12][3];
assign sum_out[4][12][3] = xor_out[20][12][3] + xor_out[21][12][3] + xor_out[22][12][3] + xor_out[23][12][3] + xor_out[24][12][3];
assign sum_out[5][12][3] = xor_out[25][12][3] + xor_out[26][12][3] + xor_out[27][12][3] + xor_out[28][12][3] + xor_out[29][12][3];
assign sum_out[6][12][3] = xor_out[30][12][3] + xor_out[31][12][3] + xor_out[32][12][3] + xor_out[33][12][3] + xor_out[34][12][3];
assign sum_out[7][12][3] = xor_out[35][12][3] + xor_out[36][12][3] + xor_out[37][12][3] + xor_out[38][12][3] + xor_out[39][12][3];
assign sum_out[8][12][3] = xor_out[40][12][3] + xor_out[41][12][3] + xor_out[42][12][3] + xor_out[43][12][3] + xor_out[44][12][3];
assign sum_out[9][12][3] = xor_out[45][12][3] + xor_out[46][12][3] + xor_out[47][12][3] + xor_out[48][12][3] + xor_out[49][12][3];
assign sum_out[10][12][3] = xor_out[50][12][3] + xor_out[51][12][3] + xor_out[52][12][3] + xor_out[53][12][3] + xor_out[54][12][3];
assign sum_out[11][12][3] = xor_out[55][12][3] + xor_out[56][12][3] + xor_out[57][12][3] + xor_out[58][12][3] + xor_out[59][12][3];
assign sum_out[12][12][3] = xor_out[60][12][3] + xor_out[61][12][3] + xor_out[62][12][3] + xor_out[63][12][3] + xor_out[64][12][3];
assign sum_out[13][12][3] = xor_out[65][12][3] + xor_out[66][12][3] + xor_out[67][12][3] + xor_out[68][12][3] + xor_out[69][12][3];
assign sum_out[14][12][3] = xor_out[70][12][3] + xor_out[71][12][3] + xor_out[72][12][3] + xor_out[73][12][3] + xor_out[74][12][3];
assign sum_out[15][12][3] = xor_out[75][12][3] + xor_out[76][12][3] + xor_out[77][12][3] + xor_out[78][12][3] + xor_out[79][12][3];
assign sum_out[16][12][3] = xor_out[80][12][3] + xor_out[81][12][3] + xor_out[82][12][3] + xor_out[83][12][3] + xor_out[84][12][3];
assign sum_out[17][12][3] = xor_out[85][12][3] + xor_out[86][12][3] + xor_out[87][12][3] + xor_out[88][12][3] + xor_out[89][12][3];
assign sum_out[18][12][3] = xor_out[90][12][3] + xor_out[91][12][3] + xor_out[92][12][3] + xor_out[93][12][3] + xor_out[94][12][3];
assign sum_out[19][12][3] = xor_out[95][12][3] + xor_out[96][12][3] + xor_out[97][12][3] + xor_out[98][12][3] + xor_out[99][12][3];

assign sum_out[0][12][4] = xor_out[0][12][4] + xor_out[1][12][4] + xor_out[2][12][4] + xor_out[3][12][4] + xor_out[4][12][4];
assign sum_out[1][12][4] = xor_out[5][12][4] + xor_out[6][12][4] + xor_out[7][12][4] + xor_out[8][12][4] + xor_out[9][12][4];
assign sum_out[2][12][4] = xor_out[10][12][4] + xor_out[11][12][4] + xor_out[12][12][4] + xor_out[13][12][4] + xor_out[14][12][4];
assign sum_out[3][12][4] = xor_out[15][12][4] + xor_out[16][12][4] + xor_out[17][12][4] + xor_out[18][12][4] + xor_out[19][12][4];
assign sum_out[4][12][4] = xor_out[20][12][4] + xor_out[21][12][4] + xor_out[22][12][4] + xor_out[23][12][4] + xor_out[24][12][4];
assign sum_out[5][12][4] = xor_out[25][12][4] + xor_out[26][12][4] + xor_out[27][12][4] + xor_out[28][12][4] + xor_out[29][12][4];
assign sum_out[6][12][4] = xor_out[30][12][4] + xor_out[31][12][4] + xor_out[32][12][4] + xor_out[33][12][4] + xor_out[34][12][4];
assign sum_out[7][12][4] = xor_out[35][12][4] + xor_out[36][12][4] + xor_out[37][12][4] + xor_out[38][12][4] + xor_out[39][12][4];
assign sum_out[8][12][4] = xor_out[40][12][4] + xor_out[41][12][4] + xor_out[42][12][4] + xor_out[43][12][4] + xor_out[44][12][4];
assign sum_out[9][12][4] = xor_out[45][12][4] + xor_out[46][12][4] + xor_out[47][12][4] + xor_out[48][12][4] + xor_out[49][12][4];
assign sum_out[10][12][4] = xor_out[50][12][4] + xor_out[51][12][4] + xor_out[52][12][4] + xor_out[53][12][4] + xor_out[54][12][4];
assign sum_out[11][12][4] = xor_out[55][12][4] + xor_out[56][12][4] + xor_out[57][12][4] + xor_out[58][12][4] + xor_out[59][12][4];
assign sum_out[12][12][4] = xor_out[60][12][4] + xor_out[61][12][4] + xor_out[62][12][4] + xor_out[63][12][4] + xor_out[64][12][4];
assign sum_out[13][12][4] = xor_out[65][12][4] + xor_out[66][12][4] + xor_out[67][12][4] + xor_out[68][12][4] + xor_out[69][12][4];
assign sum_out[14][12][4] = xor_out[70][12][4] + xor_out[71][12][4] + xor_out[72][12][4] + xor_out[73][12][4] + xor_out[74][12][4];
assign sum_out[15][12][4] = xor_out[75][12][4] + xor_out[76][12][4] + xor_out[77][12][4] + xor_out[78][12][4] + xor_out[79][12][4];
assign sum_out[16][12][4] = xor_out[80][12][4] + xor_out[81][12][4] + xor_out[82][12][4] + xor_out[83][12][4] + xor_out[84][12][4];
assign sum_out[17][12][4] = xor_out[85][12][4] + xor_out[86][12][4] + xor_out[87][12][4] + xor_out[88][12][4] + xor_out[89][12][4];
assign sum_out[18][12][4] = xor_out[90][12][4] + xor_out[91][12][4] + xor_out[92][12][4] + xor_out[93][12][4] + xor_out[94][12][4];
assign sum_out[19][12][4] = xor_out[95][12][4] + xor_out[96][12][4] + xor_out[97][12][4] + xor_out[98][12][4] + xor_out[99][12][4];

assign sum_out[0][12][5] = xor_out[0][12][5] + xor_out[1][12][5] + xor_out[2][12][5] + xor_out[3][12][5] + xor_out[4][12][5];
assign sum_out[1][12][5] = xor_out[5][12][5] + xor_out[6][12][5] + xor_out[7][12][5] + xor_out[8][12][5] + xor_out[9][12][5];
assign sum_out[2][12][5] = xor_out[10][12][5] + xor_out[11][12][5] + xor_out[12][12][5] + xor_out[13][12][5] + xor_out[14][12][5];
assign sum_out[3][12][5] = xor_out[15][12][5] + xor_out[16][12][5] + xor_out[17][12][5] + xor_out[18][12][5] + xor_out[19][12][5];
assign sum_out[4][12][5] = xor_out[20][12][5] + xor_out[21][12][5] + xor_out[22][12][5] + xor_out[23][12][5] + xor_out[24][12][5];
assign sum_out[5][12][5] = xor_out[25][12][5] + xor_out[26][12][5] + xor_out[27][12][5] + xor_out[28][12][5] + xor_out[29][12][5];
assign sum_out[6][12][5] = xor_out[30][12][5] + xor_out[31][12][5] + xor_out[32][12][5] + xor_out[33][12][5] + xor_out[34][12][5];
assign sum_out[7][12][5] = xor_out[35][12][5] + xor_out[36][12][5] + xor_out[37][12][5] + xor_out[38][12][5] + xor_out[39][12][5];
assign sum_out[8][12][5] = xor_out[40][12][5] + xor_out[41][12][5] + xor_out[42][12][5] + xor_out[43][12][5] + xor_out[44][12][5];
assign sum_out[9][12][5] = xor_out[45][12][5] + xor_out[46][12][5] + xor_out[47][12][5] + xor_out[48][12][5] + xor_out[49][12][5];
assign sum_out[10][12][5] = xor_out[50][12][5] + xor_out[51][12][5] + xor_out[52][12][5] + xor_out[53][12][5] + xor_out[54][12][5];
assign sum_out[11][12][5] = xor_out[55][12][5] + xor_out[56][12][5] + xor_out[57][12][5] + xor_out[58][12][5] + xor_out[59][12][5];
assign sum_out[12][12][5] = xor_out[60][12][5] + xor_out[61][12][5] + xor_out[62][12][5] + xor_out[63][12][5] + xor_out[64][12][5];
assign sum_out[13][12][5] = xor_out[65][12][5] + xor_out[66][12][5] + xor_out[67][12][5] + xor_out[68][12][5] + xor_out[69][12][5];
assign sum_out[14][12][5] = xor_out[70][12][5] + xor_out[71][12][5] + xor_out[72][12][5] + xor_out[73][12][5] + xor_out[74][12][5];
assign sum_out[15][12][5] = xor_out[75][12][5] + xor_out[76][12][5] + xor_out[77][12][5] + xor_out[78][12][5] + xor_out[79][12][5];
assign sum_out[16][12][5] = xor_out[80][12][5] + xor_out[81][12][5] + xor_out[82][12][5] + xor_out[83][12][5] + xor_out[84][12][5];
assign sum_out[17][12][5] = xor_out[85][12][5] + xor_out[86][12][5] + xor_out[87][12][5] + xor_out[88][12][5] + xor_out[89][12][5];
assign sum_out[18][12][5] = xor_out[90][12][5] + xor_out[91][12][5] + xor_out[92][12][5] + xor_out[93][12][5] + xor_out[94][12][5];
assign sum_out[19][12][5] = xor_out[95][12][5] + xor_out[96][12][5] + xor_out[97][12][5] + xor_out[98][12][5] + xor_out[99][12][5];

assign sum_out[0][12][6] = xor_out[0][12][6] + xor_out[1][12][6] + xor_out[2][12][6] + xor_out[3][12][6] + xor_out[4][12][6];
assign sum_out[1][12][6] = xor_out[5][12][6] + xor_out[6][12][6] + xor_out[7][12][6] + xor_out[8][12][6] + xor_out[9][12][6];
assign sum_out[2][12][6] = xor_out[10][12][6] + xor_out[11][12][6] + xor_out[12][12][6] + xor_out[13][12][6] + xor_out[14][12][6];
assign sum_out[3][12][6] = xor_out[15][12][6] + xor_out[16][12][6] + xor_out[17][12][6] + xor_out[18][12][6] + xor_out[19][12][6];
assign sum_out[4][12][6] = xor_out[20][12][6] + xor_out[21][12][6] + xor_out[22][12][6] + xor_out[23][12][6] + xor_out[24][12][6];
assign sum_out[5][12][6] = xor_out[25][12][6] + xor_out[26][12][6] + xor_out[27][12][6] + xor_out[28][12][6] + xor_out[29][12][6];
assign sum_out[6][12][6] = xor_out[30][12][6] + xor_out[31][12][6] + xor_out[32][12][6] + xor_out[33][12][6] + xor_out[34][12][6];
assign sum_out[7][12][6] = xor_out[35][12][6] + xor_out[36][12][6] + xor_out[37][12][6] + xor_out[38][12][6] + xor_out[39][12][6];
assign sum_out[8][12][6] = xor_out[40][12][6] + xor_out[41][12][6] + xor_out[42][12][6] + xor_out[43][12][6] + xor_out[44][12][6];
assign sum_out[9][12][6] = xor_out[45][12][6] + xor_out[46][12][6] + xor_out[47][12][6] + xor_out[48][12][6] + xor_out[49][12][6];
assign sum_out[10][12][6] = xor_out[50][12][6] + xor_out[51][12][6] + xor_out[52][12][6] + xor_out[53][12][6] + xor_out[54][12][6];
assign sum_out[11][12][6] = xor_out[55][12][6] + xor_out[56][12][6] + xor_out[57][12][6] + xor_out[58][12][6] + xor_out[59][12][6];
assign sum_out[12][12][6] = xor_out[60][12][6] + xor_out[61][12][6] + xor_out[62][12][6] + xor_out[63][12][6] + xor_out[64][12][6];
assign sum_out[13][12][6] = xor_out[65][12][6] + xor_out[66][12][6] + xor_out[67][12][6] + xor_out[68][12][6] + xor_out[69][12][6];
assign sum_out[14][12][6] = xor_out[70][12][6] + xor_out[71][12][6] + xor_out[72][12][6] + xor_out[73][12][6] + xor_out[74][12][6];
assign sum_out[15][12][6] = xor_out[75][12][6] + xor_out[76][12][6] + xor_out[77][12][6] + xor_out[78][12][6] + xor_out[79][12][6];
assign sum_out[16][12][6] = xor_out[80][12][6] + xor_out[81][12][6] + xor_out[82][12][6] + xor_out[83][12][6] + xor_out[84][12][6];
assign sum_out[17][12][6] = xor_out[85][12][6] + xor_out[86][12][6] + xor_out[87][12][6] + xor_out[88][12][6] + xor_out[89][12][6];
assign sum_out[18][12][6] = xor_out[90][12][6] + xor_out[91][12][6] + xor_out[92][12][6] + xor_out[93][12][6] + xor_out[94][12][6];
assign sum_out[19][12][6] = xor_out[95][12][6] + xor_out[96][12][6] + xor_out[97][12][6] + xor_out[98][12][6] + xor_out[99][12][6];

assign sum_out[0][12][7] = xor_out[0][12][7] + xor_out[1][12][7] + xor_out[2][12][7] + xor_out[3][12][7] + xor_out[4][12][7];
assign sum_out[1][12][7] = xor_out[5][12][7] + xor_out[6][12][7] + xor_out[7][12][7] + xor_out[8][12][7] + xor_out[9][12][7];
assign sum_out[2][12][7] = xor_out[10][12][7] + xor_out[11][12][7] + xor_out[12][12][7] + xor_out[13][12][7] + xor_out[14][12][7];
assign sum_out[3][12][7] = xor_out[15][12][7] + xor_out[16][12][7] + xor_out[17][12][7] + xor_out[18][12][7] + xor_out[19][12][7];
assign sum_out[4][12][7] = xor_out[20][12][7] + xor_out[21][12][7] + xor_out[22][12][7] + xor_out[23][12][7] + xor_out[24][12][7];
assign sum_out[5][12][7] = xor_out[25][12][7] + xor_out[26][12][7] + xor_out[27][12][7] + xor_out[28][12][7] + xor_out[29][12][7];
assign sum_out[6][12][7] = xor_out[30][12][7] + xor_out[31][12][7] + xor_out[32][12][7] + xor_out[33][12][7] + xor_out[34][12][7];
assign sum_out[7][12][7] = xor_out[35][12][7] + xor_out[36][12][7] + xor_out[37][12][7] + xor_out[38][12][7] + xor_out[39][12][7];
assign sum_out[8][12][7] = xor_out[40][12][7] + xor_out[41][12][7] + xor_out[42][12][7] + xor_out[43][12][7] + xor_out[44][12][7];
assign sum_out[9][12][7] = xor_out[45][12][7] + xor_out[46][12][7] + xor_out[47][12][7] + xor_out[48][12][7] + xor_out[49][12][7];
assign sum_out[10][12][7] = xor_out[50][12][7] + xor_out[51][12][7] + xor_out[52][12][7] + xor_out[53][12][7] + xor_out[54][12][7];
assign sum_out[11][12][7] = xor_out[55][12][7] + xor_out[56][12][7] + xor_out[57][12][7] + xor_out[58][12][7] + xor_out[59][12][7];
assign sum_out[12][12][7] = xor_out[60][12][7] + xor_out[61][12][7] + xor_out[62][12][7] + xor_out[63][12][7] + xor_out[64][12][7];
assign sum_out[13][12][7] = xor_out[65][12][7] + xor_out[66][12][7] + xor_out[67][12][7] + xor_out[68][12][7] + xor_out[69][12][7];
assign sum_out[14][12][7] = xor_out[70][12][7] + xor_out[71][12][7] + xor_out[72][12][7] + xor_out[73][12][7] + xor_out[74][12][7];
assign sum_out[15][12][7] = xor_out[75][12][7] + xor_out[76][12][7] + xor_out[77][12][7] + xor_out[78][12][7] + xor_out[79][12][7];
assign sum_out[16][12][7] = xor_out[80][12][7] + xor_out[81][12][7] + xor_out[82][12][7] + xor_out[83][12][7] + xor_out[84][12][7];
assign sum_out[17][12][7] = xor_out[85][12][7] + xor_out[86][12][7] + xor_out[87][12][7] + xor_out[88][12][7] + xor_out[89][12][7];
assign sum_out[18][12][7] = xor_out[90][12][7] + xor_out[91][12][7] + xor_out[92][12][7] + xor_out[93][12][7] + xor_out[94][12][7];
assign sum_out[19][12][7] = xor_out[95][12][7] + xor_out[96][12][7] + xor_out[97][12][7] + xor_out[98][12][7] + xor_out[99][12][7];

assign sum_out[0][12][8] = xor_out[0][12][8] + xor_out[1][12][8] + xor_out[2][12][8] + xor_out[3][12][8] + xor_out[4][12][8];
assign sum_out[1][12][8] = xor_out[5][12][8] + xor_out[6][12][8] + xor_out[7][12][8] + xor_out[8][12][8] + xor_out[9][12][8];
assign sum_out[2][12][8] = xor_out[10][12][8] + xor_out[11][12][8] + xor_out[12][12][8] + xor_out[13][12][8] + xor_out[14][12][8];
assign sum_out[3][12][8] = xor_out[15][12][8] + xor_out[16][12][8] + xor_out[17][12][8] + xor_out[18][12][8] + xor_out[19][12][8];
assign sum_out[4][12][8] = xor_out[20][12][8] + xor_out[21][12][8] + xor_out[22][12][8] + xor_out[23][12][8] + xor_out[24][12][8];
assign sum_out[5][12][8] = xor_out[25][12][8] + xor_out[26][12][8] + xor_out[27][12][8] + xor_out[28][12][8] + xor_out[29][12][8];
assign sum_out[6][12][8] = xor_out[30][12][8] + xor_out[31][12][8] + xor_out[32][12][8] + xor_out[33][12][8] + xor_out[34][12][8];
assign sum_out[7][12][8] = xor_out[35][12][8] + xor_out[36][12][8] + xor_out[37][12][8] + xor_out[38][12][8] + xor_out[39][12][8];
assign sum_out[8][12][8] = xor_out[40][12][8] + xor_out[41][12][8] + xor_out[42][12][8] + xor_out[43][12][8] + xor_out[44][12][8];
assign sum_out[9][12][8] = xor_out[45][12][8] + xor_out[46][12][8] + xor_out[47][12][8] + xor_out[48][12][8] + xor_out[49][12][8];
assign sum_out[10][12][8] = xor_out[50][12][8] + xor_out[51][12][8] + xor_out[52][12][8] + xor_out[53][12][8] + xor_out[54][12][8];
assign sum_out[11][12][8] = xor_out[55][12][8] + xor_out[56][12][8] + xor_out[57][12][8] + xor_out[58][12][8] + xor_out[59][12][8];
assign sum_out[12][12][8] = xor_out[60][12][8] + xor_out[61][12][8] + xor_out[62][12][8] + xor_out[63][12][8] + xor_out[64][12][8];
assign sum_out[13][12][8] = xor_out[65][12][8] + xor_out[66][12][8] + xor_out[67][12][8] + xor_out[68][12][8] + xor_out[69][12][8];
assign sum_out[14][12][8] = xor_out[70][12][8] + xor_out[71][12][8] + xor_out[72][12][8] + xor_out[73][12][8] + xor_out[74][12][8];
assign sum_out[15][12][8] = xor_out[75][12][8] + xor_out[76][12][8] + xor_out[77][12][8] + xor_out[78][12][8] + xor_out[79][12][8];
assign sum_out[16][12][8] = xor_out[80][12][8] + xor_out[81][12][8] + xor_out[82][12][8] + xor_out[83][12][8] + xor_out[84][12][8];
assign sum_out[17][12][8] = xor_out[85][12][8] + xor_out[86][12][8] + xor_out[87][12][8] + xor_out[88][12][8] + xor_out[89][12][8];
assign sum_out[18][12][8] = xor_out[90][12][8] + xor_out[91][12][8] + xor_out[92][12][8] + xor_out[93][12][8] + xor_out[94][12][8];
assign sum_out[19][12][8] = xor_out[95][12][8] + xor_out[96][12][8] + xor_out[97][12][8] + xor_out[98][12][8] + xor_out[99][12][8];

assign sum_out[0][12][9] = xor_out[0][12][9] + xor_out[1][12][9] + xor_out[2][12][9] + xor_out[3][12][9] + xor_out[4][12][9];
assign sum_out[1][12][9] = xor_out[5][12][9] + xor_out[6][12][9] + xor_out[7][12][9] + xor_out[8][12][9] + xor_out[9][12][9];
assign sum_out[2][12][9] = xor_out[10][12][9] + xor_out[11][12][9] + xor_out[12][12][9] + xor_out[13][12][9] + xor_out[14][12][9];
assign sum_out[3][12][9] = xor_out[15][12][9] + xor_out[16][12][9] + xor_out[17][12][9] + xor_out[18][12][9] + xor_out[19][12][9];
assign sum_out[4][12][9] = xor_out[20][12][9] + xor_out[21][12][9] + xor_out[22][12][9] + xor_out[23][12][9] + xor_out[24][12][9];
assign sum_out[5][12][9] = xor_out[25][12][9] + xor_out[26][12][9] + xor_out[27][12][9] + xor_out[28][12][9] + xor_out[29][12][9];
assign sum_out[6][12][9] = xor_out[30][12][9] + xor_out[31][12][9] + xor_out[32][12][9] + xor_out[33][12][9] + xor_out[34][12][9];
assign sum_out[7][12][9] = xor_out[35][12][9] + xor_out[36][12][9] + xor_out[37][12][9] + xor_out[38][12][9] + xor_out[39][12][9];
assign sum_out[8][12][9] = xor_out[40][12][9] + xor_out[41][12][9] + xor_out[42][12][9] + xor_out[43][12][9] + xor_out[44][12][9];
assign sum_out[9][12][9] = xor_out[45][12][9] + xor_out[46][12][9] + xor_out[47][12][9] + xor_out[48][12][9] + xor_out[49][12][9];
assign sum_out[10][12][9] = xor_out[50][12][9] + xor_out[51][12][9] + xor_out[52][12][9] + xor_out[53][12][9] + xor_out[54][12][9];
assign sum_out[11][12][9] = xor_out[55][12][9] + xor_out[56][12][9] + xor_out[57][12][9] + xor_out[58][12][9] + xor_out[59][12][9];
assign sum_out[12][12][9] = xor_out[60][12][9] + xor_out[61][12][9] + xor_out[62][12][9] + xor_out[63][12][9] + xor_out[64][12][9];
assign sum_out[13][12][9] = xor_out[65][12][9] + xor_out[66][12][9] + xor_out[67][12][9] + xor_out[68][12][9] + xor_out[69][12][9];
assign sum_out[14][12][9] = xor_out[70][12][9] + xor_out[71][12][9] + xor_out[72][12][9] + xor_out[73][12][9] + xor_out[74][12][9];
assign sum_out[15][12][9] = xor_out[75][12][9] + xor_out[76][12][9] + xor_out[77][12][9] + xor_out[78][12][9] + xor_out[79][12][9];
assign sum_out[16][12][9] = xor_out[80][12][9] + xor_out[81][12][9] + xor_out[82][12][9] + xor_out[83][12][9] + xor_out[84][12][9];
assign sum_out[17][12][9] = xor_out[85][12][9] + xor_out[86][12][9] + xor_out[87][12][9] + xor_out[88][12][9] + xor_out[89][12][9];
assign sum_out[18][12][9] = xor_out[90][12][9] + xor_out[91][12][9] + xor_out[92][12][9] + xor_out[93][12][9] + xor_out[94][12][9];
assign sum_out[19][12][9] = xor_out[95][12][9] + xor_out[96][12][9] + xor_out[97][12][9] + xor_out[98][12][9] + xor_out[99][12][9];

assign sum_out[0][12][10] = xor_out[0][12][10] + xor_out[1][12][10] + xor_out[2][12][10] + xor_out[3][12][10] + xor_out[4][12][10];
assign sum_out[1][12][10] = xor_out[5][12][10] + xor_out[6][12][10] + xor_out[7][12][10] + xor_out[8][12][10] + xor_out[9][12][10];
assign sum_out[2][12][10] = xor_out[10][12][10] + xor_out[11][12][10] + xor_out[12][12][10] + xor_out[13][12][10] + xor_out[14][12][10];
assign sum_out[3][12][10] = xor_out[15][12][10] + xor_out[16][12][10] + xor_out[17][12][10] + xor_out[18][12][10] + xor_out[19][12][10];
assign sum_out[4][12][10] = xor_out[20][12][10] + xor_out[21][12][10] + xor_out[22][12][10] + xor_out[23][12][10] + xor_out[24][12][10];
assign sum_out[5][12][10] = xor_out[25][12][10] + xor_out[26][12][10] + xor_out[27][12][10] + xor_out[28][12][10] + xor_out[29][12][10];
assign sum_out[6][12][10] = xor_out[30][12][10] + xor_out[31][12][10] + xor_out[32][12][10] + xor_out[33][12][10] + xor_out[34][12][10];
assign sum_out[7][12][10] = xor_out[35][12][10] + xor_out[36][12][10] + xor_out[37][12][10] + xor_out[38][12][10] + xor_out[39][12][10];
assign sum_out[8][12][10] = xor_out[40][12][10] + xor_out[41][12][10] + xor_out[42][12][10] + xor_out[43][12][10] + xor_out[44][12][10];
assign sum_out[9][12][10] = xor_out[45][12][10] + xor_out[46][12][10] + xor_out[47][12][10] + xor_out[48][12][10] + xor_out[49][12][10];
assign sum_out[10][12][10] = xor_out[50][12][10] + xor_out[51][12][10] + xor_out[52][12][10] + xor_out[53][12][10] + xor_out[54][12][10];
assign sum_out[11][12][10] = xor_out[55][12][10] + xor_out[56][12][10] + xor_out[57][12][10] + xor_out[58][12][10] + xor_out[59][12][10];
assign sum_out[12][12][10] = xor_out[60][12][10] + xor_out[61][12][10] + xor_out[62][12][10] + xor_out[63][12][10] + xor_out[64][12][10];
assign sum_out[13][12][10] = xor_out[65][12][10] + xor_out[66][12][10] + xor_out[67][12][10] + xor_out[68][12][10] + xor_out[69][12][10];
assign sum_out[14][12][10] = xor_out[70][12][10] + xor_out[71][12][10] + xor_out[72][12][10] + xor_out[73][12][10] + xor_out[74][12][10];
assign sum_out[15][12][10] = xor_out[75][12][10] + xor_out[76][12][10] + xor_out[77][12][10] + xor_out[78][12][10] + xor_out[79][12][10];
assign sum_out[16][12][10] = xor_out[80][12][10] + xor_out[81][12][10] + xor_out[82][12][10] + xor_out[83][12][10] + xor_out[84][12][10];
assign sum_out[17][12][10] = xor_out[85][12][10] + xor_out[86][12][10] + xor_out[87][12][10] + xor_out[88][12][10] + xor_out[89][12][10];
assign sum_out[18][12][10] = xor_out[90][12][10] + xor_out[91][12][10] + xor_out[92][12][10] + xor_out[93][12][10] + xor_out[94][12][10];
assign sum_out[19][12][10] = xor_out[95][12][10] + xor_out[96][12][10] + xor_out[97][12][10] + xor_out[98][12][10] + xor_out[99][12][10];

assign sum_out[0][12][11] = xor_out[0][12][11] + xor_out[1][12][11] + xor_out[2][12][11] + xor_out[3][12][11] + xor_out[4][12][11];
assign sum_out[1][12][11] = xor_out[5][12][11] + xor_out[6][12][11] + xor_out[7][12][11] + xor_out[8][12][11] + xor_out[9][12][11];
assign sum_out[2][12][11] = xor_out[10][12][11] + xor_out[11][12][11] + xor_out[12][12][11] + xor_out[13][12][11] + xor_out[14][12][11];
assign sum_out[3][12][11] = xor_out[15][12][11] + xor_out[16][12][11] + xor_out[17][12][11] + xor_out[18][12][11] + xor_out[19][12][11];
assign sum_out[4][12][11] = xor_out[20][12][11] + xor_out[21][12][11] + xor_out[22][12][11] + xor_out[23][12][11] + xor_out[24][12][11];
assign sum_out[5][12][11] = xor_out[25][12][11] + xor_out[26][12][11] + xor_out[27][12][11] + xor_out[28][12][11] + xor_out[29][12][11];
assign sum_out[6][12][11] = xor_out[30][12][11] + xor_out[31][12][11] + xor_out[32][12][11] + xor_out[33][12][11] + xor_out[34][12][11];
assign sum_out[7][12][11] = xor_out[35][12][11] + xor_out[36][12][11] + xor_out[37][12][11] + xor_out[38][12][11] + xor_out[39][12][11];
assign sum_out[8][12][11] = xor_out[40][12][11] + xor_out[41][12][11] + xor_out[42][12][11] + xor_out[43][12][11] + xor_out[44][12][11];
assign sum_out[9][12][11] = xor_out[45][12][11] + xor_out[46][12][11] + xor_out[47][12][11] + xor_out[48][12][11] + xor_out[49][12][11];
assign sum_out[10][12][11] = xor_out[50][12][11] + xor_out[51][12][11] + xor_out[52][12][11] + xor_out[53][12][11] + xor_out[54][12][11];
assign sum_out[11][12][11] = xor_out[55][12][11] + xor_out[56][12][11] + xor_out[57][12][11] + xor_out[58][12][11] + xor_out[59][12][11];
assign sum_out[12][12][11] = xor_out[60][12][11] + xor_out[61][12][11] + xor_out[62][12][11] + xor_out[63][12][11] + xor_out[64][12][11];
assign sum_out[13][12][11] = xor_out[65][12][11] + xor_out[66][12][11] + xor_out[67][12][11] + xor_out[68][12][11] + xor_out[69][12][11];
assign sum_out[14][12][11] = xor_out[70][12][11] + xor_out[71][12][11] + xor_out[72][12][11] + xor_out[73][12][11] + xor_out[74][12][11];
assign sum_out[15][12][11] = xor_out[75][12][11] + xor_out[76][12][11] + xor_out[77][12][11] + xor_out[78][12][11] + xor_out[79][12][11];
assign sum_out[16][12][11] = xor_out[80][12][11] + xor_out[81][12][11] + xor_out[82][12][11] + xor_out[83][12][11] + xor_out[84][12][11];
assign sum_out[17][12][11] = xor_out[85][12][11] + xor_out[86][12][11] + xor_out[87][12][11] + xor_out[88][12][11] + xor_out[89][12][11];
assign sum_out[18][12][11] = xor_out[90][12][11] + xor_out[91][12][11] + xor_out[92][12][11] + xor_out[93][12][11] + xor_out[94][12][11];
assign sum_out[19][12][11] = xor_out[95][12][11] + xor_out[96][12][11] + xor_out[97][12][11] + xor_out[98][12][11] + xor_out[99][12][11];

assign sum_out[0][12][12] = xor_out[0][12][12] + xor_out[1][12][12] + xor_out[2][12][12] + xor_out[3][12][12] + xor_out[4][12][12];
assign sum_out[1][12][12] = xor_out[5][12][12] + xor_out[6][12][12] + xor_out[7][12][12] + xor_out[8][12][12] + xor_out[9][12][12];
assign sum_out[2][12][12] = xor_out[10][12][12] + xor_out[11][12][12] + xor_out[12][12][12] + xor_out[13][12][12] + xor_out[14][12][12];
assign sum_out[3][12][12] = xor_out[15][12][12] + xor_out[16][12][12] + xor_out[17][12][12] + xor_out[18][12][12] + xor_out[19][12][12];
assign sum_out[4][12][12] = xor_out[20][12][12] + xor_out[21][12][12] + xor_out[22][12][12] + xor_out[23][12][12] + xor_out[24][12][12];
assign sum_out[5][12][12] = xor_out[25][12][12] + xor_out[26][12][12] + xor_out[27][12][12] + xor_out[28][12][12] + xor_out[29][12][12];
assign sum_out[6][12][12] = xor_out[30][12][12] + xor_out[31][12][12] + xor_out[32][12][12] + xor_out[33][12][12] + xor_out[34][12][12];
assign sum_out[7][12][12] = xor_out[35][12][12] + xor_out[36][12][12] + xor_out[37][12][12] + xor_out[38][12][12] + xor_out[39][12][12];
assign sum_out[8][12][12] = xor_out[40][12][12] + xor_out[41][12][12] + xor_out[42][12][12] + xor_out[43][12][12] + xor_out[44][12][12];
assign sum_out[9][12][12] = xor_out[45][12][12] + xor_out[46][12][12] + xor_out[47][12][12] + xor_out[48][12][12] + xor_out[49][12][12];
assign sum_out[10][12][12] = xor_out[50][12][12] + xor_out[51][12][12] + xor_out[52][12][12] + xor_out[53][12][12] + xor_out[54][12][12];
assign sum_out[11][12][12] = xor_out[55][12][12] + xor_out[56][12][12] + xor_out[57][12][12] + xor_out[58][12][12] + xor_out[59][12][12];
assign sum_out[12][12][12] = xor_out[60][12][12] + xor_out[61][12][12] + xor_out[62][12][12] + xor_out[63][12][12] + xor_out[64][12][12];
assign sum_out[13][12][12] = xor_out[65][12][12] + xor_out[66][12][12] + xor_out[67][12][12] + xor_out[68][12][12] + xor_out[69][12][12];
assign sum_out[14][12][12] = xor_out[70][12][12] + xor_out[71][12][12] + xor_out[72][12][12] + xor_out[73][12][12] + xor_out[74][12][12];
assign sum_out[15][12][12] = xor_out[75][12][12] + xor_out[76][12][12] + xor_out[77][12][12] + xor_out[78][12][12] + xor_out[79][12][12];
assign sum_out[16][12][12] = xor_out[80][12][12] + xor_out[81][12][12] + xor_out[82][12][12] + xor_out[83][12][12] + xor_out[84][12][12];
assign sum_out[17][12][12] = xor_out[85][12][12] + xor_out[86][12][12] + xor_out[87][12][12] + xor_out[88][12][12] + xor_out[89][12][12];
assign sum_out[18][12][12] = xor_out[90][12][12] + xor_out[91][12][12] + xor_out[92][12][12] + xor_out[93][12][12] + xor_out[94][12][12];
assign sum_out[19][12][12] = xor_out[95][12][12] + xor_out[96][12][12] + xor_out[97][12][12] + xor_out[98][12][12] + xor_out[99][12][12];

assign sum_out[0][12][13] = xor_out[0][12][13] + xor_out[1][12][13] + xor_out[2][12][13] + xor_out[3][12][13] + xor_out[4][12][13];
assign sum_out[1][12][13] = xor_out[5][12][13] + xor_out[6][12][13] + xor_out[7][12][13] + xor_out[8][12][13] + xor_out[9][12][13];
assign sum_out[2][12][13] = xor_out[10][12][13] + xor_out[11][12][13] + xor_out[12][12][13] + xor_out[13][12][13] + xor_out[14][12][13];
assign sum_out[3][12][13] = xor_out[15][12][13] + xor_out[16][12][13] + xor_out[17][12][13] + xor_out[18][12][13] + xor_out[19][12][13];
assign sum_out[4][12][13] = xor_out[20][12][13] + xor_out[21][12][13] + xor_out[22][12][13] + xor_out[23][12][13] + xor_out[24][12][13];
assign sum_out[5][12][13] = xor_out[25][12][13] + xor_out[26][12][13] + xor_out[27][12][13] + xor_out[28][12][13] + xor_out[29][12][13];
assign sum_out[6][12][13] = xor_out[30][12][13] + xor_out[31][12][13] + xor_out[32][12][13] + xor_out[33][12][13] + xor_out[34][12][13];
assign sum_out[7][12][13] = xor_out[35][12][13] + xor_out[36][12][13] + xor_out[37][12][13] + xor_out[38][12][13] + xor_out[39][12][13];
assign sum_out[8][12][13] = xor_out[40][12][13] + xor_out[41][12][13] + xor_out[42][12][13] + xor_out[43][12][13] + xor_out[44][12][13];
assign sum_out[9][12][13] = xor_out[45][12][13] + xor_out[46][12][13] + xor_out[47][12][13] + xor_out[48][12][13] + xor_out[49][12][13];
assign sum_out[10][12][13] = xor_out[50][12][13] + xor_out[51][12][13] + xor_out[52][12][13] + xor_out[53][12][13] + xor_out[54][12][13];
assign sum_out[11][12][13] = xor_out[55][12][13] + xor_out[56][12][13] + xor_out[57][12][13] + xor_out[58][12][13] + xor_out[59][12][13];
assign sum_out[12][12][13] = xor_out[60][12][13] + xor_out[61][12][13] + xor_out[62][12][13] + xor_out[63][12][13] + xor_out[64][12][13];
assign sum_out[13][12][13] = xor_out[65][12][13] + xor_out[66][12][13] + xor_out[67][12][13] + xor_out[68][12][13] + xor_out[69][12][13];
assign sum_out[14][12][13] = xor_out[70][12][13] + xor_out[71][12][13] + xor_out[72][12][13] + xor_out[73][12][13] + xor_out[74][12][13];
assign sum_out[15][12][13] = xor_out[75][12][13] + xor_out[76][12][13] + xor_out[77][12][13] + xor_out[78][12][13] + xor_out[79][12][13];
assign sum_out[16][12][13] = xor_out[80][12][13] + xor_out[81][12][13] + xor_out[82][12][13] + xor_out[83][12][13] + xor_out[84][12][13];
assign sum_out[17][12][13] = xor_out[85][12][13] + xor_out[86][12][13] + xor_out[87][12][13] + xor_out[88][12][13] + xor_out[89][12][13];
assign sum_out[18][12][13] = xor_out[90][12][13] + xor_out[91][12][13] + xor_out[92][12][13] + xor_out[93][12][13] + xor_out[94][12][13];
assign sum_out[19][12][13] = xor_out[95][12][13] + xor_out[96][12][13] + xor_out[97][12][13] + xor_out[98][12][13] + xor_out[99][12][13];

assign sum_out[0][12][14] = xor_out[0][12][14] + xor_out[1][12][14] + xor_out[2][12][14] + xor_out[3][12][14] + xor_out[4][12][14];
assign sum_out[1][12][14] = xor_out[5][12][14] + xor_out[6][12][14] + xor_out[7][12][14] + xor_out[8][12][14] + xor_out[9][12][14];
assign sum_out[2][12][14] = xor_out[10][12][14] + xor_out[11][12][14] + xor_out[12][12][14] + xor_out[13][12][14] + xor_out[14][12][14];
assign sum_out[3][12][14] = xor_out[15][12][14] + xor_out[16][12][14] + xor_out[17][12][14] + xor_out[18][12][14] + xor_out[19][12][14];
assign sum_out[4][12][14] = xor_out[20][12][14] + xor_out[21][12][14] + xor_out[22][12][14] + xor_out[23][12][14] + xor_out[24][12][14];
assign sum_out[5][12][14] = xor_out[25][12][14] + xor_out[26][12][14] + xor_out[27][12][14] + xor_out[28][12][14] + xor_out[29][12][14];
assign sum_out[6][12][14] = xor_out[30][12][14] + xor_out[31][12][14] + xor_out[32][12][14] + xor_out[33][12][14] + xor_out[34][12][14];
assign sum_out[7][12][14] = xor_out[35][12][14] + xor_out[36][12][14] + xor_out[37][12][14] + xor_out[38][12][14] + xor_out[39][12][14];
assign sum_out[8][12][14] = xor_out[40][12][14] + xor_out[41][12][14] + xor_out[42][12][14] + xor_out[43][12][14] + xor_out[44][12][14];
assign sum_out[9][12][14] = xor_out[45][12][14] + xor_out[46][12][14] + xor_out[47][12][14] + xor_out[48][12][14] + xor_out[49][12][14];
assign sum_out[10][12][14] = xor_out[50][12][14] + xor_out[51][12][14] + xor_out[52][12][14] + xor_out[53][12][14] + xor_out[54][12][14];
assign sum_out[11][12][14] = xor_out[55][12][14] + xor_out[56][12][14] + xor_out[57][12][14] + xor_out[58][12][14] + xor_out[59][12][14];
assign sum_out[12][12][14] = xor_out[60][12][14] + xor_out[61][12][14] + xor_out[62][12][14] + xor_out[63][12][14] + xor_out[64][12][14];
assign sum_out[13][12][14] = xor_out[65][12][14] + xor_out[66][12][14] + xor_out[67][12][14] + xor_out[68][12][14] + xor_out[69][12][14];
assign sum_out[14][12][14] = xor_out[70][12][14] + xor_out[71][12][14] + xor_out[72][12][14] + xor_out[73][12][14] + xor_out[74][12][14];
assign sum_out[15][12][14] = xor_out[75][12][14] + xor_out[76][12][14] + xor_out[77][12][14] + xor_out[78][12][14] + xor_out[79][12][14];
assign sum_out[16][12][14] = xor_out[80][12][14] + xor_out[81][12][14] + xor_out[82][12][14] + xor_out[83][12][14] + xor_out[84][12][14];
assign sum_out[17][12][14] = xor_out[85][12][14] + xor_out[86][12][14] + xor_out[87][12][14] + xor_out[88][12][14] + xor_out[89][12][14];
assign sum_out[18][12][14] = xor_out[90][12][14] + xor_out[91][12][14] + xor_out[92][12][14] + xor_out[93][12][14] + xor_out[94][12][14];
assign sum_out[19][12][14] = xor_out[95][12][14] + xor_out[96][12][14] + xor_out[97][12][14] + xor_out[98][12][14] + xor_out[99][12][14];

assign sum_out[0][12][15] = xor_out[0][12][15] + xor_out[1][12][15] + xor_out[2][12][15] + xor_out[3][12][15] + xor_out[4][12][15];
assign sum_out[1][12][15] = xor_out[5][12][15] + xor_out[6][12][15] + xor_out[7][12][15] + xor_out[8][12][15] + xor_out[9][12][15];
assign sum_out[2][12][15] = xor_out[10][12][15] + xor_out[11][12][15] + xor_out[12][12][15] + xor_out[13][12][15] + xor_out[14][12][15];
assign sum_out[3][12][15] = xor_out[15][12][15] + xor_out[16][12][15] + xor_out[17][12][15] + xor_out[18][12][15] + xor_out[19][12][15];
assign sum_out[4][12][15] = xor_out[20][12][15] + xor_out[21][12][15] + xor_out[22][12][15] + xor_out[23][12][15] + xor_out[24][12][15];
assign sum_out[5][12][15] = xor_out[25][12][15] + xor_out[26][12][15] + xor_out[27][12][15] + xor_out[28][12][15] + xor_out[29][12][15];
assign sum_out[6][12][15] = xor_out[30][12][15] + xor_out[31][12][15] + xor_out[32][12][15] + xor_out[33][12][15] + xor_out[34][12][15];
assign sum_out[7][12][15] = xor_out[35][12][15] + xor_out[36][12][15] + xor_out[37][12][15] + xor_out[38][12][15] + xor_out[39][12][15];
assign sum_out[8][12][15] = xor_out[40][12][15] + xor_out[41][12][15] + xor_out[42][12][15] + xor_out[43][12][15] + xor_out[44][12][15];
assign sum_out[9][12][15] = xor_out[45][12][15] + xor_out[46][12][15] + xor_out[47][12][15] + xor_out[48][12][15] + xor_out[49][12][15];
assign sum_out[10][12][15] = xor_out[50][12][15] + xor_out[51][12][15] + xor_out[52][12][15] + xor_out[53][12][15] + xor_out[54][12][15];
assign sum_out[11][12][15] = xor_out[55][12][15] + xor_out[56][12][15] + xor_out[57][12][15] + xor_out[58][12][15] + xor_out[59][12][15];
assign sum_out[12][12][15] = xor_out[60][12][15] + xor_out[61][12][15] + xor_out[62][12][15] + xor_out[63][12][15] + xor_out[64][12][15];
assign sum_out[13][12][15] = xor_out[65][12][15] + xor_out[66][12][15] + xor_out[67][12][15] + xor_out[68][12][15] + xor_out[69][12][15];
assign sum_out[14][12][15] = xor_out[70][12][15] + xor_out[71][12][15] + xor_out[72][12][15] + xor_out[73][12][15] + xor_out[74][12][15];
assign sum_out[15][12][15] = xor_out[75][12][15] + xor_out[76][12][15] + xor_out[77][12][15] + xor_out[78][12][15] + xor_out[79][12][15];
assign sum_out[16][12][15] = xor_out[80][12][15] + xor_out[81][12][15] + xor_out[82][12][15] + xor_out[83][12][15] + xor_out[84][12][15];
assign sum_out[17][12][15] = xor_out[85][12][15] + xor_out[86][12][15] + xor_out[87][12][15] + xor_out[88][12][15] + xor_out[89][12][15];
assign sum_out[18][12][15] = xor_out[90][12][15] + xor_out[91][12][15] + xor_out[92][12][15] + xor_out[93][12][15] + xor_out[94][12][15];
assign sum_out[19][12][15] = xor_out[95][12][15] + xor_out[96][12][15] + xor_out[97][12][15] + xor_out[98][12][15] + xor_out[99][12][15];

assign sum_out[0][12][16] = xor_out[0][12][16] + xor_out[1][12][16] + xor_out[2][12][16] + xor_out[3][12][16] + xor_out[4][12][16];
assign sum_out[1][12][16] = xor_out[5][12][16] + xor_out[6][12][16] + xor_out[7][12][16] + xor_out[8][12][16] + xor_out[9][12][16];
assign sum_out[2][12][16] = xor_out[10][12][16] + xor_out[11][12][16] + xor_out[12][12][16] + xor_out[13][12][16] + xor_out[14][12][16];
assign sum_out[3][12][16] = xor_out[15][12][16] + xor_out[16][12][16] + xor_out[17][12][16] + xor_out[18][12][16] + xor_out[19][12][16];
assign sum_out[4][12][16] = xor_out[20][12][16] + xor_out[21][12][16] + xor_out[22][12][16] + xor_out[23][12][16] + xor_out[24][12][16];
assign sum_out[5][12][16] = xor_out[25][12][16] + xor_out[26][12][16] + xor_out[27][12][16] + xor_out[28][12][16] + xor_out[29][12][16];
assign sum_out[6][12][16] = xor_out[30][12][16] + xor_out[31][12][16] + xor_out[32][12][16] + xor_out[33][12][16] + xor_out[34][12][16];
assign sum_out[7][12][16] = xor_out[35][12][16] + xor_out[36][12][16] + xor_out[37][12][16] + xor_out[38][12][16] + xor_out[39][12][16];
assign sum_out[8][12][16] = xor_out[40][12][16] + xor_out[41][12][16] + xor_out[42][12][16] + xor_out[43][12][16] + xor_out[44][12][16];
assign sum_out[9][12][16] = xor_out[45][12][16] + xor_out[46][12][16] + xor_out[47][12][16] + xor_out[48][12][16] + xor_out[49][12][16];
assign sum_out[10][12][16] = xor_out[50][12][16] + xor_out[51][12][16] + xor_out[52][12][16] + xor_out[53][12][16] + xor_out[54][12][16];
assign sum_out[11][12][16] = xor_out[55][12][16] + xor_out[56][12][16] + xor_out[57][12][16] + xor_out[58][12][16] + xor_out[59][12][16];
assign sum_out[12][12][16] = xor_out[60][12][16] + xor_out[61][12][16] + xor_out[62][12][16] + xor_out[63][12][16] + xor_out[64][12][16];
assign sum_out[13][12][16] = xor_out[65][12][16] + xor_out[66][12][16] + xor_out[67][12][16] + xor_out[68][12][16] + xor_out[69][12][16];
assign sum_out[14][12][16] = xor_out[70][12][16] + xor_out[71][12][16] + xor_out[72][12][16] + xor_out[73][12][16] + xor_out[74][12][16];
assign sum_out[15][12][16] = xor_out[75][12][16] + xor_out[76][12][16] + xor_out[77][12][16] + xor_out[78][12][16] + xor_out[79][12][16];
assign sum_out[16][12][16] = xor_out[80][12][16] + xor_out[81][12][16] + xor_out[82][12][16] + xor_out[83][12][16] + xor_out[84][12][16];
assign sum_out[17][12][16] = xor_out[85][12][16] + xor_out[86][12][16] + xor_out[87][12][16] + xor_out[88][12][16] + xor_out[89][12][16];
assign sum_out[18][12][16] = xor_out[90][12][16] + xor_out[91][12][16] + xor_out[92][12][16] + xor_out[93][12][16] + xor_out[94][12][16];
assign sum_out[19][12][16] = xor_out[95][12][16] + xor_out[96][12][16] + xor_out[97][12][16] + xor_out[98][12][16] + xor_out[99][12][16];

assign sum_out[0][12][17] = xor_out[0][12][17] + xor_out[1][12][17] + xor_out[2][12][17] + xor_out[3][12][17] + xor_out[4][12][17];
assign sum_out[1][12][17] = xor_out[5][12][17] + xor_out[6][12][17] + xor_out[7][12][17] + xor_out[8][12][17] + xor_out[9][12][17];
assign sum_out[2][12][17] = xor_out[10][12][17] + xor_out[11][12][17] + xor_out[12][12][17] + xor_out[13][12][17] + xor_out[14][12][17];
assign sum_out[3][12][17] = xor_out[15][12][17] + xor_out[16][12][17] + xor_out[17][12][17] + xor_out[18][12][17] + xor_out[19][12][17];
assign sum_out[4][12][17] = xor_out[20][12][17] + xor_out[21][12][17] + xor_out[22][12][17] + xor_out[23][12][17] + xor_out[24][12][17];
assign sum_out[5][12][17] = xor_out[25][12][17] + xor_out[26][12][17] + xor_out[27][12][17] + xor_out[28][12][17] + xor_out[29][12][17];
assign sum_out[6][12][17] = xor_out[30][12][17] + xor_out[31][12][17] + xor_out[32][12][17] + xor_out[33][12][17] + xor_out[34][12][17];
assign sum_out[7][12][17] = xor_out[35][12][17] + xor_out[36][12][17] + xor_out[37][12][17] + xor_out[38][12][17] + xor_out[39][12][17];
assign sum_out[8][12][17] = xor_out[40][12][17] + xor_out[41][12][17] + xor_out[42][12][17] + xor_out[43][12][17] + xor_out[44][12][17];
assign sum_out[9][12][17] = xor_out[45][12][17] + xor_out[46][12][17] + xor_out[47][12][17] + xor_out[48][12][17] + xor_out[49][12][17];
assign sum_out[10][12][17] = xor_out[50][12][17] + xor_out[51][12][17] + xor_out[52][12][17] + xor_out[53][12][17] + xor_out[54][12][17];
assign sum_out[11][12][17] = xor_out[55][12][17] + xor_out[56][12][17] + xor_out[57][12][17] + xor_out[58][12][17] + xor_out[59][12][17];
assign sum_out[12][12][17] = xor_out[60][12][17] + xor_out[61][12][17] + xor_out[62][12][17] + xor_out[63][12][17] + xor_out[64][12][17];
assign sum_out[13][12][17] = xor_out[65][12][17] + xor_out[66][12][17] + xor_out[67][12][17] + xor_out[68][12][17] + xor_out[69][12][17];
assign sum_out[14][12][17] = xor_out[70][12][17] + xor_out[71][12][17] + xor_out[72][12][17] + xor_out[73][12][17] + xor_out[74][12][17];
assign sum_out[15][12][17] = xor_out[75][12][17] + xor_out[76][12][17] + xor_out[77][12][17] + xor_out[78][12][17] + xor_out[79][12][17];
assign sum_out[16][12][17] = xor_out[80][12][17] + xor_out[81][12][17] + xor_out[82][12][17] + xor_out[83][12][17] + xor_out[84][12][17];
assign sum_out[17][12][17] = xor_out[85][12][17] + xor_out[86][12][17] + xor_out[87][12][17] + xor_out[88][12][17] + xor_out[89][12][17];
assign sum_out[18][12][17] = xor_out[90][12][17] + xor_out[91][12][17] + xor_out[92][12][17] + xor_out[93][12][17] + xor_out[94][12][17];
assign sum_out[19][12][17] = xor_out[95][12][17] + xor_out[96][12][17] + xor_out[97][12][17] + xor_out[98][12][17] + xor_out[99][12][17];

assign sum_out[0][12][18] = xor_out[0][12][18] + xor_out[1][12][18] + xor_out[2][12][18] + xor_out[3][12][18] + xor_out[4][12][18];
assign sum_out[1][12][18] = xor_out[5][12][18] + xor_out[6][12][18] + xor_out[7][12][18] + xor_out[8][12][18] + xor_out[9][12][18];
assign sum_out[2][12][18] = xor_out[10][12][18] + xor_out[11][12][18] + xor_out[12][12][18] + xor_out[13][12][18] + xor_out[14][12][18];
assign sum_out[3][12][18] = xor_out[15][12][18] + xor_out[16][12][18] + xor_out[17][12][18] + xor_out[18][12][18] + xor_out[19][12][18];
assign sum_out[4][12][18] = xor_out[20][12][18] + xor_out[21][12][18] + xor_out[22][12][18] + xor_out[23][12][18] + xor_out[24][12][18];
assign sum_out[5][12][18] = xor_out[25][12][18] + xor_out[26][12][18] + xor_out[27][12][18] + xor_out[28][12][18] + xor_out[29][12][18];
assign sum_out[6][12][18] = xor_out[30][12][18] + xor_out[31][12][18] + xor_out[32][12][18] + xor_out[33][12][18] + xor_out[34][12][18];
assign sum_out[7][12][18] = xor_out[35][12][18] + xor_out[36][12][18] + xor_out[37][12][18] + xor_out[38][12][18] + xor_out[39][12][18];
assign sum_out[8][12][18] = xor_out[40][12][18] + xor_out[41][12][18] + xor_out[42][12][18] + xor_out[43][12][18] + xor_out[44][12][18];
assign sum_out[9][12][18] = xor_out[45][12][18] + xor_out[46][12][18] + xor_out[47][12][18] + xor_out[48][12][18] + xor_out[49][12][18];
assign sum_out[10][12][18] = xor_out[50][12][18] + xor_out[51][12][18] + xor_out[52][12][18] + xor_out[53][12][18] + xor_out[54][12][18];
assign sum_out[11][12][18] = xor_out[55][12][18] + xor_out[56][12][18] + xor_out[57][12][18] + xor_out[58][12][18] + xor_out[59][12][18];
assign sum_out[12][12][18] = xor_out[60][12][18] + xor_out[61][12][18] + xor_out[62][12][18] + xor_out[63][12][18] + xor_out[64][12][18];
assign sum_out[13][12][18] = xor_out[65][12][18] + xor_out[66][12][18] + xor_out[67][12][18] + xor_out[68][12][18] + xor_out[69][12][18];
assign sum_out[14][12][18] = xor_out[70][12][18] + xor_out[71][12][18] + xor_out[72][12][18] + xor_out[73][12][18] + xor_out[74][12][18];
assign sum_out[15][12][18] = xor_out[75][12][18] + xor_out[76][12][18] + xor_out[77][12][18] + xor_out[78][12][18] + xor_out[79][12][18];
assign sum_out[16][12][18] = xor_out[80][12][18] + xor_out[81][12][18] + xor_out[82][12][18] + xor_out[83][12][18] + xor_out[84][12][18];
assign sum_out[17][12][18] = xor_out[85][12][18] + xor_out[86][12][18] + xor_out[87][12][18] + xor_out[88][12][18] + xor_out[89][12][18];
assign sum_out[18][12][18] = xor_out[90][12][18] + xor_out[91][12][18] + xor_out[92][12][18] + xor_out[93][12][18] + xor_out[94][12][18];
assign sum_out[19][12][18] = xor_out[95][12][18] + xor_out[96][12][18] + xor_out[97][12][18] + xor_out[98][12][18] + xor_out[99][12][18];

assign sum_out[0][12][19] = xor_out[0][12][19] + xor_out[1][12][19] + xor_out[2][12][19] + xor_out[3][12][19] + xor_out[4][12][19];
assign sum_out[1][12][19] = xor_out[5][12][19] + xor_out[6][12][19] + xor_out[7][12][19] + xor_out[8][12][19] + xor_out[9][12][19];
assign sum_out[2][12][19] = xor_out[10][12][19] + xor_out[11][12][19] + xor_out[12][12][19] + xor_out[13][12][19] + xor_out[14][12][19];
assign sum_out[3][12][19] = xor_out[15][12][19] + xor_out[16][12][19] + xor_out[17][12][19] + xor_out[18][12][19] + xor_out[19][12][19];
assign sum_out[4][12][19] = xor_out[20][12][19] + xor_out[21][12][19] + xor_out[22][12][19] + xor_out[23][12][19] + xor_out[24][12][19];
assign sum_out[5][12][19] = xor_out[25][12][19] + xor_out[26][12][19] + xor_out[27][12][19] + xor_out[28][12][19] + xor_out[29][12][19];
assign sum_out[6][12][19] = xor_out[30][12][19] + xor_out[31][12][19] + xor_out[32][12][19] + xor_out[33][12][19] + xor_out[34][12][19];
assign sum_out[7][12][19] = xor_out[35][12][19] + xor_out[36][12][19] + xor_out[37][12][19] + xor_out[38][12][19] + xor_out[39][12][19];
assign sum_out[8][12][19] = xor_out[40][12][19] + xor_out[41][12][19] + xor_out[42][12][19] + xor_out[43][12][19] + xor_out[44][12][19];
assign sum_out[9][12][19] = xor_out[45][12][19] + xor_out[46][12][19] + xor_out[47][12][19] + xor_out[48][12][19] + xor_out[49][12][19];
assign sum_out[10][12][19] = xor_out[50][12][19] + xor_out[51][12][19] + xor_out[52][12][19] + xor_out[53][12][19] + xor_out[54][12][19];
assign sum_out[11][12][19] = xor_out[55][12][19] + xor_out[56][12][19] + xor_out[57][12][19] + xor_out[58][12][19] + xor_out[59][12][19];
assign sum_out[12][12][19] = xor_out[60][12][19] + xor_out[61][12][19] + xor_out[62][12][19] + xor_out[63][12][19] + xor_out[64][12][19];
assign sum_out[13][12][19] = xor_out[65][12][19] + xor_out[66][12][19] + xor_out[67][12][19] + xor_out[68][12][19] + xor_out[69][12][19];
assign sum_out[14][12][19] = xor_out[70][12][19] + xor_out[71][12][19] + xor_out[72][12][19] + xor_out[73][12][19] + xor_out[74][12][19];
assign sum_out[15][12][19] = xor_out[75][12][19] + xor_out[76][12][19] + xor_out[77][12][19] + xor_out[78][12][19] + xor_out[79][12][19];
assign sum_out[16][12][19] = xor_out[80][12][19] + xor_out[81][12][19] + xor_out[82][12][19] + xor_out[83][12][19] + xor_out[84][12][19];
assign sum_out[17][12][19] = xor_out[85][12][19] + xor_out[86][12][19] + xor_out[87][12][19] + xor_out[88][12][19] + xor_out[89][12][19];
assign sum_out[18][12][19] = xor_out[90][12][19] + xor_out[91][12][19] + xor_out[92][12][19] + xor_out[93][12][19] + xor_out[94][12][19];
assign sum_out[19][12][19] = xor_out[95][12][19] + xor_out[96][12][19] + xor_out[97][12][19] + xor_out[98][12][19] + xor_out[99][12][19];

assign sum_out[0][12][20] = xor_out[0][12][20] + xor_out[1][12][20] + xor_out[2][12][20] + xor_out[3][12][20] + xor_out[4][12][20];
assign sum_out[1][12][20] = xor_out[5][12][20] + xor_out[6][12][20] + xor_out[7][12][20] + xor_out[8][12][20] + xor_out[9][12][20];
assign sum_out[2][12][20] = xor_out[10][12][20] + xor_out[11][12][20] + xor_out[12][12][20] + xor_out[13][12][20] + xor_out[14][12][20];
assign sum_out[3][12][20] = xor_out[15][12][20] + xor_out[16][12][20] + xor_out[17][12][20] + xor_out[18][12][20] + xor_out[19][12][20];
assign sum_out[4][12][20] = xor_out[20][12][20] + xor_out[21][12][20] + xor_out[22][12][20] + xor_out[23][12][20] + xor_out[24][12][20];
assign sum_out[5][12][20] = xor_out[25][12][20] + xor_out[26][12][20] + xor_out[27][12][20] + xor_out[28][12][20] + xor_out[29][12][20];
assign sum_out[6][12][20] = xor_out[30][12][20] + xor_out[31][12][20] + xor_out[32][12][20] + xor_out[33][12][20] + xor_out[34][12][20];
assign sum_out[7][12][20] = xor_out[35][12][20] + xor_out[36][12][20] + xor_out[37][12][20] + xor_out[38][12][20] + xor_out[39][12][20];
assign sum_out[8][12][20] = xor_out[40][12][20] + xor_out[41][12][20] + xor_out[42][12][20] + xor_out[43][12][20] + xor_out[44][12][20];
assign sum_out[9][12][20] = xor_out[45][12][20] + xor_out[46][12][20] + xor_out[47][12][20] + xor_out[48][12][20] + xor_out[49][12][20];
assign sum_out[10][12][20] = xor_out[50][12][20] + xor_out[51][12][20] + xor_out[52][12][20] + xor_out[53][12][20] + xor_out[54][12][20];
assign sum_out[11][12][20] = xor_out[55][12][20] + xor_out[56][12][20] + xor_out[57][12][20] + xor_out[58][12][20] + xor_out[59][12][20];
assign sum_out[12][12][20] = xor_out[60][12][20] + xor_out[61][12][20] + xor_out[62][12][20] + xor_out[63][12][20] + xor_out[64][12][20];
assign sum_out[13][12][20] = xor_out[65][12][20] + xor_out[66][12][20] + xor_out[67][12][20] + xor_out[68][12][20] + xor_out[69][12][20];
assign sum_out[14][12][20] = xor_out[70][12][20] + xor_out[71][12][20] + xor_out[72][12][20] + xor_out[73][12][20] + xor_out[74][12][20];
assign sum_out[15][12][20] = xor_out[75][12][20] + xor_out[76][12][20] + xor_out[77][12][20] + xor_out[78][12][20] + xor_out[79][12][20];
assign sum_out[16][12][20] = xor_out[80][12][20] + xor_out[81][12][20] + xor_out[82][12][20] + xor_out[83][12][20] + xor_out[84][12][20];
assign sum_out[17][12][20] = xor_out[85][12][20] + xor_out[86][12][20] + xor_out[87][12][20] + xor_out[88][12][20] + xor_out[89][12][20];
assign sum_out[18][12][20] = xor_out[90][12][20] + xor_out[91][12][20] + xor_out[92][12][20] + xor_out[93][12][20] + xor_out[94][12][20];
assign sum_out[19][12][20] = xor_out[95][12][20] + xor_out[96][12][20] + xor_out[97][12][20] + xor_out[98][12][20] + xor_out[99][12][20];

assign sum_out[0][12][21] = xor_out[0][12][21] + xor_out[1][12][21] + xor_out[2][12][21] + xor_out[3][12][21] + xor_out[4][12][21];
assign sum_out[1][12][21] = xor_out[5][12][21] + xor_out[6][12][21] + xor_out[7][12][21] + xor_out[8][12][21] + xor_out[9][12][21];
assign sum_out[2][12][21] = xor_out[10][12][21] + xor_out[11][12][21] + xor_out[12][12][21] + xor_out[13][12][21] + xor_out[14][12][21];
assign sum_out[3][12][21] = xor_out[15][12][21] + xor_out[16][12][21] + xor_out[17][12][21] + xor_out[18][12][21] + xor_out[19][12][21];
assign sum_out[4][12][21] = xor_out[20][12][21] + xor_out[21][12][21] + xor_out[22][12][21] + xor_out[23][12][21] + xor_out[24][12][21];
assign sum_out[5][12][21] = xor_out[25][12][21] + xor_out[26][12][21] + xor_out[27][12][21] + xor_out[28][12][21] + xor_out[29][12][21];
assign sum_out[6][12][21] = xor_out[30][12][21] + xor_out[31][12][21] + xor_out[32][12][21] + xor_out[33][12][21] + xor_out[34][12][21];
assign sum_out[7][12][21] = xor_out[35][12][21] + xor_out[36][12][21] + xor_out[37][12][21] + xor_out[38][12][21] + xor_out[39][12][21];
assign sum_out[8][12][21] = xor_out[40][12][21] + xor_out[41][12][21] + xor_out[42][12][21] + xor_out[43][12][21] + xor_out[44][12][21];
assign sum_out[9][12][21] = xor_out[45][12][21] + xor_out[46][12][21] + xor_out[47][12][21] + xor_out[48][12][21] + xor_out[49][12][21];
assign sum_out[10][12][21] = xor_out[50][12][21] + xor_out[51][12][21] + xor_out[52][12][21] + xor_out[53][12][21] + xor_out[54][12][21];
assign sum_out[11][12][21] = xor_out[55][12][21] + xor_out[56][12][21] + xor_out[57][12][21] + xor_out[58][12][21] + xor_out[59][12][21];
assign sum_out[12][12][21] = xor_out[60][12][21] + xor_out[61][12][21] + xor_out[62][12][21] + xor_out[63][12][21] + xor_out[64][12][21];
assign sum_out[13][12][21] = xor_out[65][12][21] + xor_out[66][12][21] + xor_out[67][12][21] + xor_out[68][12][21] + xor_out[69][12][21];
assign sum_out[14][12][21] = xor_out[70][12][21] + xor_out[71][12][21] + xor_out[72][12][21] + xor_out[73][12][21] + xor_out[74][12][21];
assign sum_out[15][12][21] = xor_out[75][12][21] + xor_out[76][12][21] + xor_out[77][12][21] + xor_out[78][12][21] + xor_out[79][12][21];
assign sum_out[16][12][21] = xor_out[80][12][21] + xor_out[81][12][21] + xor_out[82][12][21] + xor_out[83][12][21] + xor_out[84][12][21];
assign sum_out[17][12][21] = xor_out[85][12][21] + xor_out[86][12][21] + xor_out[87][12][21] + xor_out[88][12][21] + xor_out[89][12][21];
assign sum_out[18][12][21] = xor_out[90][12][21] + xor_out[91][12][21] + xor_out[92][12][21] + xor_out[93][12][21] + xor_out[94][12][21];
assign sum_out[19][12][21] = xor_out[95][12][21] + xor_out[96][12][21] + xor_out[97][12][21] + xor_out[98][12][21] + xor_out[99][12][21];

assign sum_out[0][12][22] = xor_out[0][12][22] + xor_out[1][12][22] + xor_out[2][12][22] + xor_out[3][12][22] + xor_out[4][12][22];
assign sum_out[1][12][22] = xor_out[5][12][22] + xor_out[6][12][22] + xor_out[7][12][22] + xor_out[8][12][22] + xor_out[9][12][22];
assign sum_out[2][12][22] = xor_out[10][12][22] + xor_out[11][12][22] + xor_out[12][12][22] + xor_out[13][12][22] + xor_out[14][12][22];
assign sum_out[3][12][22] = xor_out[15][12][22] + xor_out[16][12][22] + xor_out[17][12][22] + xor_out[18][12][22] + xor_out[19][12][22];
assign sum_out[4][12][22] = xor_out[20][12][22] + xor_out[21][12][22] + xor_out[22][12][22] + xor_out[23][12][22] + xor_out[24][12][22];
assign sum_out[5][12][22] = xor_out[25][12][22] + xor_out[26][12][22] + xor_out[27][12][22] + xor_out[28][12][22] + xor_out[29][12][22];
assign sum_out[6][12][22] = xor_out[30][12][22] + xor_out[31][12][22] + xor_out[32][12][22] + xor_out[33][12][22] + xor_out[34][12][22];
assign sum_out[7][12][22] = xor_out[35][12][22] + xor_out[36][12][22] + xor_out[37][12][22] + xor_out[38][12][22] + xor_out[39][12][22];
assign sum_out[8][12][22] = xor_out[40][12][22] + xor_out[41][12][22] + xor_out[42][12][22] + xor_out[43][12][22] + xor_out[44][12][22];
assign sum_out[9][12][22] = xor_out[45][12][22] + xor_out[46][12][22] + xor_out[47][12][22] + xor_out[48][12][22] + xor_out[49][12][22];
assign sum_out[10][12][22] = xor_out[50][12][22] + xor_out[51][12][22] + xor_out[52][12][22] + xor_out[53][12][22] + xor_out[54][12][22];
assign sum_out[11][12][22] = xor_out[55][12][22] + xor_out[56][12][22] + xor_out[57][12][22] + xor_out[58][12][22] + xor_out[59][12][22];
assign sum_out[12][12][22] = xor_out[60][12][22] + xor_out[61][12][22] + xor_out[62][12][22] + xor_out[63][12][22] + xor_out[64][12][22];
assign sum_out[13][12][22] = xor_out[65][12][22] + xor_out[66][12][22] + xor_out[67][12][22] + xor_out[68][12][22] + xor_out[69][12][22];
assign sum_out[14][12][22] = xor_out[70][12][22] + xor_out[71][12][22] + xor_out[72][12][22] + xor_out[73][12][22] + xor_out[74][12][22];
assign sum_out[15][12][22] = xor_out[75][12][22] + xor_out[76][12][22] + xor_out[77][12][22] + xor_out[78][12][22] + xor_out[79][12][22];
assign sum_out[16][12][22] = xor_out[80][12][22] + xor_out[81][12][22] + xor_out[82][12][22] + xor_out[83][12][22] + xor_out[84][12][22];
assign sum_out[17][12][22] = xor_out[85][12][22] + xor_out[86][12][22] + xor_out[87][12][22] + xor_out[88][12][22] + xor_out[89][12][22];
assign sum_out[18][12][22] = xor_out[90][12][22] + xor_out[91][12][22] + xor_out[92][12][22] + xor_out[93][12][22] + xor_out[94][12][22];
assign sum_out[19][12][22] = xor_out[95][12][22] + xor_out[96][12][22] + xor_out[97][12][22] + xor_out[98][12][22] + xor_out[99][12][22];

assign sum_out[0][12][23] = xor_out[0][12][23] + xor_out[1][12][23] + xor_out[2][12][23] + xor_out[3][12][23] + xor_out[4][12][23];
assign sum_out[1][12][23] = xor_out[5][12][23] + xor_out[6][12][23] + xor_out[7][12][23] + xor_out[8][12][23] + xor_out[9][12][23];
assign sum_out[2][12][23] = xor_out[10][12][23] + xor_out[11][12][23] + xor_out[12][12][23] + xor_out[13][12][23] + xor_out[14][12][23];
assign sum_out[3][12][23] = xor_out[15][12][23] + xor_out[16][12][23] + xor_out[17][12][23] + xor_out[18][12][23] + xor_out[19][12][23];
assign sum_out[4][12][23] = xor_out[20][12][23] + xor_out[21][12][23] + xor_out[22][12][23] + xor_out[23][12][23] + xor_out[24][12][23];
assign sum_out[5][12][23] = xor_out[25][12][23] + xor_out[26][12][23] + xor_out[27][12][23] + xor_out[28][12][23] + xor_out[29][12][23];
assign sum_out[6][12][23] = xor_out[30][12][23] + xor_out[31][12][23] + xor_out[32][12][23] + xor_out[33][12][23] + xor_out[34][12][23];
assign sum_out[7][12][23] = xor_out[35][12][23] + xor_out[36][12][23] + xor_out[37][12][23] + xor_out[38][12][23] + xor_out[39][12][23];
assign sum_out[8][12][23] = xor_out[40][12][23] + xor_out[41][12][23] + xor_out[42][12][23] + xor_out[43][12][23] + xor_out[44][12][23];
assign sum_out[9][12][23] = xor_out[45][12][23] + xor_out[46][12][23] + xor_out[47][12][23] + xor_out[48][12][23] + xor_out[49][12][23];
assign sum_out[10][12][23] = xor_out[50][12][23] + xor_out[51][12][23] + xor_out[52][12][23] + xor_out[53][12][23] + xor_out[54][12][23];
assign sum_out[11][12][23] = xor_out[55][12][23] + xor_out[56][12][23] + xor_out[57][12][23] + xor_out[58][12][23] + xor_out[59][12][23];
assign sum_out[12][12][23] = xor_out[60][12][23] + xor_out[61][12][23] + xor_out[62][12][23] + xor_out[63][12][23] + xor_out[64][12][23];
assign sum_out[13][12][23] = xor_out[65][12][23] + xor_out[66][12][23] + xor_out[67][12][23] + xor_out[68][12][23] + xor_out[69][12][23];
assign sum_out[14][12][23] = xor_out[70][12][23] + xor_out[71][12][23] + xor_out[72][12][23] + xor_out[73][12][23] + xor_out[74][12][23];
assign sum_out[15][12][23] = xor_out[75][12][23] + xor_out[76][12][23] + xor_out[77][12][23] + xor_out[78][12][23] + xor_out[79][12][23];
assign sum_out[16][12][23] = xor_out[80][12][23] + xor_out[81][12][23] + xor_out[82][12][23] + xor_out[83][12][23] + xor_out[84][12][23];
assign sum_out[17][12][23] = xor_out[85][12][23] + xor_out[86][12][23] + xor_out[87][12][23] + xor_out[88][12][23] + xor_out[89][12][23];
assign sum_out[18][12][23] = xor_out[90][12][23] + xor_out[91][12][23] + xor_out[92][12][23] + xor_out[93][12][23] + xor_out[94][12][23];
assign sum_out[19][12][23] = xor_out[95][12][23] + xor_out[96][12][23] + xor_out[97][12][23] + xor_out[98][12][23] + xor_out[99][12][23];

assign sum_out[0][13][0] = xor_out[0][13][0] + xor_out[1][13][0] + xor_out[2][13][0] + xor_out[3][13][0] + xor_out[4][13][0];
assign sum_out[1][13][0] = xor_out[5][13][0] + xor_out[6][13][0] + xor_out[7][13][0] + xor_out[8][13][0] + xor_out[9][13][0];
assign sum_out[2][13][0] = xor_out[10][13][0] + xor_out[11][13][0] + xor_out[12][13][0] + xor_out[13][13][0] + xor_out[14][13][0];
assign sum_out[3][13][0] = xor_out[15][13][0] + xor_out[16][13][0] + xor_out[17][13][0] + xor_out[18][13][0] + xor_out[19][13][0];
assign sum_out[4][13][0] = xor_out[20][13][0] + xor_out[21][13][0] + xor_out[22][13][0] + xor_out[23][13][0] + xor_out[24][13][0];
assign sum_out[5][13][0] = xor_out[25][13][0] + xor_out[26][13][0] + xor_out[27][13][0] + xor_out[28][13][0] + xor_out[29][13][0];
assign sum_out[6][13][0] = xor_out[30][13][0] + xor_out[31][13][0] + xor_out[32][13][0] + xor_out[33][13][0] + xor_out[34][13][0];
assign sum_out[7][13][0] = xor_out[35][13][0] + xor_out[36][13][0] + xor_out[37][13][0] + xor_out[38][13][0] + xor_out[39][13][0];
assign sum_out[8][13][0] = xor_out[40][13][0] + xor_out[41][13][0] + xor_out[42][13][0] + xor_out[43][13][0] + xor_out[44][13][0];
assign sum_out[9][13][0] = xor_out[45][13][0] + xor_out[46][13][0] + xor_out[47][13][0] + xor_out[48][13][0] + xor_out[49][13][0];
assign sum_out[10][13][0] = xor_out[50][13][0] + xor_out[51][13][0] + xor_out[52][13][0] + xor_out[53][13][0] + xor_out[54][13][0];
assign sum_out[11][13][0] = xor_out[55][13][0] + xor_out[56][13][0] + xor_out[57][13][0] + xor_out[58][13][0] + xor_out[59][13][0];
assign sum_out[12][13][0] = xor_out[60][13][0] + xor_out[61][13][0] + xor_out[62][13][0] + xor_out[63][13][0] + xor_out[64][13][0];
assign sum_out[13][13][0] = xor_out[65][13][0] + xor_out[66][13][0] + xor_out[67][13][0] + xor_out[68][13][0] + xor_out[69][13][0];
assign sum_out[14][13][0] = xor_out[70][13][0] + xor_out[71][13][0] + xor_out[72][13][0] + xor_out[73][13][0] + xor_out[74][13][0];
assign sum_out[15][13][0] = xor_out[75][13][0] + xor_out[76][13][0] + xor_out[77][13][0] + xor_out[78][13][0] + xor_out[79][13][0];
assign sum_out[16][13][0] = xor_out[80][13][0] + xor_out[81][13][0] + xor_out[82][13][0] + xor_out[83][13][0] + xor_out[84][13][0];
assign sum_out[17][13][0] = xor_out[85][13][0] + xor_out[86][13][0] + xor_out[87][13][0] + xor_out[88][13][0] + xor_out[89][13][0];
assign sum_out[18][13][0] = xor_out[90][13][0] + xor_out[91][13][0] + xor_out[92][13][0] + xor_out[93][13][0] + xor_out[94][13][0];
assign sum_out[19][13][0] = xor_out[95][13][0] + xor_out[96][13][0] + xor_out[97][13][0] + xor_out[98][13][0] + xor_out[99][13][0];

assign sum_out[0][13][1] = xor_out[0][13][1] + xor_out[1][13][1] + xor_out[2][13][1] + xor_out[3][13][1] + xor_out[4][13][1];
assign sum_out[1][13][1] = xor_out[5][13][1] + xor_out[6][13][1] + xor_out[7][13][1] + xor_out[8][13][1] + xor_out[9][13][1];
assign sum_out[2][13][1] = xor_out[10][13][1] + xor_out[11][13][1] + xor_out[12][13][1] + xor_out[13][13][1] + xor_out[14][13][1];
assign sum_out[3][13][1] = xor_out[15][13][1] + xor_out[16][13][1] + xor_out[17][13][1] + xor_out[18][13][1] + xor_out[19][13][1];
assign sum_out[4][13][1] = xor_out[20][13][1] + xor_out[21][13][1] + xor_out[22][13][1] + xor_out[23][13][1] + xor_out[24][13][1];
assign sum_out[5][13][1] = xor_out[25][13][1] + xor_out[26][13][1] + xor_out[27][13][1] + xor_out[28][13][1] + xor_out[29][13][1];
assign sum_out[6][13][1] = xor_out[30][13][1] + xor_out[31][13][1] + xor_out[32][13][1] + xor_out[33][13][1] + xor_out[34][13][1];
assign sum_out[7][13][1] = xor_out[35][13][1] + xor_out[36][13][1] + xor_out[37][13][1] + xor_out[38][13][1] + xor_out[39][13][1];
assign sum_out[8][13][1] = xor_out[40][13][1] + xor_out[41][13][1] + xor_out[42][13][1] + xor_out[43][13][1] + xor_out[44][13][1];
assign sum_out[9][13][1] = xor_out[45][13][1] + xor_out[46][13][1] + xor_out[47][13][1] + xor_out[48][13][1] + xor_out[49][13][1];
assign sum_out[10][13][1] = xor_out[50][13][1] + xor_out[51][13][1] + xor_out[52][13][1] + xor_out[53][13][1] + xor_out[54][13][1];
assign sum_out[11][13][1] = xor_out[55][13][1] + xor_out[56][13][1] + xor_out[57][13][1] + xor_out[58][13][1] + xor_out[59][13][1];
assign sum_out[12][13][1] = xor_out[60][13][1] + xor_out[61][13][1] + xor_out[62][13][1] + xor_out[63][13][1] + xor_out[64][13][1];
assign sum_out[13][13][1] = xor_out[65][13][1] + xor_out[66][13][1] + xor_out[67][13][1] + xor_out[68][13][1] + xor_out[69][13][1];
assign sum_out[14][13][1] = xor_out[70][13][1] + xor_out[71][13][1] + xor_out[72][13][1] + xor_out[73][13][1] + xor_out[74][13][1];
assign sum_out[15][13][1] = xor_out[75][13][1] + xor_out[76][13][1] + xor_out[77][13][1] + xor_out[78][13][1] + xor_out[79][13][1];
assign sum_out[16][13][1] = xor_out[80][13][1] + xor_out[81][13][1] + xor_out[82][13][1] + xor_out[83][13][1] + xor_out[84][13][1];
assign sum_out[17][13][1] = xor_out[85][13][1] + xor_out[86][13][1] + xor_out[87][13][1] + xor_out[88][13][1] + xor_out[89][13][1];
assign sum_out[18][13][1] = xor_out[90][13][1] + xor_out[91][13][1] + xor_out[92][13][1] + xor_out[93][13][1] + xor_out[94][13][1];
assign sum_out[19][13][1] = xor_out[95][13][1] + xor_out[96][13][1] + xor_out[97][13][1] + xor_out[98][13][1] + xor_out[99][13][1];

assign sum_out[0][13][2] = xor_out[0][13][2] + xor_out[1][13][2] + xor_out[2][13][2] + xor_out[3][13][2] + xor_out[4][13][2];
assign sum_out[1][13][2] = xor_out[5][13][2] + xor_out[6][13][2] + xor_out[7][13][2] + xor_out[8][13][2] + xor_out[9][13][2];
assign sum_out[2][13][2] = xor_out[10][13][2] + xor_out[11][13][2] + xor_out[12][13][2] + xor_out[13][13][2] + xor_out[14][13][2];
assign sum_out[3][13][2] = xor_out[15][13][2] + xor_out[16][13][2] + xor_out[17][13][2] + xor_out[18][13][2] + xor_out[19][13][2];
assign sum_out[4][13][2] = xor_out[20][13][2] + xor_out[21][13][2] + xor_out[22][13][2] + xor_out[23][13][2] + xor_out[24][13][2];
assign sum_out[5][13][2] = xor_out[25][13][2] + xor_out[26][13][2] + xor_out[27][13][2] + xor_out[28][13][2] + xor_out[29][13][2];
assign sum_out[6][13][2] = xor_out[30][13][2] + xor_out[31][13][2] + xor_out[32][13][2] + xor_out[33][13][2] + xor_out[34][13][2];
assign sum_out[7][13][2] = xor_out[35][13][2] + xor_out[36][13][2] + xor_out[37][13][2] + xor_out[38][13][2] + xor_out[39][13][2];
assign sum_out[8][13][2] = xor_out[40][13][2] + xor_out[41][13][2] + xor_out[42][13][2] + xor_out[43][13][2] + xor_out[44][13][2];
assign sum_out[9][13][2] = xor_out[45][13][2] + xor_out[46][13][2] + xor_out[47][13][2] + xor_out[48][13][2] + xor_out[49][13][2];
assign sum_out[10][13][2] = xor_out[50][13][2] + xor_out[51][13][2] + xor_out[52][13][2] + xor_out[53][13][2] + xor_out[54][13][2];
assign sum_out[11][13][2] = xor_out[55][13][2] + xor_out[56][13][2] + xor_out[57][13][2] + xor_out[58][13][2] + xor_out[59][13][2];
assign sum_out[12][13][2] = xor_out[60][13][2] + xor_out[61][13][2] + xor_out[62][13][2] + xor_out[63][13][2] + xor_out[64][13][2];
assign sum_out[13][13][2] = xor_out[65][13][2] + xor_out[66][13][2] + xor_out[67][13][2] + xor_out[68][13][2] + xor_out[69][13][2];
assign sum_out[14][13][2] = xor_out[70][13][2] + xor_out[71][13][2] + xor_out[72][13][2] + xor_out[73][13][2] + xor_out[74][13][2];
assign sum_out[15][13][2] = xor_out[75][13][2] + xor_out[76][13][2] + xor_out[77][13][2] + xor_out[78][13][2] + xor_out[79][13][2];
assign sum_out[16][13][2] = xor_out[80][13][2] + xor_out[81][13][2] + xor_out[82][13][2] + xor_out[83][13][2] + xor_out[84][13][2];
assign sum_out[17][13][2] = xor_out[85][13][2] + xor_out[86][13][2] + xor_out[87][13][2] + xor_out[88][13][2] + xor_out[89][13][2];
assign sum_out[18][13][2] = xor_out[90][13][2] + xor_out[91][13][2] + xor_out[92][13][2] + xor_out[93][13][2] + xor_out[94][13][2];
assign sum_out[19][13][2] = xor_out[95][13][2] + xor_out[96][13][2] + xor_out[97][13][2] + xor_out[98][13][2] + xor_out[99][13][2];

assign sum_out[0][13][3] = xor_out[0][13][3] + xor_out[1][13][3] + xor_out[2][13][3] + xor_out[3][13][3] + xor_out[4][13][3];
assign sum_out[1][13][3] = xor_out[5][13][3] + xor_out[6][13][3] + xor_out[7][13][3] + xor_out[8][13][3] + xor_out[9][13][3];
assign sum_out[2][13][3] = xor_out[10][13][3] + xor_out[11][13][3] + xor_out[12][13][3] + xor_out[13][13][3] + xor_out[14][13][3];
assign sum_out[3][13][3] = xor_out[15][13][3] + xor_out[16][13][3] + xor_out[17][13][3] + xor_out[18][13][3] + xor_out[19][13][3];
assign sum_out[4][13][3] = xor_out[20][13][3] + xor_out[21][13][3] + xor_out[22][13][3] + xor_out[23][13][3] + xor_out[24][13][3];
assign sum_out[5][13][3] = xor_out[25][13][3] + xor_out[26][13][3] + xor_out[27][13][3] + xor_out[28][13][3] + xor_out[29][13][3];
assign sum_out[6][13][3] = xor_out[30][13][3] + xor_out[31][13][3] + xor_out[32][13][3] + xor_out[33][13][3] + xor_out[34][13][3];
assign sum_out[7][13][3] = xor_out[35][13][3] + xor_out[36][13][3] + xor_out[37][13][3] + xor_out[38][13][3] + xor_out[39][13][3];
assign sum_out[8][13][3] = xor_out[40][13][3] + xor_out[41][13][3] + xor_out[42][13][3] + xor_out[43][13][3] + xor_out[44][13][3];
assign sum_out[9][13][3] = xor_out[45][13][3] + xor_out[46][13][3] + xor_out[47][13][3] + xor_out[48][13][3] + xor_out[49][13][3];
assign sum_out[10][13][3] = xor_out[50][13][3] + xor_out[51][13][3] + xor_out[52][13][3] + xor_out[53][13][3] + xor_out[54][13][3];
assign sum_out[11][13][3] = xor_out[55][13][3] + xor_out[56][13][3] + xor_out[57][13][3] + xor_out[58][13][3] + xor_out[59][13][3];
assign sum_out[12][13][3] = xor_out[60][13][3] + xor_out[61][13][3] + xor_out[62][13][3] + xor_out[63][13][3] + xor_out[64][13][3];
assign sum_out[13][13][3] = xor_out[65][13][3] + xor_out[66][13][3] + xor_out[67][13][3] + xor_out[68][13][3] + xor_out[69][13][3];
assign sum_out[14][13][3] = xor_out[70][13][3] + xor_out[71][13][3] + xor_out[72][13][3] + xor_out[73][13][3] + xor_out[74][13][3];
assign sum_out[15][13][3] = xor_out[75][13][3] + xor_out[76][13][3] + xor_out[77][13][3] + xor_out[78][13][3] + xor_out[79][13][3];
assign sum_out[16][13][3] = xor_out[80][13][3] + xor_out[81][13][3] + xor_out[82][13][3] + xor_out[83][13][3] + xor_out[84][13][3];
assign sum_out[17][13][3] = xor_out[85][13][3] + xor_out[86][13][3] + xor_out[87][13][3] + xor_out[88][13][3] + xor_out[89][13][3];
assign sum_out[18][13][3] = xor_out[90][13][3] + xor_out[91][13][3] + xor_out[92][13][3] + xor_out[93][13][3] + xor_out[94][13][3];
assign sum_out[19][13][3] = xor_out[95][13][3] + xor_out[96][13][3] + xor_out[97][13][3] + xor_out[98][13][3] + xor_out[99][13][3];

assign sum_out[0][13][4] = xor_out[0][13][4] + xor_out[1][13][4] + xor_out[2][13][4] + xor_out[3][13][4] + xor_out[4][13][4];
assign sum_out[1][13][4] = xor_out[5][13][4] + xor_out[6][13][4] + xor_out[7][13][4] + xor_out[8][13][4] + xor_out[9][13][4];
assign sum_out[2][13][4] = xor_out[10][13][4] + xor_out[11][13][4] + xor_out[12][13][4] + xor_out[13][13][4] + xor_out[14][13][4];
assign sum_out[3][13][4] = xor_out[15][13][4] + xor_out[16][13][4] + xor_out[17][13][4] + xor_out[18][13][4] + xor_out[19][13][4];
assign sum_out[4][13][4] = xor_out[20][13][4] + xor_out[21][13][4] + xor_out[22][13][4] + xor_out[23][13][4] + xor_out[24][13][4];
assign sum_out[5][13][4] = xor_out[25][13][4] + xor_out[26][13][4] + xor_out[27][13][4] + xor_out[28][13][4] + xor_out[29][13][4];
assign sum_out[6][13][4] = xor_out[30][13][4] + xor_out[31][13][4] + xor_out[32][13][4] + xor_out[33][13][4] + xor_out[34][13][4];
assign sum_out[7][13][4] = xor_out[35][13][4] + xor_out[36][13][4] + xor_out[37][13][4] + xor_out[38][13][4] + xor_out[39][13][4];
assign sum_out[8][13][4] = xor_out[40][13][4] + xor_out[41][13][4] + xor_out[42][13][4] + xor_out[43][13][4] + xor_out[44][13][4];
assign sum_out[9][13][4] = xor_out[45][13][4] + xor_out[46][13][4] + xor_out[47][13][4] + xor_out[48][13][4] + xor_out[49][13][4];
assign sum_out[10][13][4] = xor_out[50][13][4] + xor_out[51][13][4] + xor_out[52][13][4] + xor_out[53][13][4] + xor_out[54][13][4];
assign sum_out[11][13][4] = xor_out[55][13][4] + xor_out[56][13][4] + xor_out[57][13][4] + xor_out[58][13][4] + xor_out[59][13][4];
assign sum_out[12][13][4] = xor_out[60][13][4] + xor_out[61][13][4] + xor_out[62][13][4] + xor_out[63][13][4] + xor_out[64][13][4];
assign sum_out[13][13][4] = xor_out[65][13][4] + xor_out[66][13][4] + xor_out[67][13][4] + xor_out[68][13][4] + xor_out[69][13][4];
assign sum_out[14][13][4] = xor_out[70][13][4] + xor_out[71][13][4] + xor_out[72][13][4] + xor_out[73][13][4] + xor_out[74][13][4];
assign sum_out[15][13][4] = xor_out[75][13][4] + xor_out[76][13][4] + xor_out[77][13][4] + xor_out[78][13][4] + xor_out[79][13][4];
assign sum_out[16][13][4] = xor_out[80][13][4] + xor_out[81][13][4] + xor_out[82][13][4] + xor_out[83][13][4] + xor_out[84][13][4];
assign sum_out[17][13][4] = xor_out[85][13][4] + xor_out[86][13][4] + xor_out[87][13][4] + xor_out[88][13][4] + xor_out[89][13][4];
assign sum_out[18][13][4] = xor_out[90][13][4] + xor_out[91][13][4] + xor_out[92][13][4] + xor_out[93][13][4] + xor_out[94][13][4];
assign sum_out[19][13][4] = xor_out[95][13][4] + xor_out[96][13][4] + xor_out[97][13][4] + xor_out[98][13][4] + xor_out[99][13][4];

assign sum_out[0][13][5] = xor_out[0][13][5] + xor_out[1][13][5] + xor_out[2][13][5] + xor_out[3][13][5] + xor_out[4][13][5];
assign sum_out[1][13][5] = xor_out[5][13][5] + xor_out[6][13][5] + xor_out[7][13][5] + xor_out[8][13][5] + xor_out[9][13][5];
assign sum_out[2][13][5] = xor_out[10][13][5] + xor_out[11][13][5] + xor_out[12][13][5] + xor_out[13][13][5] + xor_out[14][13][5];
assign sum_out[3][13][5] = xor_out[15][13][5] + xor_out[16][13][5] + xor_out[17][13][5] + xor_out[18][13][5] + xor_out[19][13][5];
assign sum_out[4][13][5] = xor_out[20][13][5] + xor_out[21][13][5] + xor_out[22][13][5] + xor_out[23][13][5] + xor_out[24][13][5];
assign sum_out[5][13][5] = xor_out[25][13][5] + xor_out[26][13][5] + xor_out[27][13][5] + xor_out[28][13][5] + xor_out[29][13][5];
assign sum_out[6][13][5] = xor_out[30][13][5] + xor_out[31][13][5] + xor_out[32][13][5] + xor_out[33][13][5] + xor_out[34][13][5];
assign sum_out[7][13][5] = xor_out[35][13][5] + xor_out[36][13][5] + xor_out[37][13][5] + xor_out[38][13][5] + xor_out[39][13][5];
assign sum_out[8][13][5] = xor_out[40][13][5] + xor_out[41][13][5] + xor_out[42][13][5] + xor_out[43][13][5] + xor_out[44][13][5];
assign sum_out[9][13][5] = xor_out[45][13][5] + xor_out[46][13][5] + xor_out[47][13][5] + xor_out[48][13][5] + xor_out[49][13][5];
assign sum_out[10][13][5] = xor_out[50][13][5] + xor_out[51][13][5] + xor_out[52][13][5] + xor_out[53][13][5] + xor_out[54][13][5];
assign sum_out[11][13][5] = xor_out[55][13][5] + xor_out[56][13][5] + xor_out[57][13][5] + xor_out[58][13][5] + xor_out[59][13][5];
assign sum_out[12][13][5] = xor_out[60][13][5] + xor_out[61][13][5] + xor_out[62][13][5] + xor_out[63][13][5] + xor_out[64][13][5];
assign sum_out[13][13][5] = xor_out[65][13][5] + xor_out[66][13][5] + xor_out[67][13][5] + xor_out[68][13][5] + xor_out[69][13][5];
assign sum_out[14][13][5] = xor_out[70][13][5] + xor_out[71][13][5] + xor_out[72][13][5] + xor_out[73][13][5] + xor_out[74][13][5];
assign sum_out[15][13][5] = xor_out[75][13][5] + xor_out[76][13][5] + xor_out[77][13][5] + xor_out[78][13][5] + xor_out[79][13][5];
assign sum_out[16][13][5] = xor_out[80][13][5] + xor_out[81][13][5] + xor_out[82][13][5] + xor_out[83][13][5] + xor_out[84][13][5];
assign sum_out[17][13][5] = xor_out[85][13][5] + xor_out[86][13][5] + xor_out[87][13][5] + xor_out[88][13][5] + xor_out[89][13][5];
assign sum_out[18][13][5] = xor_out[90][13][5] + xor_out[91][13][5] + xor_out[92][13][5] + xor_out[93][13][5] + xor_out[94][13][5];
assign sum_out[19][13][5] = xor_out[95][13][5] + xor_out[96][13][5] + xor_out[97][13][5] + xor_out[98][13][5] + xor_out[99][13][5];

assign sum_out[0][13][6] = xor_out[0][13][6] + xor_out[1][13][6] + xor_out[2][13][6] + xor_out[3][13][6] + xor_out[4][13][6];
assign sum_out[1][13][6] = xor_out[5][13][6] + xor_out[6][13][6] + xor_out[7][13][6] + xor_out[8][13][6] + xor_out[9][13][6];
assign sum_out[2][13][6] = xor_out[10][13][6] + xor_out[11][13][6] + xor_out[12][13][6] + xor_out[13][13][6] + xor_out[14][13][6];
assign sum_out[3][13][6] = xor_out[15][13][6] + xor_out[16][13][6] + xor_out[17][13][6] + xor_out[18][13][6] + xor_out[19][13][6];
assign sum_out[4][13][6] = xor_out[20][13][6] + xor_out[21][13][6] + xor_out[22][13][6] + xor_out[23][13][6] + xor_out[24][13][6];
assign sum_out[5][13][6] = xor_out[25][13][6] + xor_out[26][13][6] + xor_out[27][13][6] + xor_out[28][13][6] + xor_out[29][13][6];
assign sum_out[6][13][6] = xor_out[30][13][6] + xor_out[31][13][6] + xor_out[32][13][6] + xor_out[33][13][6] + xor_out[34][13][6];
assign sum_out[7][13][6] = xor_out[35][13][6] + xor_out[36][13][6] + xor_out[37][13][6] + xor_out[38][13][6] + xor_out[39][13][6];
assign sum_out[8][13][6] = xor_out[40][13][6] + xor_out[41][13][6] + xor_out[42][13][6] + xor_out[43][13][6] + xor_out[44][13][6];
assign sum_out[9][13][6] = xor_out[45][13][6] + xor_out[46][13][6] + xor_out[47][13][6] + xor_out[48][13][6] + xor_out[49][13][6];
assign sum_out[10][13][6] = xor_out[50][13][6] + xor_out[51][13][6] + xor_out[52][13][6] + xor_out[53][13][6] + xor_out[54][13][6];
assign sum_out[11][13][6] = xor_out[55][13][6] + xor_out[56][13][6] + xor_out[57][13][6] + xor_out[58][13][6] + xor_out[59][13][6];
assign sum_out[12][13][6] = xor_out[60][13][6] + xor_out[61][13][6] + xor_out[62][13][6] + xor_out[63][13][6] + xor_out[64][13][6];
assign sum_out[13][13][6] = xor_out[65][13][6] + xor_out[66][13][6] + xor_out[67][13][6] + xor_out[68][13][6] + xor_out[69][13][6];
assign sum_out[14][13][6] = xor_out[70][13][6] + xor_out[71][13][6] + xor_out[72][13][6] + xor_out[73][13][6] + xor_out[74][13][6];
assign sum_out[15][13][6] = xor_out[75][13][6] + xor_out[76][13][6] + xor_out[77][13][6] + xor_out[78][13][6] + xor_out[79][13][6];
assign sum_out[16][13][6] = xor_out[80][13][6] + xor_out[81][13][6] + xor_out[82][13][6] + xor_out[83][13][6] + xor_out[84][13][6];
assign sum_out[17][13][6] = xor_out[85][13][6] + xor_out[86][13][6] + xor_out[87][13][6] + xor_out[88][13][6] + xor_out[89][13][6];
assign sum_out[18][13][6] = xor_out[90][13][6] + xor_out[91][13][6] + xor_out[92][13][6] + xor_out[93][13][6] + xor_out[94][13][6];
assign sum_out[19][13][6] = xor_out[95][13][6] + xor_out[96][13][6] + xor_out[97][13][6] + xor_out[98][13][6] + xor_out[99][13][6];

assign sum_out[0][13][7] = xor_out[0][13][7] + xor_out[1][13][7] + xor_out[2][13][7] + xor_out[3][13][7] + xor_out[4][13][7];
assign sum_out[1][13][7] = xor_out[5][13][7] + xor_out[6][13][7] + xor_out[7][13][7] + xor_out[8][13][7] + xor_out[9][13][7];
assign sum_out[2][13][7] = xor_out[10][13][7] + xor_out[11][13][7] + xor_out[12][13][7] + xor_out[13][13][7] + xor_out[14][13][7];
assign sum_out[3][13][7] = xor_out[15][13][7] + xor_out[16][13][7] + xor_out[17][13][7] + xor_out[18][13][7] + xor_out[19][13][7];
assign sum_out[4][13][7] = xor_out[20][13][7] + xor_out[21][13][7] + xor_out[22][13][7] + xor_out[23][13][7] + xor_out[24][13][7];
assign sum_out[5][13][7] = xor_out[25][13][7] + xor_out[26][13][7] + xor_out[27][13][7] + xor_out[28][13][7] + xor_out[29][13][7];
assign sum_out[6][13][7] = xor_out[30][13][7] + xor_out[31][13][7] + xor_out[32][13][7] + xor_out[33][13][7] + xor_out[34][13][7];
assign sum_out[7][13][7] = xor_out[35][13][7] + xor_out[36][13][7] + xor_out[37][13][7] + xor_out[38][13][7] + xor_out[39][13][7];
assign sum_out[8][13][7] = xor_out[40][13][7] + xor_out[41][13][7] + xor_out[42][13][7] + xor_out[43][13][7] + xor_out[44][13][7];
assign sum_out[9][13][7] = xor_out[45][13][7] + xor_out[46][13][7] + xor_out[47][13][7] + xor_out[48][13][7] + xor_out[49][13][7];
assign sum_out[10][13][7] = xor_out[50][13][7] + xor_out[51][13][7] + xor_out[52][13][7] + xor_out[53][13][7] + xor_out[54][13][7];
assign sum_out[11][13][7] = xor_out[55][13][7] + xor_out[56][13][7] + xor_out[57][13][7] + xor_out[58][13][7] + xor_out[59][13][7];
assign sum_out[12][13][7] = xor_out[60][13][7] + xor_out[61][13][7] + xor_out[62][13][7] + xor_out[63][13][7] + xor_out[64][13][7];
assign sum_out[13][13][7] = xor_out[65][13][7] + xor_out[66][13][7] + xor_out[67][13][7] + xor_out[68][13][7] + xor_out[69][13][7];
assign sum_out[14][13][7] = xor_out[70][13][7] + xor_out[71][13][7] + xor_out[72][13][7] + xor_out[73][13][7] + xor_out[74][13][7];
assign sum_out[15][13][7] = xor_out[75][13][7] + xor_out[76][13][7] + xor_out[77][13][7] + xor_out[78][13][7] + xor_out[79][13][7];
assign sum_out[16][13][7] = xor_out[80][13][7] + xor_out[81][13][7] + xor_out[82][13][7] + xor_out[83][13][7] + xor_out[84][13][7];
assign sum_out[17][13][7] = xor_out[85][13][7] + xor_out[86][13][7] + xor_out[87][13][7] + xor_out[88][13][7] + xor_out[89][13][7];
assign sum_out[18][13][7] = xor_out[90][13][7] + xor_out[91][13][7] + xor_out[92][13][7] + xor_out[93][13][7] + xor_out[94][13][7];
assign sum_out[19][13][7] = xor_out[95][13][7] + xor_out[96][13][7] + xor_out[97][13][7] + xor_out[98][13][7] + xor_out[99][13][7];

assign sum_out[0][13][8] = xor_out[0][13][8] + xor_out[1][13][8] + xor_out[2][13][8] + xor_out[3][13][8] + xor_out[4][13][8];
assign sum_out[1][13][8] = xor_out[5][13][8] + xor_out[6][13][8] + xor_out[7][13][8] + xor_out[8][13][8] + xor_out[9][13][8];
assign sum_out[2][13][8] = xor_out[10][13][8] + xor_out[11][13][8] + xor_out[12][13][8] + xor_out[13][13][8] + xor_out[14][13][8];
assign sum_out[3][13][8] = xor_out[15][13][8] + xor_out[16][13][8] + xor_out[17][13][8] + xor_out[18][13][8] + xor_out[19][13][8];
assign sum_out[4][13][8] = xor_out[20][13][8] + xor_out[21][13][8] + xor_out[22][13][8] + xor_out[23][13][8] + xor_out[24][13][8];
assign sum_out[5][13][8] = xor_out[25][13][8] + xor_out[26][13][8] + xor_out[27][13][8] + xor_out[28][13][8] + xor_out[29][13][8];
assign sum_out[6][13][8] = xor_out[30][13][8] + xor_out[31][13][8] + xor_out[32][13][8] + xor_out[33][13][8] + xor_out[34][13][8];
assign sum_out[7][13][8] = xor_out[35][13][8] + xor_out[36][13][8] + xor_out[37][13][8] + xor_out[38][13][8] + xor_out[39][13][8];
assign sum_out[8][13][8] = xor_out[40][13][8] + xor_out[41][13][8] + xor_out[42][13][8] + xor_out[43][13][8] + xor_out[44][13][8];
assign sum_out[9][13][8] = xor_out[45][13][8] + xor_out[46][13][8] + xor_out[47][13][8] + xor_out[48][13][8] + xor_out[49][13][8];
assign sum_out[10][13][8] = xor_out[50][13][8] + xor_out[51][13][8] + xor_out[52][13][8] + xor_out[53][13][8] + xor_out[54][13][8];
assign sum_out[11][13][8] = xor_out[55][13][8] + xor_out[56][13][8] + xor_out[57][13][8] + xor_out[58][13][8] + xor_out[59][13][8];
assign sum_out[12][13][8] = xor_out[60][13][8] + xor_out[61][13][8] + xor_out[62][13][8] + xor_out[63][13][8] + xor_out[64][13][8];
assign sum_out[13][13][8] = xor_out[65][13][8] + xor_out[66][13][8] + xor_out[67][13][8] + xor_out[68][13][8] + xor_out[69][13][8];
assign sum_out[14][13][8] = xor_out[70][13][8] + xor_out[71][13][8] + xor_out[72][13][8] + xor_out[73][13][8] + xor_out[74][13][8];
assign sum_out[15][13][8] = xor_out[75][13][8] + xor_out[76][13][8] + xor_out[77][13][8] + xor_out[78][13][8] + xor_out[79][13][8];
assign sum_out[16][13][8] = xor_out[80][13][8] + xor_out[81][13][8] + xor_out[82][13][8] + xor_out[83][13][8] + xor_out[84][13][8];
assign sum_out[17][13][8] = xor_out[85][13][8] + xor_out[86][13][8] + xor_out[87][13][8] + xor_out[88][13][8] + xor_out[89][13][8];
assign sum_out[18][13][8] = xor_out[90][13][8] + xor_out[91][13][8] + xor_out[92][13][8] + xor_out[93][13][8] + xor_out[94][13][8];
assign sum_out[19][13][8] = xor_out[95][13][8] + xor_out[96][13][8] + xor_out[97][13][8] + xor_out[98][13][8] + xor_out[99][13][8];

assign sum_out[0][13][9] = xor_out[0][13][9] + xor_out[1][13][9] + xor_out[2][13][9] + xor_out[3][13][9] + xor_out[4][13][9];
assign sum_out[1][13][9] = xor_out[5][13][9] + xor_out[6][13][9] + xor_out[7][13][9] + xor_out[8][13][9] + xor_out[9][13][9];
assign sum_out[2][13][9] = xor_out[10][13][9] + xor_out[11][13][9] + xor_out[12][13][9] + xor_out[13][13][9] + xor_out[14][13][9];
assign sum_out[3][13][9] = xor_out[15][13][9] + xor_out[16][13][9] + xor_out[17][13][9] + xor_out[18][13][9] + xor_out[19][13][9];
assign sum_out[4][13][9] = xor_out[20][13][9] + xor_out[21][13][9] + xor_out[22][13][9] + xor_out[23][13][9] + xor_out[24][13][9];
assign sum_out[5][13][9] = xor_out[25][13][9] + xor_out[26][13][9] + xor_out[27][13][9] + xor_out[28][13][9] + xor_out[29][13][9];
assign sum_out[6][13][9] = xor_out[30][13][9] + xor_out[31][13][9] + xor_out[32][13][9] + xor_out[33][13][9] + xor_out[34][13][9];
assign sum_out[7][13][9] = xor_out[35][13][9] + xor_out[36][13][9] + xor_out[37][13][9] + xor_out[38][13][9] + xor_out[39][13][9];
assign sum_out[8][13][9] = xor_out[40][13][9] + xor_out[41][13][9] + xor_out[42][13][9] + xor_out[43][13][9] + xor_out[44][13][9];
assign sum_out[9][13][9] = xor_out[45][13][9] + xor_out[46][13][9] + xor_out[47][13][9] + xor_out[48][13][9] + xor_out[49][13][9];
assign sum_out[10][13][9] = xor_out[50][13][9] + xor_out[51][13][9] + xor_out[52][13][9] + xor_out[53][13][9] + xor_out[54][13][9];
assign sum_out[11][13][9] = xor_out[55][13][9] + xor_out[56][13][9] + xor_out[57][13][9] + xor_out[58][13][9] + xor_out[59][13][9];
assign sum_out[12][13][9] = xor_out[60][13][9] + xor_out[61][13][9] + xor_out[62][13][9] + xor_out[63][13][9] + xor_out[64][13][9];
assign sum_out[13][13][9] = xor_out[65][13][9] + xor_out[66][13][9] + xor_out[67][13][9] + xor_out[68][13][9] + xor_out[69][13][9];
assign sum_out[14][13][9] = xor_out[70][13][9] + xor_out[71][13][9] + xor_out[72][13][9] + xor_out[73][13][9] + xor_out[74][13][9];
assign sum_out[15][13][9] = xor_out[75][13][9] + xor_out[76][13][9] + xor_out[77][13][9] + xor_out[78][13][9] + xor_out[79][13][9];
assign sum_out[16][13][9] = xor_out[80][13][9] + xor_out[81][13][9] + xor_out[82][13][9] + xor_out[83][13][9] + xor_out[84][13][9];
assign sum_out[17][13][9] = xor_out[85][13][9] + xor_out[86][13][9] + xor_out[87][13][9] + xor_out[88][13][9] + xor_out[89][13][9];
assign sum_out[18][13][9] = xor_out[90][13][9] + xor_out[91][13][9] + xor_out[92][13][9] + xor_out[93][13][9] + xor_out[94][13][9];
assign sum_out[19][13][9] = xor_out[95][13][9] + xor_out[96][13][9] + xor_out[97][13][9] + xor_out[98][13][9] + xor_out[99][13][9];

assign sum_out[0][13][10] = xor_out[0][13][10] + xor_out[1][13][10] + xor_out[2][13][10] + xor_out[3][13][10] + xor_out[4][13][10];
assign sum_out[1][13][10] = xor_out[5][13][10] + xor_out[6][13][10] + xor_out[7][13][10] + xor_out[8][13][10] + xor_out[9][13][10];
assign sum_out[2][13][10] = xor_out[10][13][10] + xor_out[11][13][10] + xor_out[12][13][10] + xor_out[13][13][10] + xor_out[14][13][10];
assign sum_out[3][13][10] = xor_out[15][13][10] + xor_out[16][13][10] + xor_out[17][13][10] + xor_out[18][13][10] + xor_out[19][13][10];
assign sum_out[4][13][10] = xor_out[20][13][10] + xor_out[21][13][10] + xor_out[22][13][10] + xor_out[23][13][10] + xor_out[24][13][10];
assign sum_out[5][13][10] = xor_out[25][13][10] + xor_out[26][13][10] + xor_out[27][13][10] + xor_out[28][13][10] + xor_out[29][13][10];
assign sum_out[6][13][10] = xor_out[30][13][10] + xor_out[31][13][10] + xor_out[32][13][10] + xor_out[33][13][10] + xor_out[34][13][10];
assign sum_out[7][13][10] = xor_out[35][13][10] + xor_out[36][13][10] + xor_out[37][13][10] + xor_out[38][13][10] + xor_out[39][13][10];
assign sum_out[8][13][10] = xor_out[40][13][10] + xor_out[41][13][10] + xor_out[42][13][10] + xor_out[43][13][10] + xor_out[44][13][10];
assign sum_out[9][13][10] = xor_out[45][13][10] + xor_out[46][13][10] + xor_out[47][13][10] + xor_out[48][13][10] + xor_out[49][13][10];
assign sum_out[10][13][10] = xor_out[50][13][10] + xor_out[51][13][10] + xor_out[52][13][10] + xor_out[53][13][10] + xor_out[54][13][10];
assign sum_out[11][13][10] = xor_out[55][13][10] + xor_out[56][13][10] + xor_out[57][13][10] + xor_out[58][13][10] + xor_out[59][13][10];
assign sum_out[12][13][10] = xor_out[60][13][10] + xor_out[61][13][10] + xor_out[62][13][10] + xor_out[63][13][10] + xor_out[64][13][10];
assign sum_out[13][13][10] = xor_out[65][13][10] + xor_out[66][13][10] + xor_out[67][13][10] + xor_out[68][13][10] + xor_out[69][13][10];
assign sum_out[14][13][10] = xor_out[70][13][10] + xor_out[71][13][10] + xor_out[72][13][10] + xor_out[73][13][10] + xor_out[74][13][10];
assign sum_out[15][13][10] = xor_out[75][13][10] + xor_out[76][13][10] + xor_out[77][13][10] + xor_out[78][13][10] + xor_out[79][13][10];
assign sum_out[16][13][10] = xor_out[80][13][10] + xor_out[81][13][10] + xor_out[82][13][10] + xor_out[83][13][10] + xor_out[84][13][10];
assign sum_out[17][13][10] = xor_out[85][13][10] + xor_out[86][13][10] + xor_out[87][13][10] + xor_out[88][13][10] + xor_out[89][13][10];
assign sum_out[18][13][10] = xor_out[90][13][10] + xor_out[91][13][10] + xor_out[92][13][10] + xor_out[93][13][10] + xor_out[94][13][10];
assign sum_out[19][13][10] = xor_out[95][13][10] + xor_out[96][13][10] + xor_out[97][13][10] + xor_out[98][13][10] + xor_out[99][13][10];

assign sum_out[0][13][11] = xor_out[0][13][11] + xor_out[1][13][11] + xor_out[2][13][11] + xor_out[3][13][11] + xor_out[4][13][11];
assign sum_out[1][13][11] = xor_out[5][13][11] + xor_out[6][13][11] + xor_out[7][13][11] + xor_out[8][13][11] + xor_out[9][13][11];
assign sum_out[2][13][11] = xor_out[10][13][11] + xor_out[11][13][11] + xor_out[12][13][11] + xor_out[13][13][11] + xor_out[14][13][11];
assign sum_out[3][13][11] = xor_out[15][13][11] + xor_out[16][13][11] + xor_out[17][13][11] + xor_out[18][13][11] + xor_out[19][13][11];
assign sum_out[4][13][11] = xor_out[20][13][11] + xor_out[21][13][11] + xor_out[22][13][11] + xor_out[23][13][11] + xor_out[24][13][11];
assign sum_out[5][13][11] = xor_out[25][13][11] + xor_out[26][13][11] + xor_out[27][13][11] + xor_out[28][13][11] + xor_out[29][13][11];
assign sum_out[6][13][11] = xor_out[30][13][11] + xor_out[31][13][11] + xor_out[32][13][11] + xor_out[33][13][11] + xor_out[34][13][11];
assign sum_out[7][13][11] = xor_out[35][13][11] + xor_out[36][13][11] + xor_out[37][13][11] + xor_out[38][13][11] + xor_out[39][13][11];
assign sum_out[8][13][11] = xor_out[40][13][11] + xor_out[41][13][11] + xor_out[42][13][11] + xor_out[43][13][11] + xor_out[44][13][11];
assign sum_out[9][13][11] = xor_out[45][13][11] + xor_out[46][13][11] + xor_out[47][13][11] + xor_out[48][13][11] + xor_out[49][13][11];
assign sum_out[10][13][11] = xor_out[50][13][11] + xor_out[51][13][11] + xor_out[52][13][11] + xor_out[53][13][11] + xor_out[54][13][11];
assign sum_out[11][13][11] = xor_out[55][13][11] + xor_out[56][13][11] + xor_out[57][13][11] + xor_out[58][13][11] + xor_out[59][13][11];
assign sum_out[12][13][11] = xor_out[60][13][11] + xor_out[61][13][11] + xor_out[62][13][11] + xor_out[63][13][11] + xor_out[64][13][11];
assign sum_out[13][13][11] = xor_out[65][13][11] + xor_out[66][13][11] + xor_out[67][13][11] + xor_out[68][13][11] + xor_out[69][13][11];
assign sum_out[14][13][11] = xor_out[70][13][11] + xor_out[71][13][11] + xor_out[72][13][11] + xor_out[73][13][11] + xor_out[74][13][11];
assign sum_out[15][13][11] = xor_out[75][13][11] + xor_out[76][13][11] + xor_out[77][13][11] + xor_out[78][13][11] + xor_out[79][13][11];
assign sum_out[16][13][11] = xor_out[80][13][11] + xor_out[81][13][11] + xor_out[82][13][11] + xor_out[83][13][11] + xor_out[84][13][11];
assign sum_out[17][13][11] = xor_out[85][13][11] + xor_out[86][13][11] + xor_out[87][13][11] + xor_out[88][13][11] + xor_out[89][13][11];
assign sum_out[18][13][11] = xor_out[90][13][11] + xor_out[91][13][11] + xor_out[92][13][11] + xor_out[93][13][11] + xor_out[94][13][11];
assign sum_out[19][13][11] = xor_out[95][13][11] + xor_out[96][13][11] + xor_out[97][13][11] + xor_out[98][13][11] + xor_out[99][13][11];

assign sum_out[0][13][12] = xor_out[0][13][12] + xor_out[1][13][12] + xor_out[2][13][12] + xor_out[3][13][12] + xor_out[4][13][12];
assign sum_out[1][13][12] = xor_out[5][13][12] + xor_out[6][13][12] + xor_out[7][13][12] + xor_out[8][13][12] + xor_out[9][13][12];
assign sum_out[2][13][12] = xor_out[10][13][12] + xor_out[11][13][12] + xor_out[12][13][12] + xor_out[13][13][12] + xor_out[14][13][12];
assign sum_out[3][13][12] = xor_out[15][13][12] + xor_out[16][13][12] + xor_out[17][13][12] + xor_out[18][13][12] + xor_out[19][13][12];
assign sum_out[4][13][12] = xor_out[20][13][12] + xor_out[21][13][12] + xor_out[22][13][12] + xor_out[23][13][12] + xor_out[24][13][12];
assign sum_out[5][13][12] = xor_out[25][13][12] + xor_out[26][13][12] + xor_out[27][13][12] + xor_out[28][13][12] + xor_out[29][13][12];
assign sum_out[6][13][12] = xor_out[30][13][12] + xor_out[31][13][12] + xor_out[32][13][12] + xor_out[33][13][12] + xor_out[34][13][12];
assign sum_out[7][13][12] = xor_out[35][13][12] + xor_out[36][13][12] + xor_out[37][13][12] + xor_out[38][13][12] + xor_out[39][13][12];
assign sum_out[8][13][12] = xor_out[40][13][12] + xor_out[41][13][12] + xor_out[42][13][12] + xor_out[43][13][12] + xor_out[44][13][12];
assign sum_out[9][13][12] = xor_out[45][13][12] + xor_out[46][13][12] + xor_out[47][13][12] + xor_out[48][13][12] + xor_out[49][13][12];
assign sum_out[10][13][12] = xor_out[50][13][12] + xor_out[51][13][12] + xor_out[52][13][12] + xor_out[53][13][12] + xor_out[54][13][12];
assign sum_out[11][13][12] = xor_out[55][13][12] + xor_out[56][13][12] + xor_out[57][13][12] + xor_out[58][13][12] + xor_out[59][13][12];
assign sum_out[12][13][12] = xor_out[60][13][12] + xor_out[61][13][12] + xor_out[62][13][12] + xor_out[63][13][12] + xor_out[64][13][12];
assign sum_out[13][13][12] = xor_out[65][13][12] + xor_out[66][13][12] + xor_out[67][13][12] + xor_out[68][13][12] + xor_out[69][13][12];
assign sum_out[14][13][12] = xor_out[70][13][12] + xor_out[71][13][12] + xor_out[72][13][12] + xor_out[73][13][12] + xor_out[74][13][12];
assign sum_out[15][13][12] = xor_out[75][13][12] + xor_out[76][13][12] + xor_out[77][13][12] + xor_out[78][13][12] + xor_out[79][13][12];
assign sum_out[16][13][12] = xor_out[80][13][12] + xor_out[81][13][12] + xor_out[82][13][12] + xor_out[83][13][12] + xor_out[84][13][12];
assign sum_out[17][13][12] = xor_out[85][13][12] + xor_out[86][13][12] + xor_out[87][13][12] + xor_out[88][13][12] + xor_out[89][13][12];
assign sum_out[18][13][12] = xor_out[90][13][12] + xor_out[91][13][12] + xor_out[92][13][12] + xor_out[93][13][12] + xor_out[94][13][12];
assign sum_out[19][13][12] = xor_out[95][13][12] + xor_out[96][13][12] + xor_out[97][13][12] + xor_out[98][13][12] + xor_out[99][13][12];

assign sum_out[0][13][13] = xor_out[0][13][13] + xor_out[1][13][13] + xor_out[2][13][13] + xor_out[3][13][13] + xor_out[4][13][13];
assign sum_out[1][13][13] = xor_out[5][13][13] + xor_out[6][13][13] + xor_out[7][13][13] + xor_out[8][13][13] + xor_out[9][13][13];
assign sum_out[2][13][13] = xor_out[10][13][13] + xor_out[11][13][13] + xor_out[12][13][13] + xor_out[13][13][13] + xor_out[14][13][13];
assign sum_out[3][13][13] = xor_out[15][13][13] + xor_out[16][13][13] + xor_out[17][13][13] + xor_out[18][13][13] + xor_out[19][13][13];
assign sum_out[4][13][13] = xor_out[20][13][13] + xor_out[21][13][13] + xor_out[22][13][13] + xor_out[23][13][13] + xor_out[24][13][13];
assign sum_out[5][13][13] = xor_out[25][13][13] + xor_out[26][13][13] + xor_out[27][13][13] + xor_out[28][13][13] + xor_out[29][13][13];
assign sum_out[6][13][13] = xor_out[30][13][13] + xor_out[31][13][13] + xor_out[32][13][13] + xor_out[33][13][13] + xor_out[34][13][13];
assign sum_out[7][13][13] = xor_out[35][13][13] + xor_out[36][13][13] + xor_out[37][13][13] + xor_out[38][13][13] + xor_out[39][13][13];
assign sum_out[8][13][13] = xor_out[40][13][13] + xor_out[41][13][13] + xor_out[42][13][13] + xor_out[43][13][13] + xor_out[44][13][13];
assign sum_out[9][13][13] = xor_out[45][13][13] + xor_out[46][13][13] + xor_out[47][13][13] + xor_out[48][13][13] + xor_out[49][13][13];
assign sum_out[10][13][13] = xor_out[50][13][13] + xor_out[51][13][13] + xor_out[52][13][13] + xor_out[53][13][13] + xor_out[54][13][13];
assign sum_out[11][13][13] = xor_out[55][13][13] + xor_out[56][13][13] + xor_out[57][13][13] + xor_out[58][13][13] + xor_out[59][13][13];
assign sum_out[12][13][13] = xor_out[60][13][13] + xor_out[61][13][13] + xor_out[62][13][13] + xor_out[63][13][13] + xor_out[64][13][13];
assign sum_out[13][13][13] = xor_out[65][13][13] + xor_out[66][13][13] + xor_out[67][13][13] + xor_out[68][13][13] + xor_out[69][13][13];
assign sum_out[14][13][13] = xor_out[70][13][13] + xor_out[71][13][13] + xor_out[72][13][13] + xor_out[73][13][13] + xor_out[74][13][13];
assign sum_out[15][13][13] = xor_out[75][13][13] + xor_out[76][13][13] + xor_out[77][13][13] + xor_out[78][13][13] + xor_out[79][13][13];
assign sum_out[16][13][13] = xor_out[80][13][13] + xor_out[81][13][13] + xor_out[82][13][13] + xor_out[83][13][13] + xor_out[84][13][13];
assign sum_out[17][13][13] = xor_out[85][13][13] + xor_out[86][13][13] + xor_out[87][13][13] + xor_out[88][13][13] + xor_out[89][13][13];
assign sum_out[18][13][13] = xor_out[90][13][13] + xor_out[91][13][13] + xor_out[92][13][13] + xor_out[93][13][13] + xor_out[94][13][13];
assign sum_out[19][13][13] = xor_out[95][13][13] + xor_out[96][13][13] + xor_out[97][13][13] + xor_out[98][13][13] + xor_out[99][13][13];

assign sum_out[0][13][14] = xor_out[0][13][14] + xor_out[1][13][14] + xor_out[2][13][14] + xor_out[3][13][14] + xor_out[4][13][14];
assign sum_out[1][13][14] = xor_out[5][13][14] + xor_out[6][13][14] + xor_out[7][13][14] + xor_out[8][13][14] + xor_out[9][13][14];
assign sum_out[2][13][14] = xor_out[10][13][14] + xor_out[11][13][14] + xor_out[12][13][14] + xor_out[13][13][14] + xor_out[14][13][14];
assign sum_out[3][13][14] = xor_out[15][13][14] + xor_out[16][13][14] + xor_out[17][13][14] + xor_out[18][13][14] + xor_out[19][13][14];
assign sum_out[4][13][14] = xor_out[20][13][14] + xor_out[21][13][14] + xor_out[22][13][14] + xor_out[23][13][14] + xor_out[24][13][14];
assign sum_out[5][13][14] = xor_out[25][13][14] + xor_out[26][13][14] + xor_out[27][13][14] + xor_out[28][13][14] + xor_out[29][13][14];
assign sum_out[6][13][14] = xor_out[30][13][14] + xor_out[31][13][14] + xor_out[32][13][14] + xor_out[33][13][14] + xor_out[34][13][14];
assign sum_out[7][13][14] = xor_out[35][13][14] + xor_out[36][13][14] + xor_out[37][13][14] + xor_out[38][13][14] + xor_out[39][13][14];
assign sum_out[8][13][14] = xor_out[40][13][14] + xor_out[41][13][14] + xor_out[42][13][14] + xor_out[43][13][14] + xor_out[44][13][14];
assign sum_out[9][13][14] = xor_out[45][13][14] + xor_out[46][13][14] + xor_out[47][13][14] + xor_out[48][13][14] + xor_out[49][13][14];
assign sum_out[10][13][14] = xor_out[50][13][14] + xor_out[51][13][14] + xor_out[52][13][14] + xor_out[53][13][14] + xor_out[54][13][14];
assign sum_out[11][13][14] = xor_out[55][13][14] + xor_out[56][13][14] + xor_out[57][13][14] + xor_out[58][13][14] + xor_out[59][13][14];
assign sum_out[12][13][14] = xor_out[60][13][14] + xor_out[61][13][14] + xor_out[62][13][14] + xor_out[63][13][14] + xor_out[64][13][14];
assign sum_out[13][13][14] = xor_out[65][13][14] + xor_out[66][13][14] + xor_out[67][13][14] + xor_out[68][13][14] + xor_out[69][13][14];
assign sum_out[14][13][14] = xor_out[70][13][14] + xor_out[71][13][14] + xor_out[72][13][14] + xor_out[73][13][14] + xor_out[74][13][14];
assign sum_out[15][13][14] = xor_out[75][13][14] + xor_out[76][13][14] + xor_out[77][13][14] + xor_out[78][13][14] + xor_out[79][13][14];
assign sum_out[16][13][14] = xor_out[80][13][14] + xor_out[81][13][14] + xor_out[82][13][14] + xor_out[83][13][14] + xor_out[84][13][14];
assign sum_out[17][13][14] = xor_out[85][13][14] + xor_out[86][13][14] + xor_out[87][13][14] + xor_out[88][13][14] + xor_out[89][13][14];
assign sum_out[18][13][14] = xor_out[90][13][14] + xor_out[91][13][14] + xor_out[92][13][14] + xor_out[93][13][14] + xor_out[94][13][14];
assign sum_out[19][13][14] = xor_out[95][13][14] + xor_out[96][13][14] + xor_out[97][13][14] + xor_out[98][13][14] + xor_out[99][13][14];

assign sum_out[0][13][15] = xor_out[0][13][15] + xor_out[1][13][15] + xor_out[2][13][15] + xor_out[3][13][15] + xor_out[4][13][15];
assign sum_out[1][13][15] = xor_out[5][13][15] + xor_out[6][13][15] + xor_out[7][13][15] + xor_out[8][13][15] + xor_out[9][13][15];
assign sum_out[2][13][15] = xor_out[10][13][15] + xor_out[11][13][15] + xor_out[12][13][15] + xor_out[13][13][15] + xor_out[14][13][15];
assign sum_out[3][13][15] = xor_out[15][13][15] + xor_out[16][13][15] + xor_out[17][13][15] + xor_out[18][13][15] + xor_out[19][13][15];
assign sum_out[4][13][15] = xor_out[20][13][15] + xor_out[21][13][15] + xor_out[22][13][15] + xor_out[23][13][15] + xor_out[24][13][15];
assign sum_out[5][13][15] = xor_out[25][13][15] + xor_out[26][13][15] + xor_out[27][13][15] + xor_out[28][13][15] + xor_out[29][13][15];
assign sum_out[6][13][15] = xor_out[30][13][15] + xor_out[31][13][15] + xor_out[32][13][15] + xor_out[33][13][15] + xor_out[34][13][15];
assign sum_out[7][13][15] = xor_out[35][13][15] + xor_out[36][13][15] + xor_out[37][13][15] + xor_out[38][13][15] + xor_out[39][13][15];
assign sum_out[8][13][15] = xor_out[40][13][15] + xor_out[41][13][15] + xor_out[42][13][15] + xor_out[43][13][15] + xor_out[44][13][15];
assign sum_out[9][13][15] = xor_out[45][13][15] + xor_out[46][13][15] + xor_out[47][13][15] + xor_out[48][13][15] + xor_out[49][13][15];
assign sum_out[10][13][15] = xor_out[50][13][15] + xor_out[51][13][15] + xor_out[52][13][15] + xor_out[53][13][15] + xor_out[54][13][15];
assign sum_out[11][13][15] = xor_out[55][13][15] + xor_out[56][13][15] + xor_out[57][13][15] + xor_out[58][13][15] + xor_out[59][13][15];
assign sum_out[12][13][15] = xor_out[60][13][15] + xor_out[61][13][15] + xor_out[62][13][15] + xor_out[63][13][15] + xor_out[64][13][15];
assign sum_out[13][13][15] = xor_out[65][13][15] + xor_out[66][13][15] + xor_out[67][13][15] + xor_out[68][13][15] + xor_out[69][13][15];
assign sum_out[14][13][15] = xor_out[70][13][15] + xor_out[71][13][15] + xor_out[72][13][15] + xor_out[73][13][15] + xor_out[74][13][15];
assign sum_out[15][13][15] = xor_out[75][13][15] + xor_out[76][13][15] + xor_out[77][13][15] + xor_out[78][13][15] + xor_out[79][13][15];
assign sum_out[16][13][15] = xor_out[80][13][15] + xor_out[81][13][15] + xor_out[82][13][15] + xor_out[83][13][15] + xor_out[84][13][15];
assign sum_out[17][13][15] = xor_out[85][13][15] + xor_out[86][13][15] + xor_out[87][13][15] + xor_out[88][13][15] + xor_out[89][13][15];
assign sum_out[18][13][15] = xor_out[90][13][15] + xor_out[91][13][15] + xor_out[92][13][15] + xor_out[93][13][15] + xor_out[94][13][15];
assign sum_out[19][13][15] = xor_out[95][13][15] + xor_out[96][13][15] + xor_out[97][13][15] + xor_out[98][13][15] + xor_out[99][13][15];

assign sum_out[0][13][16] = xor_out[0][13][16] + xor_out[1][13][16] + xor_out[2][13][16] + xor_out[3][13][16] + xor_out[4][13][16];
assign sum_out[1][13][16] = xor_out[5][13][16] + xor_out[6][13][16] + xor_out[7][13][16] + xor_out[8][13][16] + xor_out[9][13][16];
assign sum_out[2][13][16] = xor_out[10][13][16] + xor_out[11][13][16] + xor_out[12][13][16] + xor_out[13][13][16] + xor_out[14][13][16];
assign sum_out[3][13][16] = xor_out[15][13][16] + xor_out[16][13][16] + xor_out[17][13][16] + xor_out[18][13][16] + xor_out[19][13][16];
assign sum_out[4][13][16] = xor_out[20][13][16] + xor_out[21][13][16] + xor_out[22][13][16] + xor_out[23][13][16] + xor_out[24][13][16];
assign sum_out[5][13][16] = xor_out[25][13][16] + xor_out[26][13][16] + xor_out[27][13][16] + xor_out[28][13][16] + xor_out[29][13][16];
assign sum_out[6][13][16] = xor_out[30][13][16] + xor_out[31][13][16] + xor_out[32][13][16] + xor_out[33][13][16] + xor_out[34][13][16];
assign sum_out[7][13][16] = xor_out[35][13][16] + xor_out[36][13][16] + xor_out[37][13][16] + xor_out[38][13][16] + xor_out[39][13][16];
assign sum_out[8][13][16] = xor_out[40][13][16] + xor_out[41][13][16] + xor_out[42][13][16] + xor_out[43][13][16] + xor_out[44][13][16];
assign sum_out[9][13][16] = xor_out[45][13][16] + xor_out[46][13][16] + xor_out[47][13][16] + xor_out[48][13][16] + xor_out[49][13][16];
assign sum_out[10][13][16] = xor_out[50][13][16] + xor_out[51][13][16] + xor_out[52][13][16] + xor_out[53][13][16] + xor_out[54][13][16];
assign sum_out[11][13][16] = xor_out[55][13][16] + xor_out[56][13][16] + xor_out[57][13][16] + xor_out[58][13][16] + xor_out[59][13][16];
assign sum_out[12][13][16] = xor_out[60][13][16] + xor_out[61][13][16] + xor_out[62][13][16] + xor_out[63][13][16] + xor_out[64][13][16];
assign sum_out[13][13][16] = xor_out[65][13][16] + xor_out[66][13][16] + xor_out[67][13][16] + xor_out[68][13][16] + xor_out[69][13][16];
assign sum_out[14][13][16] = xor_out[70][13][16] + xor_out[71][13][16] + xor_out[72][13][16] + xor_out[73][13][16] + xor_out[74][13][16];
assign sum_out[15][13][16] = xor_out[75][13][16] + xor_out[76][13][16] + xor_out[77][13][16] + xor_out[78][13][16] + xor_out[79][13][16];
assign sum_out[16][13][16] = xor_out[80][13][16] + xor_out[81][13][16] + xor_out[82][13][16] + xor_out[83][13][16] + xor_out[84][13][16];
assign sum_out[17][13][16] = xor_out[85][13][16] + xor_out[86][13][16] + xor_out[87][13][16] + xor_out[88][13][16] + xor_out[89][13][16];
assign sum_out[18][13][16] = xor_out[90][13][16] + xor_out[91][13][16] + xor_out[92][13][16] + xor_out[93][13][16] + xor_out[94][13][16];
assign sum_out[19][13][16] = xor_out[95][13][16] + xor_out[96][13][16] + xor_out[97][13][16] + xor_out[98][13][16] + xor_out[99][13][16];

assign sum_out[0][13][17] = xor_out[0][13][17] + xor_out[1][13][17] + xor_out[2][13][17] + xor_out[3][13][17] + xor_out[4][13][17];
assign sum_out[1][13][17] = xor_out[5][13][17] + xor_out[6][13][17] + xor_out[7][13][17] + xor_out[8][13][17] + xor_out[9][13][17];
assign sum_out[2][13][17] = xor_out[10][13][17] + xor_out[11][13][17] + xor_out[12][13][17] + xor_out[13][13][17] + xor_out[14][13][17];
assign sum_out[3][13][17] = xor_out[15][13][17] + xor_out[16][13][17] + xor_out[17][13][17] + xor_out[18][13][17] + xor_out[19][13][17];
assign sum_out[4][13][17] = xor_out[20][13][17] + xor_out[21][13][17] + xor_out[22][13][17] + xor_out[23][13][17] + xor_out[24][13][17];
assign sum_out[5][13][17] = xor_out[25][13][17] + xor_out[26][13][17] + xor_out[27][13][17] + xor_out[28][13][17] + xor_out[29][13][17];
assign sum_out[6][13][17] = xor_out[30][13][17] + xor_out[31][13][17] + xor_out[32][13][17] + xor_out[33][13][17] + xor_out[34][13][17];
assign sum_out[7][13][17] = xor_out[35][13][17] + xor_out[36][13][17] + xor_out[37][13][17] + xor_out[38][13][17] + xor_out[39][13][17];
assign sum_out[8][13][17] = xor_out[40][13][17] + xor_out[41][13][17] + xor_out[42][13][17] + xor_out[43][13][17] + xor_out[44][13][17];
assign sum_out[9][13][17] = xor_out[45][13][17] + xor_out[46][13][17] + xor_out[47][13][17] + xor_out[48][13][17] + xor_out[49][13][17];
assign sum_out[10][13][17] = xor_out[50][13][17] + xor_out[51][13][17] + xor_out[52][13][17] + xor_out[53][13][17] + xor_out[54][13][17];
assign sum_out[11][13][17] = xor_out[55][13][17] + xor_out[56][13][17] + xor_out[57][13][17] + xor_out[58][13][17] + xor_out[59][13][17];
assign sum_out[12][13][17] = xor_out[60][13][17] + xor_out[61][13][17] + xor_out[62][13][17] + xor_out[63][13][17] + xor_out[64][13][17];
assign sum_out[13][13][17] = xor_out[65][13][17] + xor_out[66][13][17] + xor_out[67][13][17] + xor_out[68][13][17] + xor_out[69][13][17];
assign sum_out[14][13][17] = xor_out[70][13][17] + xor_out[71][13][17] + xor_out[72][13][17] + xor_out[73][13][17] + xor_out[74][13][17];
assign sum_out[15][13][17] = xor_out[75][13][17] + xor_out[76][13][17] + xor_out[77][13][17] + xor_out[78][13][17] + xor_out[79][13][17];
assign sum_out[16][13][17] = xor_out[80][13][17] + xor_out[81][13][17] + xor_out[82][13][17] + xor_out[83][13][17] + xor_out[84][13][17];
assign sum_out[17][13][17] = xor_out[85][13][17] + xor_out[86][13][17] + xor_out[87][13][17] + xor_out[88][13][17] + xor_out[89][13][17];
assign sum_out[18][13][17] = xor_out[90][13][17] + xor_out[91][13][17] + xor_out[92][13][17] + xor_out[93][13][17] + xor_out[94][13][17];
assign sum_out[19][13][17] = xor_out[95][13][17] + xor_out[96][13][17] + xor_out[97][13][17] + xor_out[98][13][17] + xor_out[99][13][17];

assign sum_out[0][13][18] = xor_out[0][13][18] + xor_out[1][13][18] + xor_out[2][13][18] + xor_out[3][13][18] + xor_out[4][13][18];
assign sum_out[1][13][18] = xor_out[5][13][18] + xor_out[6][13][18] + xor_out[7][13][18] + xor_out[8][13][18] + xor_out[9][13][18];
assign sum_out[2][13][18] = xor_out[10][13][18] + xor_out[11][13][18] + xor_out[12][13][18] + xor_out[13][13][18] + xor_out[14][13][18];
assign sum_out[3][13][18] = xor_out[15][13][18] + xor_out[16][13][18] + xor_out[17][13][18] + xor_out[18][13][18] + xor_out[19][13][18];
assign sum_out[4][13][18] = xor_out[20][13][18] + xor_out[21][13][18] + xor_out[22][13][18] + xor_out[23][13][18] + xor_out[24][13][18];
assign sum_out[5][13][18] = xor_out[25][13][18] + xor_out[26][13][18] + xor_out[27][13][18] + xor_out[28][13][18] + xor_out[29][13][18];
assign sum_out[6][13][18] = xor_out[30][13][18] + xor_out[31][13][18] + xor_out[32][13][18] + xor_out[33][13][18] + xor_out[34][13][18];
assign sum_out[7][13][18] = xor_out[35][13][18] + xor_out[36][13][18] + xor_out[37][13][18] + xor_out[38][13][18] + xor_out[39][13][18];
assign sum_out[8][13][18] = xor_out[40][13][18] + xor_out[41][13][18] + xor_out[42][13][18] + xor_out[43][13][18] + xor_out[44][13][18];
assign sum_out[9][13][18] = xor_out[45][13][18] + xor_out[46][13][18] + xor_out[47][13][18] + xor_out[48][13][18] + xor_out[49][13][18];
assign sum_out[10][13][18] = xor_out[50][13][18] + xor_out[51][13][18] + xor_out[52][13][18] + xor_out[53][13][18] + xor_out[54][13][18];
assign sum_out[11][13][18] = xor_out[55][13][18] + xor_out[56][13][18] + xor_out[57][13][18] + xor_out[58][13][18] + xor_out[59][13][18];
assign sum_out[12][13][18] = xor_out[60][13][18] + xor_out[61][13][18] + xor_out[62][13][18] + xor_out[63][13][18] + xor_out[64][13][18];
assign sum_out[13][13][18] = xor_out[65][13][18] + xor_out[66][13][18] + xor_out[67][13][18] + xor_out[68][13][18] + xor_out[69][13][18];
assign sum_out[14][13][18] = xor_out[70][13][18] + xor_out[71][13][18] + xor_out[72][13][18] + xor_out[73][13][18] + xor_out[74][13][18];
assign sum_out[15][13][18] = xor_out[75][13][18] + xor_out[76][13][18] + xor_out[77][13][18] + xor_out[78][13][18] + xor_out[79][13][18];
assign sum_out[16][13][18] = xor_out[80][13][18] + xor_out[81][13][18] + xor_out[82][13][18] + xor_out[83][13][18] + xor_out[84][13][18];
assign sum_out[17][13][18] = xor_out[85][13][18] + xor_out[86][13][18] + xor_out[87][13][18] + xor_out[88][13][18] + xor_out[89][13][18];
assign sum_out[18][13][18] = xor_out[90][13][18] + xor_out[91][13][18] + xor_out[92][13][18] + xor_out[93][13][18] + xor_out[94][13][18];
assign sum_out[19][13][18] = xor_out[95][13][18] + xor_out[96][13][18] + xor_out[97][13][18] + xor_out[98][13][18] + xor_out[99][13][18];

assign sum_out[0][13][19] = xor_out[0][13][19] + xor_out[1][13][19] + xor_out[2][13][19] + xor_out[3][13][19] + xor_out[4][13][19];
assign sum_out[1][13][19] = xor_out[5][13][19] + xor_out[6][13][19] + xor_out[7][13][19] + xor_out[8][13][19] + xor_out[9][13][19];
assign sum_out[2][13][19] = xor_out[10][13][19] + xor_out[11][13][19] + xor_out[12][13][19] + xor_out[13][13][19] + xor_out[14][13][19];
assign sum_out[3][13][19] = xor_out[15][13][19] + xor_out[16][13][19] + xor_out[17][13][19] + xor_out[18][13][19] + xor_out[19][13][19];
assign sum_out[4][13][19] = xor_out[20][13][19] + xor_out[21][13][19] + xor_out[22][13][19] + xor_out[23][13][19] + xor_out[24][13][19];
assign sum_out[5][13][19] = xor_out[25][13][19] + xor_out[26][13][19] + xor_out[27][13][19] + xor_out[28][13][19] + xor_out[29][13][19];
assign sum_out[6][13][19] = xor_out[30][13][19] + xor_out[31][13][19] + xor_out[32][13][19] + xor_out[33][13][19] + xor_out[34][13][19];
assign sum_out[7][13][19] = xor_out[35][13][19] + xor_out[36][13][19] + xor_out[37][13][19] + xor_out[38][13][19] + xor_out[39][13][19];
assign sum_out[8][13][19] = xor_out[40][13][19] + xor_out[41][13][19] + xor_out[42][13][19] + xor_out[43][13][19] + xor_out[44][13][19];
assign sum_out[9][13][19] = xor_out[45][13][19] + xor_out[46][13][19] + xor_out[47][13][19] + xor_out[48][13][19] + xor_out[49][13][19];
assign sum_out[10][13][19] = xor_out[50][13][19] + xor_out[51][13][19] + xor_out[52][13][19] + xor_out[53][13][19] + xor_out[54][13][19];
assign sum_out[11][13][19] = xor_out[55][13][19] + xor_out[56][13][19] + xor_out[57][13][19] + xor_out[58][13][19] + xor_out[59][13][19];
assign sum_out[12][13][19] = xor_out[60][13][19] + xor_out[61][13][19] + xor_out[62][13][19] + xor_out[63][13][19] + xor_out[64][13][19];
assign sum_out[13][13][19] = xor_out[65][13][19] + xor_out[66][13][19] + xor_out[67][13][19] + xor_out[68][13][19] + xor_out[69][13][19];
assign sum_out[14][13][19] = xor_out[70][13][19] + xor_out[71][13][19] + xor_out[72][13][19] + xor_out[73][13][19] + xor_out[74][13][19];
assign sum_out[15][13][19] = xor_out[75][13][19] + xor_out[76][13][19] + xor_out[77][13][19] + xor_out[78][13][19] + xor_out[79][13][19];
assign sum_out[16][13][19] = xor_out[80][13][19] + xor_out[81][13][19] + xor_out[82][13][19] + xor_out[83][13][19] + xor_out[84][13][19];
assign sum_out[17][13][19] = xor_out[85][13][19] + xor_out[86][13][19] + xor_out[87][13][19] + xor_out[88][13][19] + xor_out[89][13][19];
assign sum_out[18][13][19] = xor_out[90][13][19] + xor_out[91][13][19] + xor_out[92][13][19] + xor_out[93][13][19] + xor_out[94][13][19];
assign sum_out[19][13][19] = xor_out[95][13][19] + xor_out[96][13][19] + xor_out[97][13][19] + xor_out[98][13][19] + xor_out[99][13][19];

assign sum_out[0][13][20] = xor_out[0][13][20] + xor_out[1][13][20] + xor_out[2][13][20] + xor_out[3][13][20] + xor_out[4][13][20];
assign sum_out[1][13][20] = xor_out[5][13][20] + xor_out[6][13][20] + xor_out[7][13][20] + xor_out[8][13][20] + xor_out[9][13][20];
assign sum_out[2][13][20] = xor_out[10][13][20] + xor_out[11][13][20] + xor_out[12][13][20] + xor_out[13][13][20] + xor_out[14][13][20];
assign sum_out[3][13][20] = xor_out[15][13][20] + xor_out[16][13][20] + xor_out[17][13][20] + xor_out[18][13][20] + xor_out[19][13][20];
assign sum_out[4][13][20] = xor_out[20][13][20] + xor_out[21][13][20] + xor_out[22][13][20] + xor_out[23][13][20] + xor_out[24][13][20];
assign sum_out[5][13][20] = xor_out[25][13][20] + xor_out[26][13][20] + xor_out[27][13][20] + xor_out[28][13][20] + xor_out[29][13][20];
assign sum_out[6][13][20] = xor_out[30][13][20] + xor_out[31][13][20] + xor_out[32][13][20] + xor_out[33][13][20] + xor_out[34][13][20];
assign sum_out[7][13][20] = xor_out[35][13][20] + xor_out[36][13][20] + xor_out[37][13][20] + xor_out[38][13][20] + xor_out[39][13][20];
assign sum_out[8][13][20] = xor_out[40][13][20] + xor_out[41][13][20] + xor_out[42][13][20] + xor_out[43][13][20] + xor_out[44][13][20];
assign sum_out[9][13][20] = xor_out[45][13][20] + xor_out[46][13][20] + xor_out[47][13][20] + xor_out[48][13][20] + xor_out[49][13][20];
assign sum_out[10][13][20] = xor_out[50][13][20] + xor_out[51][13][20] + xor_out[52][13][20] + xor_out[53][13][20] + xor_out[54][13][20];
assign sum_out[11][13][20] = xor_out[55][13][20] + xor_out[56][13][20] + xor_out[57][13][20] + xor_out[58][13][20] + xor_out[59][13][20];
assign sum_out[12][13][20] = xor_out[60][13][20] + xor_out[61][13][20] + xor_out[62][13][20] + xor_out[63][13][20] + xor_out[64][13][20];
assign sum_out[13][13][20] = xor_out[65][13][20] + xor_out[66][13][20] + xor_out[67][13][20] + xor_out[68][13][20] + xor_out[69][13][20];
assign sum_out[14][13][20] = xor_out[70][13][20] + xor_out[71][13][20] + xor_out[72][13][20] + xor_out[73][13][20] + xor_out[74][13][20];
assign sum_out[15][13][20] = xor_out[75][13][20] + xor_out[76][13][20] + xor_out[77][13][20] + xor_out[78][13][20] + xor_out[79][13][20];
assign sum_out[16][13][20] = xor_out[80][13][20] + xor_out[81][13][20] + xor_out[82][13][20] + xor_out[83][13][20] + xor_out[84][13][20];
assign sum_out[17][13][20] = xor_out[85][13][20] + xor_out[86][13][20] + xor_out[87][13][20] + xor_out[88][13][20] + xor_out[89][13][20];
assign sum_out[18][13][20] = xor_out[90][13][20] + xor_out[91][13][20] + xor_out[92][13][20] + xor_out[93][13][20] + xor_out[94][13][20];
assign sum_out[19][13][20] = xor_out[95][13][20] + xor_out[96][13][20] + xor_out[97][13][20] + xor_out[98][13][20] + xor_out[99][13][20];

assign sum_out[0][13][21] = xor_out[0][13][21] + xor_out[1][13][21] + xor_out[2][13][21] + xor_out[3][13][21] + xor_out[4][13][21];
assign sum_out[1][13][21] = xor_out[5][13][21] + xor_out[6][13][21] + xor_out[7][13][21] + xor_out[8][13][21] + xor_out[9][13][21];
assign sum_out[2][13][21] = xor_out[10][13][21] + xor_out[11][13][21] + xor_out[12][13][21] + xor_out[13][13][21] + xor_out[14][13][21];
assign sum_out[3][13][21] = xor_out[15][13][21] + xor_out[16][13][21] + xor_out[17][13][21] + xor_out[18][13][21] + xor_out[19][13][21];
assign sum_out[4][13][21] = xor_out[20][13][21] + xor_out[21][13][21] + xor_out[22][13][21] + xor_out[23][13][21] + xor_out[24][13][21];
assign sum_out[5][13][21] = xor_out[25][13][21] + xor_out[26][13][21] + xor_out[27][13][21] + xor_out[28][13][21] + xor_out[29][13][21];
assign sum_out[6][13][21] = xor_out[30][13][21] + xor_out[31][13][21] + xor_out[32][13][21] + xor_out[33][13][21] + xor_out[34][13][21];
assign sum_out[7][13][21] = xor_out[35][13][21] + xor_out[36][13][21] + xor_out[37][13][21] + xor_out[38][13][21] + xor_out[39][13][21];
assign sum_out[8][13][21] = xor_out[40][13][21] + xor_out[41][13][21] + xor_out[42][13][21] + xor_out[43][13][21] + xor_out[44][13][21];
assign sum_out[9][13][21] = xor_out[45][13][21] + xor_out[46][13][21] + xor_out[47][13][21] + xor_out[48][13][21] + xor_out[49][13][21];
assign sum_out[10][13][21] = xor_out[50][13][21] + xor_out[51][13][21] + xor_out[52][13][21] + xor_out[53][13][21] + xor_out[54][13][21];
assign sum_out[11][13][21] = xor_out[55][13][21] + xor_out[56][13][21] + xor_out[57][13][21] + xor_out[58][13][21] + xor_out[59][13][21];
assign sum_out[12][13][21] = xor_out[60][13][21] + xor_out[61][13][21] + xor_out[62][13][21] + xor_out[63][13][21] + xor_out[64][13][21];
assign sum_out[13][13][21] = xor_out[65][13][21] + xor_out[66][13][21] + xor_out[67][13][21] + xor_out[68][13][21] + xor_out[69][13][21];
assign sum_out[14][13][21] = xor_out[70][13][21] + xor_out[71][13][21] + xor_out[72][13][21] + xor_out[73][13][21] + xor_out[74][13][21];
assign sum_out[15][13][21] = xor_out[75][13][21] + xor_out[76][13][21] + xor_out[77][13][21] + xor_out[78][13][21] + xor_out[79][13][21];
assign sum_out[16][13][21] = xor_out[80][13][21] + xor_out[81][13][21] + xor_out[82][13][21] + xor_out[83][13][21] + xor_out[84][13][21];
assign sum_out[17][13][21] = xor_out[85][13][21] + xor_out[86][13][21] + xor_out[87][13][21] + xor_out[88][13][21] + xor_out[89][13][21];
assign sum_out[18][13][21] = xor_out[90][13][21] + xor_out[91][13][21] + xor_out[92][13][21] + xor_out[93][13][21] + xor_out[94][13][21];
assign sum_out[19][13][21] = xor_out[95][13][21] + xor_out[96][13][21] + xor_out[97][13][21] + xor_out[98][13][21] + xor_out[99][13][21];

assign sum_out[0][13][22] = xor_out[0][13][22] + xor_out[1][13][22] + xor_out[2][13][22] + xor_out[3][13][22] + xor_out[4][13][22];
assign sum_out[1][13][22] = xor_out[5][13][22] + xor_out[6][13][22] + xor_out[7][13][22] + xor_out[8][13][22] + xor_out[9][13][22];
assign sum_out[2][13][22] = xor_out[10][13][22] + xor_out[11][13][22] + xor_out[12][13][22] + xor_out[13][13][22] + xor_out[14][13][22];
assign sum_out[3][13][22] = xor_out[15][13][22] + xor_out[16][13][22] + xor_out[17][13][22] + xor_out[18][13][22] + xor_out[19][13][22];
assign sum_out[4][13][22] = xor_out[20][13][22] + xor_out[21][13][22] + xor_out[22][13][22] + xor_out[23][13][22] + xor_out[24][13][22];
assign sum_out[5][13][22] = xor_out[25][13][22] + xor_out[26][13][22] + xor_out[27][13][22] + xor_out[28][13][22] + xor_out[29][13][22];
assign sum_out[6][13][22] = xor_out[30][13][22] + xor_out[31][13][22] + xor_out[32][13][22] + xor_out[33][13][22] + xor_out[34][13][22];
assign sum_out[7][13][22] = xor_out[35][13][22] + xor_out[36][13][22] + xor_out[37][13][22] + xor_out[38][13][22] + xor_out[39][13][22];
assign sum_out[8][13][22] = xor_out[40][13][22] + xor_out[41][13][22] + xor_out[42][13][22] + xor_out[43][13][22] + xor_out[44][13][22];
assign sum_out[9][13][22] = xor_out[45][13][22] + xor_out[46][13][22] + xor_out[47][13][22] + xor_out[48][13][22] + xor_out[49][13][22];
assign sum_out[10][13][22] = xor_out[50][13][22] + xor_out[51][13][22] + xor_out[52][13][22] + xor_out[53][13][22] + xor_out[54][13][22];
assign sum_out[11][13][22] = xor_out[55][13][22] + xor_out[56][13][22] + xor_out[57][13][22] + xor_out[58][13][22] + xor_out[59][13][22];
assign sum_out[12][13][22] = xor_out[60][13][22] + xor_out[61][13][22] + xor_out[62][13][22] + xor_out[63][13][22] + xor_out[64][13][22];
assign sum_out[13][13][22] = xor_out[65][13][22] + xor_out[66][13][22] + xor_out[67][13][22] + xor_out[68][13][22] + xor_out[69][13][22];
assign sum_out[14][13][22] = xor_out[70][13][22] + xor_out[71][13][22] + xor_out[72][13][22] + xor_out[73][13][22] + xor_out[74][13][22];
assign sum_out[15][13][22] = xor_out[75][13][22] + xor_out[76][13][22] + xor_out[77][13][22] + xor_out[78][13][22] + xor_out[79][13][22];
assign sum_out[16][13][22] = xor_out[80][13][22] + xor_out[81][13][22] + xor_out[82][13][22] + xor_out[83][13][22] + xor_out[84][13][22];
assign sum_out[17][13][22] = xor_out[85][13][22] + xor_out[86][13][22] + xor_out[87][13][22] + xor_out[88][13][22] + xor_out[89][13][22];
assign sum_out[18][13][22] = xor_out[90][13][22] + xor_out[91][13][22] + xor_out[92][13][22] + xor_out[93][13][22] + xor_out[94][13][22];
assign sum_out[19][13][22] = xor_out[95][13][22] + xor_out[96][13][22] + xor_out[97][13][22] + xor_out[98][13][22] + xor_out[99][13][22];

assign sum_out[0][13][23] = xor_out[0][13][23] + xor_out[1][13][23] + xor_out[2][13][23] + xor_out[3][13][23] + xor_out[4][13][23];
assign sum_out[1][13][23] = xor_out[5][13][23] + xor_out[6][13][23] + xor_out[7][13][23] + xor_out[8][13][23] + xor_out[9][13][23];
assign sum_out[2][13][23] = xor_out[10][13][23] + xor_out[11][13][23] + xor_out[12][13][23] + xor_out[13][13][23] + xor_out[14][13][23];
assign sum_out[3][13][23] = xor_out[15][13][23] + xor_out[16][13][23] + xor_out[17][13][23] + xor_out[18][13][23] + xor_out[19][13][23];
assign sum_out[4][13][23] = xor_out[20][13][23] + xor_out[21][13][23] + xor_out[22][13][23] + xor_out[23][13][23] + xor_out[24][13][23];
assign sum_out[5][13][23] = xor_out[25][13][23] + xor_out[26][13][23] + xor_out[27][13][23] + xor_out[28][13][23] + xor_out[29][13][23];
assign sum_out[6][13][23] = xor_out[30][13][23] + xor_out[31][13][23] + xor_out[32][13][23] + xor_out[33][13][23] + xor_out[34][13][23];
assign sum_out[7][13][23] = xor_out[35][13][23] + xor_out[36][13][23] + xor_out[37][13][23] + xor_out[38][13][23] + xor_out[39][13][23];
assign sum_out[8][13][23] = xor_out[40][13][23] + xor_out[41][13][23] + xor_out[42][13][23] + xor_out[43][13][23] + xor_out[44][13][23];
assign sum_out[9][13][23] = xor_out[45][13][23] + xor_out[46][13][23] + xor_out[47][13][23] + xor_out[48][13][23] + xor_out[49][13][23];
assign sum_out[10][13][23] = xor_out[50][13][23] + xor_out[51][13][23] + xor_out[52][13][23] + xor_out[53][13][23] + xor_out[54][13][23];
assign sum_out[11][13][23] = xor_out[55][13][23] + xor_out[56][13][23] + xor_out[57][13][23] + xor_out[58][13][23] + xor_out[59][13][23];
assign sum_out[12][13][23] = xor_out[60][13][23] + xor_out[61][13][23] + xor_out[62][13][23] + xor_out[63][13][23] + xor_out[64][13][23];
assign sum_out[13][13][23] = xor_out[65][13][23] + xor_out[66][13][23] + xor_out[67][13][23] + xor_out[68][13][23] + xor_out[69][13][23];
assign sum_out[14][13][23] = xor_out[70][13][23] + xor_out[71][13][23] + xor_out[72][13][23] + xor_out[73][13][23] + xor_out[74][13][23];
assign sum_out[15][13][23] = xor_out[75][13][23] + xor_out[76][13][23] + xor_out[77][13][23] + xor_out[78][13][23] + xor_out[79][13][23];
assign sum_out[16][13][23] = xor_out[80][13][23] + xor_out[81][13][23] + xor_out[82][13][23] + xor_out[83][13][23] + xor_out[84][13][23];
assign sum_out[17][13][23] = xor_out[85][13][23] + xor_out[86][13][23] + xor_out[87][13][23] + xor_out[88][13][23] + xor_out[89][13][23];
assign sum_out[18][13][23] = xor_out[90][13][23] + xor_out[91][13][23] + xor_out[92][13][23] + xor_out[93][13][23] + xor_out[94][13][23];
assign sum_out[19][13][23] = xor_out[95][13][23] + xor_out[96][13][23] + xor_out[97][13][23] + xor_out[98][13][23] + xor_out[99][13][23];

assign sum_out[0][14][0] = xor_out[0][14][0] + xor_out[1][14][0] + xor_out[2][14][0] + xor_out[3][14][0] + xor_out[4][14][0];
assign sum_out[1][14][0] = xor_out[5][14][0] + xor_out[6][14][0] + xor_out[7][14][0] + xor_out[8][14][0] + xor_out[9][14][0];
assign sum_out[2][14][0] = xor_out[10][14][0] + xor_out[11][14][0] + xor_out[12][14][0] + xor_out[13][14][0] + xor_out[14][14][0];
assign sum_out[3][14][0] = xor_out[15][14][0] + xor_out[16][14][0] + xor_out[17][14][0] + xor_out[18][14][0] + xor_out[19][14][0];
assign sum_out[4][14][0] = xor_out[20][14][0] + xor_out[21][14][0] + xor_out[22][14][0] + xor_out[23][14][0] + xor_out[24][14][0];
assign sum_out[5][14][0] = xor_out[25][14][0] + xor_out[26][14][0] + xor_out[27][14][0] + xor_out[28][14][0] + xor_out[29][14][0];
assign sum_out[6][14][0] = xor_out[30][14][0] + xor_out[31][14][0] + xor_out[32][14][0] + xor_out[33][14][0] + xor_out[34][14][0];
assign sum_out[7][14][0] = xor_out[35][14][0] + xor_out[36][14][0] + xor_out[37][14][0] + xor_out[38][14][0] + xor_out[39][14][0];
assign sum_out[8][14][0] = xor_out[40][14][0] + xor_out[41][14][0] + xor_out[42][14][0] + xor_out[43][14][0] + xor_out[44][14][0];
assign sum_out[9][14][0] = xor_out[45][14][0] + xor_out[46][14][0] + xor_out[47][14][0] + xor_out[48][14][0] + xor_out[49][14][0];
assign sum_out[10][14][0] = xor_out[50][14][0] + xor_out[51][14][0] + xor_out[52][14][0] + xor_out[53][14][0] + xor_out[54][14][0];
assign sum_out[11][14][0] = xor_out[55][14][0] + xor_out[56][14][0] + xor_out[57][14][0] + xor_out[58][14][0] + xor_out[59][14][0];
assign sum_out[12][14][0] = xor_out[60][14][0] + xor_out[61][14][0] + xor_out[62][14][0] + xor_out[63][14][0] + xor_out[64][14][0];
assign sum_out[13][14][0] = xor_out[65][14][0] + xor_out[66][14][0] + xor_out[67][14][0] + xor_out[68][14][0] + xor_out[69][14][0];
assign sum_out[14][14][0] = xor_out[70][14][0] + xor_out[71][14][0] + xor_out[72][14][0] + xor_out[73][14][0] + xor_out[74][14][0];
assign sum_out[15][14][0] = xor_out[75][14][0] + xor_out[76][14][0] + xor_out[77][14][0] + xor_out[78][14][0] + xor_out[79][14][0];
assign sum_out[16][14][0] = xor_out[80][14][0] + xor_out[81][14][0] + xor_out[82][14][0] + xor_out[83][14][0] + xor_out[84][14][0];
assign sum_out[17][14][0] = xor_out[85][14][0] + xor_out[86][14][0] + xor_out[87][14][0] + xor_out[88][14][0] + xor_out[89][14][0];
assign sum_out[18][14][0] = xor_out[90][14][0] + xor_out[91][14][0] + xor_out[92][14][0] + xor_out[93][14][0] + xor_out[94][14][0];
assign sum_out[19][14][0] = xor_out[95][14][0] + xor_out[96][14][0] + xor_out[97][14][0] + xor_out[98][14][0] + xor_out[99][14][0];

assign sum_out[0][14][1] = xor_out[0][14][1] + xor_out[1][14][1] + xor_out[2][14][1] + xor_out[3][14][1] + xor_out[4][14][1];
assign sum_out[1][14][1] = xor_out[5][14][1] + xor_out[6][14][1] + xor_out[7][14][1] + xor_out[8][14][1] + xor_out[9][14][1];
assign sum_out[2][14][1] = xor_out[10][14][1] + xor_out[11][14][1] + xor_out[12][14][1] + xor_out[13][14][1] + xor_out[14][14][1];
assign sum_out[3][14][1] = xor_out[15][14][1] + xor_out[16][14][1] + xor_out[17][14][1] + xor_out[18][14][1] + xor_out[19][14][1];
assign sum_out[4][14][1] = xor_out[20][14][1] + xor_out[21][14][1] + xor_out[22][14][1] + xor_out[23][14][1] + xor_out[24][14][1];
assign sum_out[5][14][1] = xor_out[25][14][1] + xor_out[26][14][1] + xor_out[27][14][1] + xor_out[28][14][1] + xor_out[29][14][1];
assign sum_out[6][14][1] = xor_out[30][14][1] + xor_out[31][14][1] + xor_out[32][14][1] + xor_out[33][14][1] + xor_out[34][14][1];
assign sum_out[7][14][1] = xor_out[35][14][1] + xor_out[36][14][1] + xor_out[37][14][1] + xor_out[38][14][1] + xor_out[39][14][1];
assign sum_out[8][14][1] = xor_out[40][14][1] + xor_out[41][14][1] + xor_out[42][14][1] + xor_out[43][14][1] + xor_out[44][14][1];
assign sum_out[9][14][1] = xor_out[45][14][1] + xor_out[46][14][1] + xor_out[47][14][1] + xor_out[48][14][1] + xor_out[49][14][1];
assign sum_out[10][14][1] = xor_out[50][14][1] + xor_out[51][14][1] + xor_out[52][14][1] + xor_out[53][14][1] + xor_out[54][14][1];
assign sum_out[11][14][1] = xor_out[55][14][1] + xor_out[56][14][1] + xor_out[57][14][1] + xor_out[58][14][1] + xor_out[59][14][1];
assign sum_out[12][14][1] = xor_out[60][14][1] + xor_out[61][14][1] + xor_out[62][14][1] + xor_out[63][14][1] + xor_out[64][14][1];
assign sum_out[13][14][1] = xor_out[65][14][1] + xor_out[66][14][1] + xor_out[67][14][1] + xor_out[68][14][1] + xor_out[69][14][1];
assign sum_out[14][14][1] = xor_out[70][14][1] + xor_out[71][14][1] + xor_out[72][14][1] + xor_out[73][14][1] + xor_out[74][14][1];
assign sum_out[15][14][1] = xor_out[75][14][1] + xor_out[76][14][1] + xor_out[77][14][1] + xor_out[78][14][1] + xor_out[79][14][1];
assign sum_out[16][14][1] = xor_out[80][14][1] + xor_out[81][14][1] + xor_out[82][14][1] + xor_out[83][14][1] + xor_out[84][14][1];
assign sum_out[17][14][1] = xor_out[85][14][1] + xor_out[86][14][1] + xor_out[87][14][1] + xor_out[88][14][1] + xor_out[89][14][1];
assign sum_out[18][14][1] = xor_out[90][14][1] + xor_out[91][14][1] + xor_out[92][14][1] + xor_out[93][14][1] + xor_out[94][14][1];
assign sum_out[19][14][1] = xor_out[95][14][1] + xor_out[96][14][1] + xor_out[97][14][1] + xor_out[98][14][1] + xor_out[99][14][1];

assign sum_out[0][14][2] = xor_out[0][14][2] + xor_out[1][14][2] + xor_out[2][14][2] + xor_out[3][14][2] + xor_out[4][14][2];
assign sum_out[1][14][2] = xor_out[5][14][2] + xor_out[6][14][2] + xor_out[7][14][2] + xor_out[8][14][2] + xor_out[9][14][2];
assign sum_out[2][14][2] = xor_out[10][14][2] + xor_out[11][14][2] + xor_out[12][14][2] + xor_out[13][14][2] + xor_out[14][14][2];
assign sum_out[3][14][2] = xor_out[15][14][2] + xor_out[16][14][2] + xor_out[17][14][2] + xor_out[18][14][2] + xor_out[19][14][2];
assign sum_out[4][14][2] = xor_out[20][14][2] + xor_out[21][14][2] + xor_out[22][14][2] + xor_out[23][14][2] + xor_out[24][14][2];
assign sum_out[5][14][2] = xor_out[25][14][2] + xor_out[26][14][2] + xor_out[27][14][2] + xor_out[28][14][2] + xor_out[29][14][2];
assign sum_out[6][14][2] = xor_out[30][14][2] + xor_out[31][14][2] + xor_out[32][14][2] + xor_out[33][14][2] + xor_out[34][14][2];
assign sum_out[7][14][2] = xor_out[35][14][2] + xor_out[36][14][2] + xor_out[37][14][2] + xor_out[38][14][2] + xor_out[39][14][2];
assign sum_out[8][14][2] = xor_out[40][14][2] + xor_out[41][14][2] + xor_out[42][14][2] + xor_out[43][14][2] + xor_out[44][14][2];
assign sum_out[9][14][2] = xor_out[45][14][2] + xor_out[46][14][2] + xor_out[47][14][2] + xor_out[48][14][2] + xor_out[49][14][2];
assign sum_out[10][14][2] = xor_out[50][14][2] + xor_out[51][14][2] + xor_out[52][14][2] + xor_out[53][14][2] + xor_out[54][14][2];
assign sum_out[11][14][2] = xor_out[55][14][2] + xor_out[56][14][2] + xor_out[57][14][2] + xor_out[58][14][2] + xor_out[59][14][2];
assign sum_out[12][14][2] = xor_out[60][14][2] + xor_out[61][14][2] + xor_out[62][14][2] + xor_out[63][14][2] + xor_out[64][14][2];
assign sum_out[13][14][2] = xor_out[65][14][2] + xor_out[66][14][2] + xor_out[67][14][2] + xor_out[68][14][2] + xor_out[69][14][2];
assign sum_out[14][14][2] = xor_out[70][14][2] + xor_out[71][14][2] + xor_out[72][14][2] + xor_out[73][14][2] + xor_out[74][14][2];
assign sum_out[15][14][2] = xor_out[75][14][2] + xor_out[76][14][2] + xor_out[77][14][2] + xor_out[78][14][2] + xor_out[79][14][2];
assign sum_out[16][14][2] = xor_out[80][14][2] + xor_out[81][14][2] + xor_out[82][14][2] + xor_out[83][14][2] + xor_out[84][14][2];
assign sum_out[17][14][2] = xor_out[85][14][2] + xor_out[86][14][2] + xor_out[87][14][2] + xor_out[88][14][2] + xor_out[89][14][2];
assign sum_out[18][14][2] = xor_out[90][14][2] + xor_out[91][14][2] + xor_out[92][14][2] + xor_out[93][14][2] + xor_out[94][14][2];
assign sum_out[19][14][2] = xor_out[95][14][2] + xor_out[96][14][2] + xor_out[97][14][2] + xor_out[98][14][2] + xor_out[99][14][2];

assign sum_out[0][14][3] = xor_out[0][14][3] + xor_out[1][14][3] + xor_out[2][14][3] + xor_out[3][14][3] + xor_out[4][14][3];
assign sum_out[1][14][3] = xor_out[5][14][3] + xor_out[6][14][3] + xor_out[7][14][3] + xor_out[8][14][3] + xor_out[9][14][3];
assign sum_out[2][14][3] = xor_out[10][14][3] + xor_out[11][14][3] + xor_out[12][14][3] + xor_out[13][14][3] + xor_out[14][14][3];
assign sum_out[3][14][3] = xor_out[15][14][3] + xor_out[16][14][3] + xor_out[17][14][3] + xor_out[18][14][3] + xor_out[19][14][3];
assign sum_out[4][14][3] = xor_out[20][14][3] + xor_out[21][14][3] + xor_out[22][14][3] + xor_out[23][14][3] + xor_out[24][14][3];
assign sum_out[5][14][3] = xor_out[25][14][3] + xor_out[26][14][3] + xor_out[27][14][3] + xor_out[28][14][3] + xor_out[29][14][3];
assign sum_out[6][14][3] = xor_out[30][14][3] + xor_out[31][14][3] + xor_out[32][14][3] + xor_out[33][14][3] + xor_out[34][14][3];
assign sum_out[7][14][3] = xor_out[35][14][3] + xor_out[36][14][3] + xor_out[37][14][3] + xor_out[38][14][3] + xor_out[39][14][3];
assign sum_out[8][14][3] = xor_out[40][14][3] + xor_out[41][14][3] + xor_out[42][14][3] + xor_out[43][14][3] + xor_out[44][14][3];
assign sum_out[9][14][3] = xor_out[45][14][3] + xor_out[46][14][3] + xor_out[47][14][3] + xor_out[48][14][3] + xor_out[49][14][3];
assign sum_out[10][14][3] = xor_out[50][14][3] + xor_out[51][14][3] + xor_out[52][14][3] + xor_out[53][14][3] + xor_out[54][14][3];
assign sum_out[11][14][3] = xor_out[55][14][3] + xor_out[56][14][3] + xor_out[57][14][3] + xor_out[58][14][3] + xor_out[59][14][3];
assign sum_out[12][14][3] = xor_out[60][14][3] + xor_out[61][14][3] + xor_out[62][14][3] + xor_out[63][14][3] + xor_out[64][14][3];
assign sum_out[13][14][3] = xor_out[65][14][3] + xor_out[66][14][3] + xor_out[67][14][3] + xor_out[68][14][3] + xor_out[69][14][3];
assign sum_out[14][14][3] = xor_out[70][14][3] + xor_out[71][14][3] + xor_out[72][14][3] + xor_out[73][14][3] + xor_out[74][14][3];
assign sum_out[15][14][3] = xor_out[75][14][3] + xor_out[76][14][3] + xor_out[77][14][3] + xor_out[78][14][3] + xor_out[79][14][3];
assign sum_out[16][14][3] = xor_out[80][14][3] + xor_out[81][14][3] + xor_out[82][14][3] + xor_out[83][14][3] + xor_out[84][14][3];
assign sum_out[17][14][3] = xor_out[85][14][3] + xor_out[86][14][3] + xor_out[87][14][3] + xor_out[88][14][3] + xor_out[89][14][3];
assign sum_out[18][14][3] = xor_out[90][14][3] + xor_out[91][14][3] + xor_out[92][14][3] + xor_out[93][14][3] + xor_out[94][14][3];
assign sum_out[19][14][3] = xor_out[95][14][3] + xor_out[96][14][3] + xor_out[97][14][3] + xor_out[98][14][3] + xor_out[99][14][3];

assign sum_out[0][14][4] = xor_out[0][14][4] + xor_out[1][14][4] + xor_out[2][14][4] + xor_out[3][14][4] + xor_out[4][14][4];
assign sum_out[1][14][4] = xor_out[5][14][4] + xor_out[6][14][4] + xor_out[7][14][4] + xor_out[8][14][4] + xor_out[9][14][4];
assign sum_out[2][14][4] = xor_out[10][14][4] + xor_out[11][14][4] + xor_out[12][14][4] + xor_out[13][14][4] + xor_out[14][14][4];
assign sum_out[3][14][4] = xor_out[15][14][4] + xor_out[16][14][4] + xor_out[17][14][4] + xor_out[18][14][4] + xor_out[19][14][4];
assign sum_out[4][14][4] = xor_out[20][14][4] + xor_out[21][14][4] + xor_out[22][14][4] + xor_out[23][14][4] + xor_out[24][14][4];
assign sum_out[5][14][4] = xor_out[25][14][4] + xor_out[26][14][4] + xor_out[27][14][4] + xor_out[28][14][4] + xor_out[29][14][4];
assign sum_out[6][14][4] = xor_out[30][14][4] + xor_out[31][14][4] + xor_out[32][14][4] + xor_out[33][14][4] + xor_out[34][14][4];
assign sum_out[7][14][4] = xor_out[35][14][4] + xor_out[36][14][4] + xor_out[37][14][4] + xor_out[38][14][4] + xor_out[39][14][4];
assign sum_out[8][14][4] = xor_out[40][14][4] + xor_out[41][14][4] + xor_out[42][14][4] + xor_out[43][14][4] + xor_out[44][14][4];
assign sum_out[9][14][4] = xor_out[45][14][4] + xor_out[46][14][4] + xor_out[47][14][4] + xor_out[48][14][4] + xor_out[49][14][4];
assign sum_out[10][14][4] = xor_out[50][14][4] + xor_out[51][14][4] + xor_out[52][14][4] + xor_out[53][14][4] + xor_out[54][14][4];
assign sum_out[11][14][4] = xor_out[55][14][4] + xor_out[56][14][4] + xor_out[57][14][4] + xor_out[58][14][4] + xor_out[59][14][4];
assign sum_out[12][14][4] = xor_out[60][14][4] + xor_out[61][14][4] + xor_out[62][14][4] + xor_out[63][14][4] + xor_out[64][14][4];
assign sum_out[13][14][4] = xor_out[65][14][4] + xor_out[66][14][4] + xor_out[67][14][4] + xor_out[68][14][4] + xor_out[69][14][4];
assign sum_out[14][14][4] = xor_out[70][14][4] + xor_out[71][14][4] + xor_out[72][14][4] + xor_out[73][14][4] + xor_out[74][14][4];
assign sum_out[15][14][4] = xor_out[75][14][4] + xor_out[76][14][4] + xor_out[77][14][4] + xor_out[78][14][4] + xor_out[79][14][4];
assign sum_out[16][14][4] = xor_out[80][14][4] + xor_out[81][14][4] + xor_out[82][14][4] + xor_out[83][14][4] + xor_out[84][14][4];
assign sum_out[17][14][4] = xor_out[85][14][4] + xor_out[86][14][4] + xor_out[87][14][4] + xor_out[88][14][4] + xor_out[89][14][4];
assign sum_out[18][14][4] = xor_out[90][14][4] + xor_out[91][14][4] + xor_out[92][14][4] + xor_out[93][14][4] + xor_out[94][14][4];
assign sum_out[19][14][4] = xor_out[95][14][4] + xor_out[96][14][4] + xor_out[97][14][4] + xor_out[98][14][4] + xor_out[99][14][4];

assign sum_out[0][14][5] = xor_out[0][14][5] + xor_out[1][14][5] + xor_out[2][14][5] + xor_out[3][14][5] + xor_out[4][14][5];
assign sum_out[1][14][5] = xor_out[5][14][5] + xor_out[6][14][5] + xor_out[7][14][5] + xor_out[8][14][5] + xor_out[9][14][5];
assign sum_out[2][14][5] = xor_out[10][14][5] + xor_out[11][14][5] + xor_out[12][14][5] + xor_out[13][14][5] + xor_out[14][14][5];
assign sum_out[3][14][5] = xor_out[15][14][5] + xor_out[16][14][5] + xor_out[17][14][5] + xor_out[18][14][5] + xor_out[19][14][5];
assign sum_out[4][14][5] = xor_out[20][14][5] + xor_out[21][14][5] + xor_out[22][14][5] + xor_out[23][14][5] + xor_out[24][14][5];
assign sum_out[5][14][5] = xor_out[25][14][5] + xor_out[26][14][5] + xor_out[27][14][5] + xor_out[28][14][5] + xor_out[29][14][5];
assign sum_out[6][14][5] = xor_out[30][14][5] + xor_out[31][14][5] + xor_out[32][14][5] + xor_out[33][14][5] + xor_out[34][14][5];
assign sum_out[7][14][5] = xor_out[35][14][5] + xor_out[36][14][5] + xor_out[37][14][5] + xor_out[38][14][5] + xor_out[39][14][5];
assign sum_out[8][14][5] = xor_out[40][14][5] + xor_out[41][14][5] + xor_out[42][14][5] + xor_out[43][14][5] + xor_out[44][14][5];
assign sum_out[9][14][5] = xor_out[45][14][5] + xor_out[46][14][5] + xor_out[47][14][5] + xor_out[48][14][5] + xor_out[49][14][5];
assign sum_out[10][14][5] = xor_out[50][14][5] + xor_out[51][14][5] + xor_out[52][14][5] + xor_out[53][14][5] + xor_out[54][14][5];
assign sum_out[11][14][5] = xor_out[55][14][5] + xor_out[56][14][5] + xor_out[57][14][5] + xor_out[58][14][5] + xor_out[59][14][5];
assign sum_out[12][14][5] = xor_out[60][14][5] + xor_out[61][14][5] + xor_out[62][14][5] + xor_out[63][14][5] + xor_out[64][14][5];
assign sum_out[13][14][5] = xor_out[65][14][5] + xor_out[66][14][5] + xor_out[67][14][5] + xor_out[68][14][5] + xor_out[69][14][5];
assign sum_out[14][14][5] = xor_out[70][14][5] + xor_out[71][14][5] + xor_out[72][14][5] + xor_out[73][14][5] + xor_out[74][14][5];
assign sum_out[15][14][5] = xor_out[75][14][5] + xor_out[76][14][5] + xor_out[77][14][5] + xor_out[78][14][5] + xor_out[79][14][5];
assign sum_out[16][14][5] = xor_out[80][14][5] + xor_out[81][14][5] + xor_out[82][14][5] + xor_out[83][14][5] + xor_out[84][14][5];
assign sum_out[17][14][5] = xor_out[85][14][5] + xor_out[86][14][5] + xor_out[87][14][5] + xor_out[88][14][5] + xor_out[89][14][5];
assign sum_out[18][14][5] = xor_out[90][14][5] + xor_out[91][14][5] + xor_out[92][14][5] + xor_out[93][14][5] + xor_out[94][14][5];
assign sum_out[19][14][5] = xor_out[95][14][5] + xor_out[96][14][5] + xor_out[97][14][5] + xor_out[98][14][5] + xor_out[99][14][5];

assign sum_out[0][14][6] = xor_out[0][14][6] + xor_out[1][14][6] + xor_out[2][14][6] + xor_out[3][14][6] + xor_out[4][14][6];
assign sum_out[1][14][6] = xor_out[5][14][6] + xor_out[6][14][6] + xor_out[7][14][6] + xor_out[8][14][6] + xor_out[9][14][6];
assign sum_out[2][14][6] = xor_out[10][14][6] + xor_out[11][14][6] + xor_out[12][14][6] + xor_out[13][14][6] + xor_out[14][14][6];
assign sum_out[3][14][6] = xor_out[15][14][6] + xor_out[16][14][6] + xor_out[17][14][6] + xor_out[18][14][6] + xor_out[19][14][6];
assign sum_out[4][14][6] = xor_out[20][14][6] + xor_out[21][14][6] + xor_out[22][14][6] + xor_out[23][14][6] + xor_out[24][14][6];
assign sum_out[5][14][6] = xor_out[25][14][6] + xor_out[26][14][6] + xor_out[27][14][6] + xor_out[28][14][6] + xor_out[29][14][6];
assign sum_out[6][14][6] = xor_out[30][14][6] + xor_out[31][14][6] + xor_out[32][14][6] + xor_out[33][14][6] + xor_out[34][14][6];
assign sum_out[7][14][6] = xor_out[35][14][6] + xor_out[36][14][6] + xor_out[37][14][6] + xor_out[38][14][6] + xor_out[39][14][6];
assign sum_out[8][14][6] = xor_out[40][14][6] + xor_out[41][14][6] + xor_out[42][14][6] + xor_out[43][14][6] + xor_out[44][14][6];
assign sum_out[9][14][6] = xor_out[45][14][6] + xor_out[46][14][6] + xor_out[47][14][6] + xor_out[48][14][6] + xor_out[49][14][6];
assign sum_out[10][14][6] = xor_out[50][14][6] + xor_out[51][14][6] + xor_out[52][14][6] + xor_out[53][14][6] + xor_out[54][14][6];
assign sum_out[11][14][6] = xor_out[55][14][6] + xor_out[56][14][6] + xor_out[57][14][6] + xor_out[58][14][6] + xor_out[59][14][6];
assign sum_out[12][14][6] = xor_out[60][14][6] + xor_out[61][14][6] + xor_out[62][14][6] + xor_out[63][14][6] + xor_out[64][14][6];
assign sum_out[13][14][6] = xor_out[65][14][6] + xor_out[66][14][6] + xor_out[67][14][6] + xor_out[68][14][6] + xor_out[69][14][6];
assign sum_out[14][14][6] = xor_out[70][14][6] + xor_out[71][14][6] + xor_out[72][14][6] + xor_out[73][14][6] + xor_out[74][14][6];
assign sum_out[15][14][6] = xor_out[75][14][6] + xor_out[76][14][6] + xor_out[77][14][6] + xor_out[78][14][6] + xor_out[79][14][6];
assign sum_out[16][14][6] = xor_out[80][14][6] + xor_out[81][14][6] + xor_out[82][14][6] + xor_out[83][14][6] + xor_out[84][14][6];
assign sum_out[17][14][6] = xor_out[85][14][6] + xor_out[86][14][6] + xor_out[87][14][6] + xor_out[88][14][6] + xor_out[89][14][6];
assign sum_out[18][14][6] = xor_out[90][14][6] + xor_out[91][14][6] + xor_out[92][14][6] + xor_out[93][14][6] + xor_out[94][14][6];
assign sum_out[19][14][6] = xor_out[95][14][6] + xor_out[96][14][6] + xor_out[97][14][6] + xor_out[98][14][6] + xor_out[99][14][6];

assign sum_out[0][14][7] = xor_out[0][14][7] + xor_out[1][14][7] + xor_out[2][14][7] + xor_out[3][14][7] + xor_out[4][14][7];
assign sum_out[1][14][7] = xor_out[5][14][7] + xor_out[6][14][7] + xor_out[7][14][7] + xor_out[8][14][7] + xor_out[9][14][7];
assign sum_out[2][14][7] = xor_out[10][14][7] + xor_out[11][14][7] + xor_out[12][14][7] + xor_out[13][14][7] + xor_out[14][14][7];
assign sum_out[3][14][7] = xor_out[15][14][7] + xor_out[16][14][7] + xor_out[17][14][7] + xor_out[18][14][7] + xor_out[19][14][7];
assign sum_out[4][14][7] = xor_out[20][14][7] + xor_out[21][14][7] + xor_out[22][14][7] + xor_out[23][14][7] + xor_out[24][14][7];
assign sum_out[5][14][7] = xor_out[25][14][7] + xor_out[26][14][7] + xor_out[27][14][7] + xor_out[28][14][7] + xor_out[29][14][7];
assign sum_out[6][14][7] = xor_out[30][14][7] + xor_out[31][14][7] + xor_out[32][14][7] + xor_out[33][14][7] + xor_out[34][14][7];
assign sum_out[7][14][7] = xor_out[35][14][7] + xor_out[36][14][7] + xor_out[37][14][7] + xor_out[38][14][7] + xor_out[39][14][7];
assign sum_out[8][14][7] = xor_out[40][14][7] + xor_out[41][14][7] + xor_out[42][14][7] + xor_out[43][14][7] + xor_out[44][14][7];
assign sum_out[9][14][7] = xor_out[45][14][7] + xor_out[46][14][7] + xor_out[47][14][7] + xor_out[48][14][7] + xor_out[49][14][7];
assign sum_out[10][14][7] = xor_out[50][14][7] + xor_out[51][14][7] + xor_out[52][14][7] + xor_out[53][14][7] + xor_out[54][14][7];
assign sum_out[11][14][7] = xor_out[55][14][7] + xor_out[56][14][7] + xor_out[57][14][7] + xor_out[58][14][7] + xor_out[59][14][7];
assign sum_out[12][14][7] = xor_out[60][14][7] + xor_out[61][14][7] + xor_out[62][14][7] + xor_out[63][14][7] + xor_out[64][14][7];
assign sum_out[13][14][7] = xor_out[65][14][7] + xor_out[66][14][7] + xor_out[67][14][7] + xor_out[68][14][7] + xor_out[69][14][7];
assign sum_out[14][14][7] = xor_out[70][14][7] + xor_out[71][14][7] + xor_out[72][14][7] + xor_out[73][14][7] + xor_out[74][14][7];
assign sum_out[15][14][7] = xor_out[75][14][7] + xor_out[76][14][7] + xor_out[77][14][7] + xor_out[78][14][7] + xor_out[79][14][7];
assign sum_out[16][14][7] = xor_out[80][14][7] + xor_out[81][14][7] + xor_out[82][14][7] + xor_out[83][14][7] + xor_out[84][14][7];
assign sum_out[17][14][7] = xor_out[85][14][7] + xor_out[86][14][7] + xor_out[87][14][7] + xor_out[88][14][7] + xor_out[89][14][7];
assign sum_out[18][14][7] = xor_out[90][14][7] + xor_out[91][14][7] + xor_out[92][14][7] + xor_out[93][14][7] + xor_out[94][14][7];
assign sum_out[19][14][7] = xor_out[95][14][7] + xor_out[96][14][7] + xor_out[97][14][7] + xor_out[98][14][7] + xor_out[99][14][7];

assign sum_out[0][14][8] = xor_out[0][14][8] + xor_out[1][14][8] + xor_out[2][14][8] + xor_out[3][14][8] + xor_out[4][14][8];
assign sum_out[1][14][8] = xor_out[5][14][8] + xor_out[6][14][8] + xor_out[7][14][8] + xor_out[8][14][8] + xor_out[9][14][8];
assign sum_out[2][14][8] = xor_out[10][14][8] + xor_out[11][14][8] + xor_out[12][14][8] + xor_out[13][14][8] + xor_out[14][14][8];
assign sum_out[3][14][8] = xor_out[15][14][8] + xor_out[16][14][8] + xor_out[17][14][8] + xor_out[18][14][8] + xor_out[19][14][8];
assign sum_out[4][14][8] = xor_out[20][14][8] + xor_out[21][14][8] + xor_out[22][14][8] + xor_out[23][14][8] + xor_out[24][14][8];
assign sum_out[5][14][8] = xor_out[25][14][8] + xor_out[26][14][8] + xor_out[27][14][8] + xor_out[28][14][8] + xor_out[29][14][8];
assign sum_out[6][14][8] = xor_out[30][14][8] + xor_out[31][14][8] + xor_out[32][14][8] + xor_out[33][14][8] + xor_out[34][14][8];
assign sum_out[7][14][8] = xor_out[35][14][8] + xor_out[36][14][8] + xor_out[37][14][8] + xor_out[38][14][8] + xor_out[39][14][8];
assign sum_out[8][14][8] = xor_out[40][14][8] + xor_out[41][14][8] + xor_out[42][14][8] + xor_out[43][14][8] + xor_out[44][14][8];
assign sum_out[9][14][8] = xor_out[45][14][8] + xor_out[46][14][8] + xor_out[47][14][8] + xor_out[48][14][8] + xor_out[49][14][8];
assign sum_out[10][14][8] = xor_out[50][14][8] + xor_out[51][14][8] + xor_out[52][14][8] + xor_out[53][14][8] + xor_out[54][14][8];
assign sum_out[11][14][8] = xor_out[55][14][8] + xor_out[56][14][8] + xor_out[57][14][8] + xor_out[58][14][8] + xor_out[59][14][8];
assign sum_out[12][14][8] = xor_out[60][14][8] + xor_out[61][14][8] + xor_out[62][14][8] + xor_out[63][14][8] + xor_out[64][14][8];
assign sum_out[13][14][8] = xor_out[65][14][8] + xor_out[66][14][8] + xor_out[67][14][8] + xor_out[68][14][8] + xor_out[69][14][8];
assign sum_out[14][14][8] = xor_out[70][14][8] + xor_out[71][14][8] + xor_out[72][14][8] + xor_out[73][14][8] + xor_out[74][14][8];
assign sum_out[15][14][8] = xor_out[75][14][8] + xor_out[76][14][8] + xor_out[77][14][8] + xor_out[78][14][8] + xor_out[79][14][8];
assign sum_out[16][14][8] = xor_out[80][14][8] + xor_out[81][14][8] + xor_out[82][14][8] + xor_out[83][14][8] + xor_out[84][14][8];
assign sum_out[17][14][8] = xor_out[85][14][8] + xor_out[86][14][8] + xor_out[87][14][8] + xor_out[88][14][8] + xor_out[89][14][8];
assign sum_out[18][14][8] = xor_out[90][14][8] + xor_out[91][14][8] + xor_out[92][14][8] + xor_out[93][14][8] + xor_out[94][14][8];
assign sum_out[19][14][8] = xor_out[95][14][8] + xor_out[96][14][8] + xor_out[97][14][8] + xor_out[98][14][8] + xor_out[99][14][8];

assign sum_out[0][14][9] = xor_out[0][14][9] + xor_out[1][14][9] + xor_out[2][14][9] + xor_out[3][14][9] + xor_out[4][14][9];
assign sum_out[1][14][9] = xor_out[5][14][9] + xor_out[6][14][9] + xor_out[7][14][9] + xor_out[8][14][9] + xor_out[9][14][9];
assign sum_out[2][14][9] = xor_out[10][14][9] + xor_out[11][14][9] + xor_out[12][14][9] + xor_out[13][14][9] + xor_out[14][14][9];
assign sum_out[3][14][9] = xor_out[15][14][9] + xor_out[16][14][9] + xor_out[17][14][9] + xor_out[18][14][9] + xor_out[19][14][9];
assign sum_out[4][14][9] = xor_out[20][14][9] + xor_out[21][14][9] + xor_out[22][14][9] + xor_out[23][14][9] + xor_out[24][14][9];
assign sum_out[5][14][9] = xor_out[25][14][9] + xor_out[26][14][9] + xor_out[27][14][9] + xor_out[28][14][9] + xor_out[29][14][9];
assign sum_out[6][14][9] = xor_out[30][14][9] + xor_out[31][14][9] + xor_out[32][14][9] + xor_out[33][14][9] + xor_out[34][14][9];
assign sum_out[7][14][9] = xor_out[35][14][9] + xor_out[36][14][9] + xor_out[37][14][9] + xor_out[38][14][9] + xor_out[39][14][9];
assign sum_out[8][14][9] = xor_out[40][14][9] + xor_out[41][14][9] + xor_out[42][14][9] + xor_out[43][14][9] + xor_out[44][14][9];
assign sum_out[9][14][9] = xor_out[45][14][9] + xor_out[46][14][9] + xor_out[47][14][9] + xor_out[48][14][9] + xor_out[49][14][9];
assign sum_out[10][14][9] = xor_out[50][14][9] + xor_out[51][14][9] + xor_out[52][14][9] + xor_out[53][14][9] + xor_out[54][14][9];
assign sum_out[11][14][9] = xor_out[55][14][9] + xor_out[56][14][9] + xor_out[57][14][9] + xor_out[58][14][9] + xor_out[59][14][9];
assign sum_out[12][14][9] = xor_out[60][14][9] + xor_out[61][14][9] + xor_out[62][14][9] + xor_out[63][14][9] + xor_out[64][14][9];
assign sum_out[13][14][9] = xor_out[65][14][9] + xor_out[66][14][9] + xor_out[67][14][9] + xor_out[68][14][9] + xor_out[69][14][9];
assign sum_out[14][14][9] = xor_out[70][14][9] + xor_out[71][14][9] + xor_out[72][14][9] + xor_out[73][14][9] + xor_out[74][14][9];
assign sum_out[15][14][9] = xor_out[75][14][9] + xor_out[76][14][9] + xor_out[77][14][9] + xor_out[78][14][9] + xor_out[79][14][9];
assign sum_out[16][14][9] = xor_out[80][14][9] + xor_out[81][14][9] + xor_out[82][14][9] + xor_out[83][14][9] + xor_out[84][14][9];
assign sum_out[17][14][9] = xor_out[85][14][9] + xor_out[86][14][9] + xor_out[87][14][9] + xor_out[88][14][9] + xor_out[89][14][9];
assign sum_out[18][14][9] = xor_out[90][14][9] + xor_out[91][14][9] + xor_out[92][14][9] + xor_out[93][14][9] + xor_out[94][14][9];
assign sum_out[19][14][9] = xor_out[95][14][9] + xor_out[96][14][9] + xor_out[97][14][9] + xor_out[98][14][9] + xor_out[99][14][9];

assign sum_out[0][14][10] = xor_out[0][14][10] + xor_out[1][14][10] + xor_out[2][14][10] + xor_out[3][14][10] + xor_out[4][14][10];
assign sum_out[1][14][10] = xor_out[5][14][10] + xor_out[6][14][10] + xor_out[7][14][10] + xor_out[8][14][10] + xor_out[9][14][10];
assign sum_out[2][14][10] = xor_out[10][14][10] + xor_out[11][14][10] + xor_out[12][14][10] + xor_out[13][14][10] + xor_out[14][14][10];
assign sum_out[3][14][10] = xor_out[15][14][10] + xor_out[16][14][10] + xor_out[17][14][10] + xor_out[18][14][10] + xor_out[19][14][10];
assign sum_out[4][14][10] = xor_out[20][14][10] + xor_out[21][14][10] + xor_out[22][14][10] + xor_out[23][14][10] + xor_out[24][14][10];
assign sum_out[5][14][10] = xor_out[25][14][10] + xor_out[26][14][10] + xor_out[27][14][10] + xor_out[28][14][10] + xor_out[29][14][10];
assign sum_out[6][14][10] = xor_out[30][14][10] + xor_out[31][14][10] + xor_out[32][14][10] + xor_out[33][14][10] + xor_out[34][14][10];
assign sum_out[7][14][10] = xor_out[35][14][10] + xor_out[36][14][10] + xor_out[37][14][10] + xor_out[38][14][10] + xor_out[39][14][10];
assign sum_out[8][14][10] = xor_out[40][14][10] + xor_out[41][14][10] + xor_out[42][14][10] + xor_out[43][14][10] + xor_out[44][14][10];
assign sum_out[9][14][10] = xor_out[45][14][10] + xor_out[46][14][10] + xor_out[47][14][10] + xor_out[48][14][10] + xor_out[49][14][10];
assign sum_out[10][14][10] = xor_out[50][14][10] + xor_out[51][14][10] + xor_out[52][14][10] + xor_out[53][14][10] + xor_out[54][14][10];
assign sum_out[11][14][10] = xor_out[55][14][10] + xor_out[56][14][10] + xor_out[57][14][10] + xor_out[58][14][10] + xor_out[59][14][10];
assign sum_out[12][14][10] = xor_out[60][14][10] + xor_out[61][14][10] + xor_out[62][14][10] + xor_out[63][14][10] + xor_out[64][14][10];
assign sum_out[13][14][10] = xor_out[65][14][10] + xor_out[66][14][10] + xor_out[67][14][10] + xor_out[68][14][10] + xor_out[69][14][10];
assign sum_out[14][14][10] = xor_out[70][14][10] + xor_out[71][14][10] + xor_out[72][14][10] + xor_out[73][14][10] + xor_out[74][14][10];
assign sum_out[15][14][10] = xor_out[75][14][10] + xor_out[76][14][10] + xor_out[77][14][10] + xor_out[78][14][10] + xor_out[79][14][10];
assign sum_out[16][14][10] = xor_out[80][14][10] + xor_out[81][14][10] + xor_out[82][14][10] + xor_out[83][14][10] + xor_out[84][14][10];
assign sum_out[17][14][10] = xor_out[85][14][10] + xor_out[86][14][10] + xor_out[87][14][10] + xor_out[88][14][10] + xor_out[89][14][10];
assign sum_out[18][14][10] = xor_out[90][14][10] + xor_out[91][14][10] + xor_out[92][14][10] + xor_out[93][14][10] + xor_out[94][14][10];
assign sum_out[19][14][10] = xor_out[95][14][10] + xor_out[96][14][10] + xor_out[97][14][10] + xor_out[98][14][10] + xor_out[99][14][10];

assign sum_out[0][14][11] = xor_out[0][14][11] + xor_out[1][14][11] + xor_out[2][14][11] + xor_out[3][14][11] + xor_out[4][14][11];
assign sum_out[1][14][11] = xor_out[5][14][11] + xor_out[6][14][11] + xor_out[7][14][11] + xor_out[8][14][11] + xor_out[9][14][11];
assign sum_out[2][14][11] = xor_out[10][14][11] + xor_out[11][14][11] + xor_out[12][14][11] + xor_out[13][14][11] + xor_out[14][14][11];
assign sum_out[3][14][11] = xor_out[15][14][11] + xor_out[16][14][11] + xor_out[17][14][11] + xor_out[18][14][11] + xor_out[19][14][11];
assign sum_out[4][14][11] = xor_out[20][14][11] + xor_out[21][14][11] + xor_out[22][14][11] + xor_out[23][14][11] + xor_out[24][14][11];
assign sum_out[5][14][11] = xor_out[25][14][11] + xor_out[26][14][11] + xor_out[27][14][11] + xor_out[28][14][11] + xor_out[29][14][11];
assign sum_out[6][14][11] = xor_out[30][14][11] + xor_out[31][14][11] + xor_out[32][14][11] + xor_out[33][14][11] + xor_out[34][14][11];
assign sum_out[7][14][11] = xor_out[35][14][11] + xor_out[36][14][11] + xor_out[37][14][11] + xor_out[38][14][11] + xor_out[39][14][11];
assign sum_out[8][14][11] = xor_out[40][14][11] + xor_out[41][14][11] + xor_out[42][14][11] + xor_out[43][14][11] + xor_out[44][14][11];
assign sum_out[9][14][11] = xor_out[45][14][11] + xor_out[46][14][11] + xor_out[47][14][11] + xor_out[48][14][11] + xor_out[49][14][11];
assign sum_out[10][14][11] = xor_out[50][14][11] + xor_out[51][14][11] + xor_out[52][14][11] + xor_out[53][14][11] + xor_out[54][14][11];
assign sum_out[11][14][11] = xor_out[55][14][11] + xor_out[56][14][11] + xor_out[57][14][11] + xor_out[58][14][11] + xor_out[59][14][11];
assign sum_out[12][14][11] = xor_out[60][14][11] + xor_out[61][14][11] + xor_out[62][14][11] + xor_out[63][14][11] + xor_out[64][14][11];
assign sum_out[13][14][11] = xor_out[65][14][11] + xor_out[66][14][11] + xor_out[67][14][11] + xor_out[68][14][11] + xor_out[69][14][11];
assign sum_out[14][14][11] = xor_out[70][14][11] + xor_out[71][14][11] + xor_out[72][14][11] + xor_out[73][14][11] + xor_out[74][14][11];
assign sum_out[15][14][11] = xor_out[75][14][11] + xor_out[76][14][11] + xor_out[77][14][11] + xor_out[78][14][11] + xor_out[79][14][11];
assign sum_out[16][14][11] = xor_out[80][14][11] + xor_out[81][14][11] + xor_out[82][14][11] + xor_out[83][14][11] + xor_out[84][14][11];
assign sum_out[17][14][11] = xor_out[85][14][11] + xor_out[86][14][11] + xor_out[87][14][11] + xor_out[88][14][11] + xor_out[89][14][11];
assign sum_out[18][14][11] = xor_out[90][14][11] + xor_out[91][14][11] + xor_out[92][14][11] + xor_out[93][14][11] + xor_out[94][14][11];
assign sum_out[19][14][11] = xor_out[95][14][11] + xor_out[96][14][11] + xor_out[97][14][11] + xor_out[98][14][11] + xor_out[99][14][11];

assign sum_out[0][14][12] = xor_out[0][14][12] + xor_out[1][14][12] + xor_out[2][14][12] + xor_out[3][14][12] + xor_out[4][14][12];
assign sum_out[1][14][12] = xor_out[5][14][12] + xor_out[6][14][12] + xor_out[7][14][12] + xor_out[8][14][12] + xor_out[9][14][12];
assign sum_out[2][14][12] = xor_out[10][14][12] + xor_out[11][14][12] + xor_out[12][14][12] + xor_out[13][14][12] + xor_out[14][14][12];
assign sum_out[3][14][12] = xor_out[15][14][12] + xor_out[16][14][12] + xor_out[17][14][12] + xor_out[18][14][12] + xor_out[19][14][12];
assign sum_out[4][14][12] = xor_out[20][14][12] + xor_out[21][14][12] + xor_out[22][14][12] + xor_out[23][14][12] + xor_out[24][14][12];
assign sum_out[5][14][12] = xor_out[25][14][12] + xor_out[26][14][12] + xor_out[27][14][12] + xor_out[28][14][12] + xor_out[29][14][12];
assign sum_out[6][14][12] = xor_out[30][14][12] + xor_out[31][14][12] + xor_out[32][14][12] + xor_out[33][14][12] + xor_out[34][14][12];
assign sum_out[7][14][12] = xor_out[35][14][12] + xor_out[36][14][12] + xor_out[37][14][12] + xor_out[38][14][12] + xor_out[39][14][12];
assign sum_out[8][14][12] = xor_out[40][14][12] + xor_out[41][14][12] + xor_out[42][14][12] + xor_out[43][14][12] + xor_out[44][14][12];
assign sum_out[9][14][12] = xor_out[45][14][12] + xor_out[46][14][12] + xor_out[47][14][12] + xor_out[48][14][12] + xor_out[49][14][12];
assign sum_out[10][14][12] = xor_out[50][14][12] + xor_out[51][14][12] + xor_out[52][14][12] + xor_out[53][14][12] + xor_out[54][14][12];
assign sum_out[11][14][12] = xor_out[55][14][12] + xor_out[56][14][12] + xor_out[57][14][12] + xor_out[58][14][12] + xor_out[59][14][12];
assign sum_out[12][14][12] = xor_out[60][14][12] + xor_out[61][14][12] + xor_out[62][14][12] + xor_out[63][14][12] + xor_out[64][14][12];
assign sum_out[13][14][12] = xor_out[65][14][12] + xor_out[66][14][12] + xor_out[67][14][12] + xor_out[68][14][12] + xor_out[69][14][12];
assign sum_out[14][14][12] = xor_out[70][14][12] + xor_out[71][14][12] + xor_out[72][14][12] + xor_out[73][14][12] + xor_out[74][14][12];
assign sum_out[15][14][12] = xor_out[75][14][12] + xor_out[76][14][12] + xor_out[77][14][12] + xor_out[78][14][12] + xor_out[79][14][12];
assign sum_out[16][14][12] = xor_out[80][14][12] + xor_out[81][14][12] + xor_out[82][14][12] + xor_out[83][14][12] + xor_out[84][14][12];
assign sum_out[17][14][12] = xor_out[85][14][12] + xor_out[86][14][12] + xor_out[87][14][12] + xor_out[88][14][12] + xor_out[89][14][12];
assign sum_out[18][14][12] = xor_out[90][14][12] + xor_out[91][14][12] + xor_out[92][14][12] + xor_out[93][14][12] + xor_out[94][14][12];
assign sum_out[19][14][12] = xor_out[95][14][12] + xor_out[96][14][12] + xor_out[97][14][12] + xor_out[98][14][12] + xor_out[99][14][12];

assign sum_out[0][14][13] = xor_out[0][14][13] + xor_out[1][14][13] + xor_out[2][14][13] + xor_out[3][14][13] + xor_out[4][14][13];
assign sum_out[1][14][13] = xor_out[5][14][13] + xor_out[6][14][13] + xor_out[7][14][13] + xor_out[8][14][13] + xor_out[9][14][13];
assign sum_out[2][14][13] = xor_out[10][14][13] + xor_out[11][14][13] + xor_out[12][14][13] + xor_out[13][14][13] + xor_out[14][14][13];
assign sum_out[3][14][13] = xor_out[15][14][13] + xor_out[16][14][13] + xor_out[17][14][13] + xor_out[18][14][13] + xor_out[19][14][13];
assign sum_out[4][14][13] = xor_out[20][14][13] + xor_out[21][14][13] + xor_out[22][14][13] + xor_out[23][14][13] + xor_out[24][14][13];
assign sum_out[5][14][13] = xor_out[25][14][13] + xor_out[26][14][13] + xor_out[27][14][13] + xor_out[28][14][13] + xor_out[29][14][13];
assign sum_out[6][14][13] = xor_out[30][14][13] + xor_out[31][14][13] + xor_out[32][14][13] + xor_out[33][14][13] + xor_out[34][14][13];
assign sum_out[7][14][13] = xor_out[35][14][13] + xor_out[36][14][13] + xor_out[37][14][13] + xor_out[38][14][13] + xor_out[39][14][13];
assign sum_out[8][14][13] = xor_out[40][14][13] + xor_out[41][14][13] + xor_out[42][14][13] + xor_out[43][14][13] + xor_out[44][14][13];
assign sum_out[9][14][13] = xor_out[45][14][13] + xor_out[46][14][13] + xor_out[47][14][13] + xor_out[48][14][13] + xor_out[49][14][13];
assign sum_out[10][14][13] = xor_out[50][14][13] + xor_out[51][14][13] + xor_out[52][14][13] + xor_out[53][14][13] + xor_out[54][14][13];
assign sum_out[11][14][13] = xor_out[55][14][13] + xor_out[56][14][13] + xor_out[57][14][13] + xor_out[58][14][13] + xor_out[59][14][13];
assign sum_out[12][14][13] = xor_out[60][14][13] + xor_out[61][14][13] + xor_out[62][14][13] + xor_out[63][14][13] + xor_out[64][14][13];
assign sum_out[13][14][13] = xor_out[65][14][13] + xor_out[66][14][13] + xor_out[67][14][13] + xor_out[68][14][13] + xor_out[69][14][13];
assign sum_out[14][14][13] = xor_out[70][14][13] + xor_out[71][14][13] + xor_out[72][14][13] + xor_out[73][14][13] + xor_out[74][14][13];
assign sum_out[15][14][13] = xor_out[75][14][13] + xor_out[76][14][13] + xor_out[77][14][13] + xor_out[78][14][13] + xor_out[79][14][13];
assign sum_out[16][14][13] = xor_out[80][14][13] + xor_out[81][14][13] + xor_out[82][14][13] + xor_out[83][14][13] + xor_out[84][14][13];
assign sum_out[17][14][13] = xor_out[85][14][13] + xor_out[86][14][13] + xor_out[87][14][13] + xor_out[88][14][13] + xor_out[89][14][13];
assign sum_out[18][14][13] = xor_out[90][14][13] + xor_out[91][14][13] + xor_out[92][14][13] + xor_out[93][14][13] + xor_out[94][14][13];
assign sum_out[19][14][13] = xor_out[95][14][13] + xor_out[96][14][13] + xor_out[97][14][13] + xor_out[98][14][13] + xor_out[99][14][13];

assign sum_out[0][14][14] = xor_out[0][14][14] + xor_out[1][14][14] + xor_out[2][14][14] + xor_out[3][14][14] + xor_out[4][14][14];
assign sum_out[1][14][14] = xor_out[5][14][14] + xor_out[6][14][14] + xor_out[7][14][14] + xor_out[8][14][14] + xor_out[9][14][14];
assign sum_out[2][14][14] = xor_out[10][14][14] + xor_out[11][14][14] + xor_out[12][14][14] + xor_out[13][14][14] + xor_out[14][14][14];
assign sum_out[3][14][14] = xor_out[15][14][14] + xor_out[16][14][14] + xor_out[17][14][14] + xor_out[18][14][14] + xor_out[19][14][14];
assign sum_out[4][14][14] = xor_out[20][14][14] + xor_out[21][14][14] + xor_out[22][14][14] + xor_out[23][14][14] + xor_out[24][14][14];
assign sum_out[5][14][14] = xor_out[25][14][14] + xor_out[26][14][14] + xor_out[27][14][14] + xor_out[28][14][14] + xor_out[29][14][14];
assign sum_out[6][14][14] = xor_out[30][14][14] + xor_out[31][14][14] + xor_out[32][14][14] + xor_out[33][14][14] + xor_out[34][14][14];
assign sum_out[7][14][14] = xor_out[35][14][14] + xor_out[36][14][14] + xor_out[37][14][14] + xor_out[38][14][14] + xor_out[39][14][14];
assign sum_out[8][14][14] = xor_out[40][14][14] + xor_out[41][14][14] + xor_out[42][14][14] + xor_out[43][14][14] + xor_out[44][14][14];
assign sum_out[9][14][14] = xor_out[45][14][14] + xor_out[46][14][14] + xor_out[47][14][14] + xor_out[48][14][14] + xor_out[49][14][14];
assign sum_out[10][14][14] = xor_out[50][14][14] + xor_out[51][14][14] + xor_out[52][14][14] + xor_out[53][14][14] + xor_out[54][14][14];
assign sum_out[11][14][14] = xor_out[55][14][14] + xor_out[56][14][14] + xor_out[57][14][14] + xor_out[58][14][14] + xor_out[59][14][14];
assign sum_out[12][14][14] = xor_out[60][14][14] + xor_out[61][14][14] + xor_out[62][14][14] + xor_out[63][14][14] + xor_out[64][14][14];
assign sum_out[13][14][14] = xor_out[65][14][14] + xor_out[66][14][14] + xor_out[67][14][14] + xor_out[68][14][14] + xor_out[69][14][14];
assign sum_out[14][14][14] = xor_out[70][14][14] + xor_out[71][14][14] + xor_out[72][14][14] + xor_out[73][14][14] + xor_out[74][14][14];
assign sum_out[15][14][14] = xor_out[75][14][14] + xor_out[76][14][14] + xor_out[77][14][14] + xor_out[78][14][14] + xor_out[79][14][14];
assign sum_out[16][14][14] = xor_out[80][14][14] + xor_out[81][14][14] + xor_out[82][14][14] + xor_out[83][14][14] + xor_out[84][14][14];
assign sum_out[17][14][14] = xor_out[85][14][14] + xor_out[86][14][14] + xor_out[87][14][14] + xor_out[88][14][14] + xor_out[89][14][14];
assign sum_out[18][14][14] = xor_out[90][14][14] + xor_out[91][14][14] + xor_out[92][14][14] + xor_out[93][14][14] + xor_out[94][14][14];
assign sum_out[19][14][14] = xor_out[95][14][14] + xor_out[96][14][14] + xor_out[97][14][14] + xor_out[98][14][14] + xor_out[99][14][14];

assign sum_out[0][14][15] = xor_out[0][14][15] + xor_out[1][14][15] + xor_out[2][14][15] + xor_out[3][14][15] + xor_out[4][14][15];
assign sum_out[1][14][15] = xor_out[5][14][15] + xor_out[6][14][15] + xor_out[7][14][15] + xor_out[8][14][15] + xor_out[9][14][15];
assign sum_out[2][14][15] = xor_out[10][14][15] + xor_out[11][14][15] + xor_out[12][14][15] + xor_out[13][14][15] + xor_out[14][14][15];
assign sum_out[3][14][15] = xor_out[15][14][15] + xor_out[16][14][15] + xor_out[17][14][15] + xor_out[18][14][15] + xor_out[19][14][15];
assign sum_out[4][14][15] = xor_out[20][14][15] + xor_out[21][14][15] + xor_out[22][14][15] + xor_out[23][14][15] + xor_out[24][14][15];
assign sum_out[5][14][15] = xor_out[25][14][15] + xor_out[26][14][15] + xor_out[27][14][15] + xor_out[28][14][15] + xor_out[29][14][15];
assign sum_out[6][14][15] = xor_out[30][14][15] + xor_out[31][14][15] + xor_out[32][14][15] + xor_out[33][14][15] + xor_out[34][14][15];
assign sum_out[7][14][15] = xor_out[35][14][15] + xor_out[36][14][15] + xor_out[37][14][15] + xor_out[38][14][15] + xor_out[39][14][15];
assign sum_out[8][14][15] = xor_out[40][14][15] + xor_out[41][14][15] + xor_out[42][14][15] + xor_out[43][14][15] + xor_out[44][14][15];
assign sum_out[9][14][15] = xor_out[45][14][15] + xor_out[46][14][15] + xor_out[47][14][15] + xor_out[48][14][15] + xor_out[49][14][15];
assign sum_out[10][14][15] = xor_out[50][14][15] + xor_out[51][14][15] + xor_out[52][14][15] + xor_out[53][14][15] + xor_out[54][14][15];
assign sum_out[11][14][15] = xor_out[55][14][15] + xor_out[56][14][15] + xor_out[57][14][15] + xor_out[58][14][15] + xor_out[59][14][15];
assign sum_out[12][14][15] = xor_out[60][14][15] + xor_out[61][14][15] + xor_out[62][14][15] + xor_out[63][14][15] + xor_out[64][14][15];
assign sum_out[13][14][15] = xor_out[65][14][15] + xor_out[66][14][15] + xor_out[67][14][15] + xor_out[68][14][15] + xor_out[69][14][15];
assign sum_out[14][14][15] = xor_out[70][14][15] + xor_out[71][14][15] + xor_out[72][14][15] + xor_out[73][14][15] + xor_out[74][14][15];
assign sum_out[15][14][15] = xor_out[75][14][15] + xor_out[76][14][15] + xor_out[77][14][15] + xor_out[78][14][15] + xor_out[79][14][15];
assign sum_out[16][14][15] = xor_out[80][14][15] + xor_out[81][14][15] + xor_out[82][14][15] + xor_out[83][14][15] + xor_out[84][14][15];
assign sum_out[17][14][15] = xor_out[85][14][15] + xor_out[86][14][15] + xor_out[87][14][15] + xor_out[88][14][15] + xor_out[89][14][15];
assign sum_out[18][14][15] = xor_out[90][14][15] + xor_out[91][14][15] + xor_out[92][14][15] + xor_out[93][14][15] + xor_out[94][14][15];
assign sum_out[19][14][15] = xor_out[95][14][15] + xor_out[96][14][15] + xor_out[97][14][15] + xor_out[98][14][15] + xor_out[99][14][15];

assign sum_out[0][14][16] = xor_out[0][14][16] + xor_out[1][14][16] + xor_out[2][14][16] + xor_out[3][14][16] + xor_out[4][14][16];
assign sum_out[1][14][16] = xor_out[5][14][16] + xor_out[6][14][16] + xor_out[7][14][16] + xor_out[8][14][16] + xor_out[9][14][16];
assign sum_out[2][14][16] = xor_out[10][14][16] + xor_out[11][14][16] + xor_out[12][14][16] + xor_out[13][14][16] + xor_out[14][14][16];
assign sum_out[3][14][16] = xor_out[15][14][16] + xor_out[16][14][16] + xor_out[17][14][16] + xor_out[18][14][16] + xor_out[19][14][16];
assign sum_out[4][14][16] = xor_out[20][14][16] + xor_out[21][14][16] + xor_out[22][14][16] + xor_out[23][14][16] + xor_out[24][14][16];
assign sum_out[5][14][16] = xor_out[25][14][16] + xor_out[26][14][16] + xor_out[27][14][16] + xor_out[28][14][16] + xor_out[29][14][16];
assign sum_out[6][14][16] = xor_out[30][14][16] + xor_out[31][14][16] + xor_out[32][14][16] + xor_out[33][14][16] + xor_out[34][14][16];
assign sum_out[7][14][16] = xor_out[35][14][16] + xor_out[36][14][16] + xor_out[37][14][16] + xor_out[38][14][16] + xor_out[39][14][16];
assign sum_out[8][14][16] = xor_out[40][14][16] + xor_out[41][14][16] + xor_out[42][14][16] + xor_out[43][14][16] + xor_out[44][14][16];
assign sum_out[9][14][16] = xor_out[45][14][16] + xor_out[46][14][16] + xor_out[47][14][16] + xor_out[48][14][16] + xor_out[49][14][16];
assign sum_out[10][14][16] = xor_out[50][14][16] + xor_out[51][14][16] + xor_out[52][14][16] + xor_out[53][14][16] + xor_out[54][14][16];
assign sum_out[11][14][16] = xor_out[55][14][16] + xor_out[56][14][16] + xor_out[57][14][16] + xor_out[58][14][16] + xor_out[59][14][16];
assign sum_out[12][14][16] = xor_out[60][14][16] + xor_out[61][14][16] + xor_out[62][14][16] + xor_out[63][14][16] + xor_out[64][14][16];
assign sum_out[13][14][16] = xor_out[65][14][16] + xor_out[66][14][16] + xor_out[67][14][16] + xor_out[68][14][16] + xor_out[69][14][16];
assign sum_out[14][14][16] = xor_out[70][14][16] + xor_out[71][14][16] + xor_out[72][14][16] + xor_out[73][14][16] + xor_out[74][14][16];
assign sum_out[15][14][16] = xor_out[75][14][16] + xor_out[76][14][16] + xor_out[77][14][16] + xor_out[78][14][16] + xor_out[79][14][16];
assign sum_out[16][14][16] = xor_out[80][14][16] + xor_out[81][14][16] + xor_out[82][14][16] + xor_out[83][14][16] + xor_out[84][14][16];
assign sum_out[17][14][16] = xor_out[85][14][16] + xor_out[86][14][16] + xor_out[87][14][16] + xor_out[88][14][16] + xor_out[89][14][16];
assign sum_out[18][14][16] = xor_out[90][14][16] + xor_out[91][14][16] + xor_out[92][14][16] + xor_out[93][14][16] + xor_out[94][14][16];
assign sum_out[19][14][16] = xor_out[95][14][16] + xor_out[96][14][16] + xor_out[97][14][16] + xor_out[98][14][16] + xor_out[99][14][16];

assign sum_out[0][14][17] = xor_out[0][14][17] + xor_out[1][14][17] + xor_out[2][14][17] + xor_out[3][14][17] + xor_out[4][14][17];
assign sum_out[1][14][17] = xor_out[5][14][17] + xor_out[6][14][17] + xor_out[7][14][17] + xor_out[8][14][17] + xor_out[9][14][17];
assign sum_out[2][14][17] = xor_out[10][14][17] + xor_out[11][14][17] + xor_out[12][14][17] + xor_out[13][14][17] + xor_out[14][14][17];
assign sum_out[3][14][17] = xor_out[15][14][17] + xor_out[16][14][17] + xor_out[17][14][17] + xor_out[18][14][17] + xor_out[19][14][17];
assign sum_out[4][14][17] = xor_out[20][14][17] + xor_out[21][14][17] + xor_out[22][14][17] + xor_out[23][14][17] + xor_out[24][14][17];
assign sum_out[5][14][17] = xor_out[25][14][17] + xor_out[26][14][17] + xor_out[27][14][17] + xor_out[28][14][17] + xor_out[29][14][17];
assign sum_out[6][14][17] = xor_out[30][14][17] + xor_out[31][14][17] + xor_out[32][14][17] + xor_out[33][14][17] + xor_out[34][14][17];
assign sum_out[7][14][17] = xor_out[35][14][17] + xor_out[36][14][17] + xor_out[37][14][17] + xor_out[38][14][17] + xor_out[39][14][17];
assign sum_out[8][14][17] = xor_out[40][14][17] + xor_out[41][14][17] + xor_out[42][14][17] + xor_out[43][14][17] + xor_out[44][14][17];
assign sum_out[9][14][17] = xor_out[45][14][17] + xor_out[46][14][17] + xor_out[47][14][17] + xor_out[48][14][17] + xor_out[49][14][17];
assign sum_out[10][14][17] = xor_out[50][14][17] + xor_out[51][14][17] + xor_out[52][14][17] + xor_out[53][14][17] + xor_out[54][14][17];
assign sum_out[11][14][17] = xor_out[55][14][17] + xor_out[56][14][17] + xor_out[57][14][17] + xor_out[58][14][17] + xor_out[59][14][17];
assign sum_out[12][14][17] = xor_out[60][14][17] + xor_out[61][14][17] + xor_out[62][14][17] + xor_out[63][14][17] + xor_out[64][14][17];
assign sum_out[13][14][17] = xor_out[65][14][17] + xor_out[66][14][17] + xor_out[67][14][17] + xor_out[68][14][17] + xor_out[69][14][17];
assign sum_out[14][14][17] = xor_out[70][14][17] + xor_out[71][14][17] + xor_out[72][14][17] + xor_out[73][14][17] + xor_out[74][14][17];
assign sum_out[15][14][17] = xor_out[75][14][17] + xor_out[76][14][17] + xor_out[77][14][17] + xor_out[78][14][17] + xor_out[79][14][17];
assign sum_out[16][14][17] = xor_out[80][14][17] + xor_out[81][14][17] + xor_out[82][14][17] + xor_out[83][14][17] + xor_out[84][14][17];
assign sum_out[17][14][17] = xor_out[85][14][17] + xor_out[86][14][17] + xor_out[87][14][17] + xor_out[88][14][17] + xor_out[89][14][17];
assign sum_out[18][14][17] = xor_out[90][14][17] + xor_out[91][14][17] + xor_out[92][14][17] + xor_out[93][14][17] + xor_out[94][14][17];
assign sum_out[19][14][17] = xor_out[95][14][17] + xor_out[96][14][17] + xor_out[97][14][17] + xor_out[98][14][17] + xor_out[99][14][17];

assign sum_out[0][14][18] = xor_out[0][14][18] + xor_out[1][14][18] + xor_out[2][14][18] + xor_out[3][14][18] + xor_out[4][14][18];
assign sum_out[1][14][18] = xor_out[5][14][18] + xor_out[6][14][18] + xor_out[7][14][18] + xor_out[8][14][18] + xor_out[9][14][18];
assign sum_out[2][14][18] = xor_out[10][14][18] + xor_out[11][14][18] + xor_out[12][14][18] + xor_out[13][14][18] + xor_out[14][14][18];
assign sum_out[3][14][18] = xor_out[15][14][18] + xor_out[16][14][18] + xor_out[17][14][18] + xor_out[18][14][18] + xor_out[19][14][18];
assign sum_out[4][14][18] = xor_out[20][14][18] + xor_out[21][14][18] + xor_out[22][14][18] + xor_out[23][14][18] + xor_out[24][14][18];
assign sum_out[5][14][18] = xor_out[25][14][18] + xor_out[26][14][18] + xor_out[27][14][18] + xor_out[28][14][18] + xor_out[29][14][18];
assign sum_out[6][14][18] = xor_out[30][14][18] + xor_out[31][14][18] + xor_out[32][14][18] + xor_out[33][14][18] + xor_out[34][14][18];
assign sum_out[7][14][18] = xor_out[35][14][18] + xor_out[36][14][18] + xor_out[37][14][18] + xor_out[38][14][18] + xor_out[39][14][18];
assign sum_out[8][14][18] = xor_out[40][14][18] + xor_out[41][14][18] + xor_out[42][14][18] + xor_out[43][14][18] + xor_out[44][14][18];
assign sum_out[9][14][18] = xor_out[45][14][18] + xor_out[46][14][18] + xor_out[47][14][18] + xor_out[48][14][18] + xor_out[49][14][18];
assign sum_out[10][14][18] = xor_out[50][14][18] + xor_out[51][14][18] + xor_out[52][14][18] + xor_out[53][14][18] + xor_out[54][14][18];
assign sum_out[11][14][18] = xor_out[55][14][18] + xor_out[56][14][18] + xor_out[57][14][18] + xor_out[58][14][18] + xor_out[59][14][18];
assign sum_out[12][14][18] = xor_out[60][14][18] + xor_out[61][14][18] + xor_out[62][14][18] + xor_out[63][14][18] + xor_out[64][14][18];
assign sum_out[13][14][18] = xor_out[65][14][18] + xor_out[66][14][18] + xor_out[67][14][18] + xor_out[68][14][18] + xor_out[69][14][18];
assign sum_out[14][14][18] = xor_out[70][14][18] + xor_out[71][14][18] + xor_out[72][14][18] + xor_out[73][14][18] + xor_out[74][14][18];
assign sum_out[15][14][18] = xor_out[75][14][18] + xor_out[76][14][18] + xor_out[77][14][18] + xor_out[78][14][18] + xor_out[79][14][18];
assign sum_out[16][14][18] = xor_out[80][14][18] + xor_out[81][14][18] + xor_out[82][14][18] + xor_out[83][14][18] + xor_out[84][14][18];
assign sum_out[17][14][18] = xor_out[85][14][18] + xor_out[86][14][18] + xor_out[87][14][18] + xor_out[88][14][18] + xor_out[89][14][18];
assign sum_out[18][14][18] = xor_out[90][14][18] + xor_out[91][14][18] + xor_out[92][14][18] + xor_out[93][14][18] + xor_out[94][14][18];
assign sum_out[19][14][18] = xor_out[95][14][18] + xor_out[96][14][18] + xor_out[97][14][18] + xor_out[98][14][18] + xor_out[99][14][18];

assign sum_out[0][14][19] = xor_out[0][14][19] + xor_out[1][14][19] + xor_out[2][14][19] + xor_out[3][14][19] + xor_out[4][14][19];
assign sum_out[1][14][19] = xor_out[5][14][19] + xor_out[6][14][19] + xor_out[7][14][19] + xor_out[8][14][19] + xor_out[9][14][19];
assign sum_out[2][14][19] = xor_out[10][14][19] + xor_out[11][14][19] + xor_out[12][14][19] + xor_out[13][14][19] + xor_out[14][14][19];
assign sum_out[3][14][19] = xor_out[15][14][19] + xor_out[16][14][19] + xor_out[17][14][19] + xor_out[18][14][19] + xor_out[19][14][19];
assign sum_out[4][14][19] = xor_out[20][14][19] + xor_out[21][14][19] + xor_out[22][14][19] + xor_out[23][14][19] + xor_out[24][14][19];
assign sum_out[5][14][19] = xor_out[25][14][19] + xor_out[26][14][19] + xor_out[27][14][19] + xor_out[28][14][19] + xor_out[29][14][19];
assign sum_out[6][14][19] = xor_out[30][14][19] + xor_out[31][14][19] + xor_out[32][14][19] + xor_out[33][14][19] + xor_out[34][14][19];
assign sum_out[7][14][19] = xor_out[35][14][19] + xor_out[36][14][19] + xor_out[37][14][19] + xor_out[38][14][19] + xor_out[39][14][19];
assign sum_out[8][14][19] = xor_out[40][14][19] + xor_out[41][14][19] + xor_out[42][14][19] + xor_out[43][14][19] + xor_out[44][14][19];
assign sum_out[9][14][19] = xor_out[45][14][19] + xor_out[46][14][19] + xor_out[47][14][19] + xor_out[48][14][19] + xor_out[49][14][19];
assign sum_out[10][14][19] = xor_out[50][14][19] + xor_out[51][14][19] + xor_out[52][14][19] + xor_out[53][14][19] + xor_out[54][14][19];
assign sum_out[11][14][19] = xor_out[55][14][19] + xor_out[56][14][19] + xor_out[57][14][19] + xor_out[58][14][19] + xor_out[59][14][19];
assign sum_out[12][14][19] = xor_out[60][14][19] + xor_out[61][14][19] + xor_out[62][14][19] + xor_out[63][14][19] + xor_out[64][14][19];
assign sum_out[13][14][19] = xor_out[65][14][19] + xor_out[66][14][19] + xor_out[67][14][19] + xor_out[68][14][19] + xor_out[69][14][19];
assign sum_out[14][14][19] = xor_out[70][14][19] + xor_out[71][14][19] + xor_out[72][14][19] + xor_out[73][14][19] + xor_out[74][14][19];
assign sum_out[15][14][19] = xor_out[75][14][19] + xor_out[76][14][19] + xor_out[77][14][19] + xor_out[78][14][19] + xor_out[79][14][19];
assign sum_out[16][14][19] = xor_out[80][14][19] + xor_out[81][14][19] + xor_out[82][14][19] + xor_out[83][14][19] + xor_out[84][14][19];
assign sum_out[17][14][19] = xor_out[85][14][19] + xor_out[86][14][19] + xor_out[87][14][19] + xor_out[88][14][19] + xor_out[89][14][19];
assign sum_out[18][14][19] = xor_out[90][14][19] + xor_out[91][14][19] + xor_out[92][14][19] + xor_out[93][14][19] + xor_out[94][14][19];
assign sum_out[19][14][19] = xor_out[95][14][19] + xor_out[96][14][19] + xor_out[97][14][19] + xor_out[98][14][19] + xor_out[99][14][19];

assign sum_out[0][14][20] = xor_out[0][14][20] + xor_out[1][14][20] + xor_out[2][14][20] + xor_out[3][14][20] + xor_out[4][14][20];
assign sum_out[1][14][20] = xor_out[5][14][20] + xor_out[6][14][20] + xor_out[7][14][20] + xor_out[8][14][20] + xor_out[9][14][20];
assign sum_out[2][14][20] = xor_out[10][14][20] + xor_out[11][14][20] + xor_out[12][14][20] + xor_out[13][14][20] + xor_out[14][14][20];
assign sum_out[3][14][20] = xor_out[15][14][20] + xor_out[16][14][20] + xor_out[17][14][20] + xor_out[18][14][20] + xor_out[19][14][20];
assign sum_out[4][14][20] = xor_out[20][14][20] + xor_out[21][14][20] + xor_out[22][14][20] + xor_out[23][14][20] + xor_out[24][14][20];
assign sum_out[5][14][20] = xor_out[25][14][20] + xor_out[26][14][20] + xor_out[27][14][20] + xor_out[28][14][20] + xor_out[29][14][20];
assign sum_out[6][14][20] = xor_out[30][14][20] + xor_out[31][14][20] + xor_out[32][14][20] + xor_out[33][14][20] + xor_out[34][14][20];
assign sum_out[7][14][20] = xor_out[35][14][20] + xor_out[36][14][20] + xor_out[37][14][20] + xor_out[38][14][20] + xor_out[39][14][20];
assign sum_out[8][14][20] = xor_out[40][14][20] + xor_out[41][14][20] + xor_out[42][14][20] + xor_out[43][14][20] + xor_out[44][14][20];
assign sum_out[9][14][20] = xor_out[45][14][20] + xor_out[46][14][20] + xor_out[47][14][20] + xor_out[48][14][20] + xor_out[49][14][20];
assign sum_out[10][14][20] = xor_out[50][14][20] + xor_out[51][14][20] + xor_out[52][14][20] + xor_out[53][14][20] + xor_out[54][14][20];
assign sum_out[11][14][20] = xor_out[55][14][20] + xor_out[56][14][20] + xor_out[57][14][20] + xor_out[58][14][20] + xor_out[59][14][20];
assign sum_out[12][14][20] = xor_out[60][14][20] + xor_out[61][14][20] + xor_out[62][14][20] + xor_out[63][14][20] + xor_out[64][14][20];
assign sum_out[13][14][20] = xor_out[65][14][20] + xor_out[66][14][20] + xor_out[67][14][20] + xor_out[68][14][20] + xor_out[69][14][20];
assign sum_out[14][14][20] = xor_out[70][14][20] + xor_out[71][14][20] + xor_out[72][14][20] + xor_out[73][14][20] + xor_out[74][14][20];
assign sum_out[15][14][20] = xor_out[75][14][20] + xor_out[76][14][20] + xor_out[77][14][20] + xor_out[78][14][20] + xor_out[79][14][20];
assign sum_out[16][14][20] = xor_out[80][14][20] + xor_out[81][14][20] + xor_out[82][14][20] + xor_out[83][14][20] + xor_out[84][14][20];
assign sum_out[17][14][20] = xor_out[85][14][20] + xor_out[86][14][20] + xor_out[87][14][20] + xor_out[88][14][20] + xor_out[89][14][20];
assign sum_out[18][14][20] = xor_out[90][14][20] + xor_out[91][14][20] + xor_out[92][14][20] + xor_out[93][14][20] + xor_out[94][14][20];
assign sum_out[19][14][20] = xor_out[95][14][20] + xor_out[96][14][20] + xor_out[97][14][20] + xor_out[98][14][20] + xor_out[99][14][20];

assign sum_out[0][14][21] = xor_out[0][14][21] + xor_out[1][14][21] + xor_out[2][14][21] + xor_out[3][14][21] + xor_out[4][14][21];
assign sum_out[1][14][21] = xor_out[5][14][21] + xor_out[6][14][21] + xor_out[7][14][21] + xor_out[8][14][21] + xor_out[9][14][21];
assign sum_out[2][14][21] = xor_out[10][14][21] + xor_out[11][14][21] + xor_out[12][14][21] + xor_out[13][14][21] + xor_out[14][14][21];
assign sum_out[3][14][21] = xor_out[15][14][21] + xor_out[16][14][21] + xor_out[17][14][21] + xor_out[18][14][21] + xor_out[19][14][21];
assign sum_out[4][14][21] = xor_out[20][14][21] + xor_out[21][14][21] + xor_out[22][14][21] + xor_out[23][14][21] + xor_out[24][14][21];
assign sum_out[5][14][21] = xor_out[25][14][21] + xor_out[26][14][21] + xor_out[27][14][21] + xor_out[28][14][21] + xor_out[29][14][21];
assign sum_out[6][14][21] = xor_out[30][14][21] + xor_out[31][14][21] + xor_out[32][14][21] + xor_out[33][14][21] + xor_out[34][14][21];
assign sum_out[7][14][21] = xor_out[35][14][21] + xor_out[36][14][21] + xor_out[37][14][21] + xor_out[38][14][21] + xor_out[39][14][21];
assign sum_out[8][14][21] = xor_out[40][14][21] + xor_out[41][14][21] + xor_out[42][14][21] + xor_out[43][14][21] + xor_out[44][14][21];
assign sum_out[9][14][21] = xor_out[45][14][21] + xor_out[46][14][21] + xor_out[47][14][21] + xor_out[48][14][21] + xor_out[49][14][21];
assign sum_out[10][14][21] = xor_out[50][14][21] + xor_out[51][14][21] + xor_out[52][14][21] + xor_out[53][14][21] + xor_out[54][14][21];
assign sum_out[11][14][21] = xor_out[55][14][21] + xor_out[56][14][21] + xor_out[57][14][21] + xor_out[58][14][21] + xor_out[59][14][21];
assign sum_out[12][14][21] = xor_out[60][14][21] + xor_out[61][14][21] + xor_out[62][14][21] + xor_out[63][14][21] + xor_out[64][14][21];
assign sum_out[13][14][21] = xor_out[65][14][21] + xor_out[66][14][21] + xor_out[67][14][21] + xor_out[68][14][21] + xor_out[69][14][21];
assign sum_out[14][14][21] = xor_out[70][14][21] + xor_out[71][14][21] + xor_out[72][14][21] + xor_out[73][14][21] + xor_out[74][14][21];
assign sum_out[15][14][21] = xor_out[75][14][21] + xor_out[76][14][21] + xor_out[77][14][21] + xor_out[78][14][21] + xor_out[79][14][21];
assign sum_out[16][14][21] = xor_out[80][14][21] + xor_out[81][14][21] + xor_out[82][14][21] + xor_out[83][14][21] + xor_out[84][14][21];
assign sum_out[17][14][21] = xor_out[85][14][21] + xor_out[86][14][21] + xor_out[87][14][21] + xor_out[88][14][21] + xor_out[89][14][21];
assign sum_out[18][14][21] = xor_out[90][14][21] + xor_out[91][14][21] + xor_out[92][14][21] + xor_out[93][14][21] + xor_out[94][14][21];
assign sum_out[19][14][21] = xor_out[95][14][21] + xor_out[96][14][21] + xor_out[97][14][21] + xor_out[98][14][21] + xor_out[99][14][21];

assign sum_out[0][14][22] = xor_out[0][14][22] + xor_out[1][14][22] + xor_out[2][14][22] + xor_out[3][14][22] + xor_out[4][14][22];
assign sum_out[1][14][22] = xor_out[5][14][22] + xor_out[6][14][22] + xor_out[7][14][22] + xor_out[8][14][22] + xor_out[9][14][22];
assign sum_out[2][14][22] = xor_out[10][14][22] + xor_out[11][14][22] + xor_out[12][14][22] + xor_out[13][14][22] + xor_out[14][14][22];
assign sum_out[3][14][22] = xor_out[15][14][22] + xor_out[16][14][22] + xor_out[17][14][22] + xor_out[18][14][22] + xor_out[19][14][22];
assign sum_out[4][14][22] = xor_out[20][14][22] + xor_out[21][14][22] + xor_out[22][14][22] + xor_out[23][14][22] + xor_out[24][14][22];
assign sum_out[5][14][22] = xor_out[25][14][22] + xor_out[26][14][22] + xor_out[27][14][22] + xor_out[28][14][22] + xor_out[29][14][22];
assign sum_out[6][14][22] = xor_out[30][14][22] + xor_out[31][14][22] + xor_out[32][14][22] + xor_out[33][14][22] + xor_out[34][14][22];
assign sum_out[7][14][22] = xor_out[35][14][22] + xor_out[36][14][22] + xor_out[37][14][22] + xor_out[38][14][22] + xor_out[39][14][22];
assign sum_out[8][14][22] = xor_out[40][14][22] + xor_out[41][14][22] + xor_out[42][14][22] + xor_out[43][14][22] + xor_out[44][14][22];
assign sum_out[9][14][22] = xor_out[45][14][22] + xor_out[46][14][22] + xor_out[47][14][22] + xor_out[48][14][22] + xor_out[49][14][22];
assign sum_out[10][14][22] = xor_out[50][14][22] + xor_out[51][14][22] + xor_out[52][14][22] + xor_out[53][14][22] + xor_out[54][14][22];
assign sum_out[11][14][22] = xor_out[55][14][22] + xor_out[56][14][22] + xor_out[57][14][22] + xor_out[58][14][22] + xor_out[59][14][22];
assign sum_out[12][14][22] = xor_out[60][14][22] + xor_out[61][14][22] + xor_out[62][14][22] + xor_out[63][14][22] + xor_out[64][14][22];
assign sum_out[13][14][22] = xor_out[65][14][22] + xor_out[66][14][22] + xor_out[67][14][22] + xor_out[68][14][22] + xor_out[69][14][22];
assign sum_out[14][14][22] = xor_out[70][14][22] + xor_out[71][14][22] + xor_out[72][14][22] + xor_out[73][14][22] + xor_out[74][14][22];
assign sum_out[15][14][22] = xor_out[75][14][22] + xor_out[76][14][22] + xor_out[77][14][22] + xor_out[78][14][22] + xor_out[79][14][22];
assign sum_out[16][14][22] = xor_out[80][14][22] + xor_out[81][14][22] + xor_out[82][14][22] + xor_out[83][14][22] + xor_out[84][14][22];
assign sum_out[17][14][22] = xor_out[85][14][22] + xor_out[86][14][22] + xor_out[87][14][22] + xor_out[88][14][22] + xor_out[89][14][22];
assign sum_out[18][14][22] = xor_out[90][14][22] + xor_out[91][14][22] + xor_out[92][14][22] + xor_out[93][14][22] + xor_out[94][14][22];
assign sum_out[19][14][22] = xor_out[95][14][22] + xor_out[96][14][22] + xor_out[97][14][22] + xor_out[98][14][22] + xor_out[99][14][22];

assign sum_out[0][14][23] = xor_out[0][14][23] + xor_out[1][14][23] + xor_out[2][14][23] + xor_out[3][14][23] + xor_out[4][14][23];
assign sum_out[1][14][23] = xor_out[5][14][23] + xor_out[6][14][23] + xor_out[7][14][23] + xor_out[8][14][23] + xor_out[9][14][23];
assign sum_out[2][14][23] = xor_out[10][14][23] + xor_out[11][14][23] + xor_out[12][14][23] + xor_out[13][14][23] + xor_out[14][14][23];
assign sum_out[3][14][23] = xor_out[15][14][23] + xor_out[16][14][23] + xor_out[17][14][23] + xor_out[18][14][23] + xor_out[19][14][23];
assign sum_out[4][14][23] = xor_out[20][14][23] + xor_out[21][14][23] + xor_out[22][14][23] + xor_out[23][14][23] + xor_out[24][14][23];
assign sum_out[5][14][23] = xor_out[25][14][23] + xor_out[26][14][23] + xor_out[27][14][23] + xor_out[28][14][23] + xor_out[29][14][23];
assign sum_out[6][14][23] = xor_out[30][14][23] + xor_out[31][14][23] + xor_out[32][14][23] + xor_out[33][14][23] + xor_out[34][14][23];
assign sum_out[7][14][23] = xor_out[35][14][23] + xor_out[36][14][23] + xor_out[37][14][23] + xor_out[38][14][23] + xor_out[39][14][23];
assign sum_out[8][14][23] = xor_out[40][14][23] + xor_out[41][14][23] + xor_out[42][14][23] + xor_out[43][14][23] + xor_out[44][14][23];
assign sum_out[9][14][23] = xor_out[45][14][23] + xor_out[46][14][23] + xor_out[47][14][23] + xor_out[48][14][23] + xor_out[49][14][23];
assign sum_out[10][14][23] = xor_out[50][14][23] + xor_out[51][14][23] + xor_out[52][14][23] + xor_out[53][14][23] + xor_out[54][14][23];
assign sum_out[11][14][23] = xor_out[55][14][23] + xor_out[56][14][23] + xor_out[57][14][23] + xor_out[58][14][23] + xor_out[59][14][23];
assign sum_out[12][14][23] = xor_out[60][14][23] + xor_out[61][14][23] + xor_out[62][14][23] + xor_out[63][14][23] + xor_out[64][14][23];
assign sum_out[13][14][23] = xor_out[65][14][23] + xor_out[66][14][23] + xor_out[67][14][23] + xor_out[68][14][23] + xor_out[69][14][23];
assign sum_out[14][14][23] = xor_out[70][14][23] + xor_out[71][14][23] + xor_out[72][14][23] + xor_out[73][14][23] + xor_out[74][14][23];
assign sum_out[15][14][23] = xor_out[75][14][23] + xor_out[76][14][23] + xor_out[77][14][23] + xor_out[78][14][23] + xor_out[79][14][23];
assign sum_out[16][14][23] = xor_out[80][14][23] + xor_out[81][14][23] + xor_out[82][14][23] + xor_out[83][14][23] + xor_out[84][14][23];
assign sum_out[17][14][23] = xor_out[85][14][23] + xor_out[86][14][23] + xor_out[87][14][23] + xor_out[88][14][23] + xor_out[89][14][23];
assign sum_out[18][14][23] = xor_out[90][14][23] + xor_out[91][14][23] + xor_out[92][14][23] + xor_out[93][14][23] + xor_out[94][14][23];
assign sum_out[19][14][23] = xor_out[95][14][23] + xor_out[96][14][23] + xor_out[97][14][23] + xor_out[98][14][23] + xor_out[99][14][23];

assign sum_out[0][15][0] = xor_out[0][15][0] + xor_out[1][15][0] + xor_out[2][15][0] + xor_out[3][15][0] + xor_out[4][15][0];
assign sum_out[1][15][0] = xor_out[5][15][0] + xor_out[6][15][0] + xor_out[7][15][0] + xor_out[8][15][0] + xor_out[9][15][0];
assign sum_out[2][15][0] = xor_out[10][15][0] + xor_out[11][15][0] + xor_out[12][15][0] + xor_out[13][15][0] + xor_out[14][15][0];
assign sum_out[3][15][0] = xor_out[15][15][0] + xor_out[16][15][0] + xor_out[17][15][0] + xor_out[18][15][0] + xor_out[19][15][0];
assign sum_out[4][15][0] = xor_out[20][15][0] + xor_out[21][15][0] + xor_out[22][15][0] + xor_out[23][15][0] + xor_out[24][15][0];
assign sum_out[5][15][0] = xor_out[25][15][0] + xor_out[26][15][0] + xor_out[27][15][0] + xor_out[28][15][0] + xor_out[29][15][0];
assign sum_out[6][15][0] = xor_out[30][15][0] + xor_out[31][15][0] + xor_out[32][15][0] + xor_out[33][15][0] + xor_out[34][15][0];
assign sum_out[7][15][0] = xor_out[35][15][0] + xor_out[36][15][0] + xor_out[37][15][0] + xor_out[38][15][0] + xor_out[39][15][0];
assign sum_out[8][15][0] = xor_out[40][15][0] + xor_out[41][15][0] + xor_out[42][15][0] + xor_out[43][15][0] + xor_out[44][15][0];
assign sum_out[9][15][0] = xor_out[45][15][0] + xor_out[46][15][0] + xor_out[47][15][0] + xor_out[48][15][0] + xor_out[49][15][0];
assign sum_out[10][15][0] = xor_out[50][15][0] + xor_out[51][15][0] + xor_out[52][15][0] + xor_out[53][15][0] + xor_out[54][15][0];
assign sum_out[11][15][0] = xor_out[55][15][0] + xor_out[56][15][0] + xor_out[57][15][0] + xor_out[58][15][0] + xor_out[59][15][0];
assign sum_out[12][15][0] = xor_out[60][15][0] + xor_out[61][15][0] + xor_out[62][15][0] + xor_out[63][15][0] + xor_out[64][15][0];
assign sum_out[13][15][0] = xor_out[65][15][0] + xor_out[66][15][0] + xor_out[67][15][0] + xor_out[68][15][0] + xor_out[69][15][0];
assign sum_out[14][15][0] = xor_out[70][15][0] + xor_out[71][15][0] + xor_out[72][15][0] + xor_out[73][15][0] + xor_out[74][15][0];
assign sum_out[15][15][0] = xor_out[75][15][0] + xor_out[76][15][0] + xor_out[77][15][0] + xor_out[78][15][0] + xor_out[79][15][0];
assign sum_out[16][15][0] = xor_out[80][15][0] + xor_out[81][15][0] + xor_out[82][15][0] + xor_out[83][15][0] + xor_out[84][15][0];
assign sum_out[17][15][0] = xor_out[85][15][0] + xor_out[86][15][0] + xor_out[87][15][0] + xor_out[88][15][0] + xor_out[89][15][0];
assign sum_out[18][15][0] = xor_out[90][15][0] + xor_out[91][15][0] + xor_out[92][15][0] + xor_out[93][15][0] + xor_out[94][15][0];
assign sum_out[19][15][0] = xor_out[95][15][0] + xor_out[96][15][0] + xor_out[97][15][0] + xor_out[98][15][0] + xor_out[99][15][0];

assign sum_out[0][15][1] = xor_out[0][15][1] + xor_out[1][15][1] + xor_out[2][15][1] + xor_out[3][15][1] + xor_out[4][15][1];
assign sum_out[1][15][1] = xor_out[5][15][1] + xor_out[6][15][1] + xor_out[7][15][1] + xor_out[8][15][1] + xor_out[9][15][1];
assign sum_out[2][15][1] = xor_out[10][15][1] + xor_out[11][15][1] + xor_out[12][15][1] + xor_out[13][15][1] + xor_out[14][15][1];
assign sum_out[3][15][1] = xor_out[15][15][1] + xor_out[16][15][1] + xor_out[17][15][1] + xor_out[18][15][1] + xor_out[19][15][1];
assign sum_out[4][15][1] = xor_out[20][15][1] + xor_out[21][15][1] + xor_out[22][15][1] + xor_out[23][15][1] + xor_out[24][15][1];
assign sum_out[5][15][1] = xor_out[25][15][1] + xor_out[26][15][1] + xor_out[27][15][1] + xor_out[28][15][1] + xor_out[29][15][1];
assign sum_out[6][15][1] = xor_out[30][15][1] + xor_out[31][15][1] + xor_out[32][15][1] + xor_out[33][15][1] + xor_out[34][15][1];
assign sum_out[7][15][1] = xor_out[35][15][1] + xor_out[36][15][1] + xor_out[37][15][1] + xor_out[38][15][1] + xor_out[39][15][1];
assign sum_out[8][15][1] = xor_out[40][15][1] + xor_out[41][15][1] + xor_out[42][15][1] + xor_out[43][15][1] + xor_out[44][15][1];
assign sum_out[9][15][1] = xor_out[45][15][1] + xor_out[46][15][1] + xor_out[47][15][1] + xor_out[48][15][1] + xor_out[49][15][1];
assign sum_out[10][15][1] = xor_out[50][15][1] + xor_out[51][15][1] + xor_out[52][15][1] + xor_out[53][15][1] + xor_out[54][15][1];
assign sum_out[11][15][1] = xor_out[55][15][1] + xor_out[56][15][1] + xor_out[57][15][1] + xor_out[58][15][1] + xor_out[59][15][1];
assign sum_out[12][15][1] = xor_out[60][15][1] + xor_out[61][15][1] + xor_out[62][15][1] + xor_out[63][15][1] + xor_out[64][15][1];
assign sum_out[13][15][1] = xor_out[65][15][1] + xor_out[66][15][1] + xor_out[67][15][1] + xor_out[68][15][1] + xor_out[69][15][1];
assign sum_out[14][15][1] = xor_out[70][15][1] + xor_out[71][15][1] + xor_out[72][15][1] + xor_out[73][15][1] + xor_out[74][15][1];
assign sum_out[15][15][1] = xor_out[75][15][1] + xor_out[76][15][1] + xor_out[77][15][1] + xor_out[78][15][1] + xor_out[79][15][1];
assign sum_out[16][15][1] = xor_out[80][15][1] + xor_out[81][15][1] + xor_out[82][15][1] + xor_out[83][15][1] + xor_out[84][15][1];
assign sum_out[17][15][1] = xor_out[85][15][1] + xor_out[86][15][1] + xor_out[87][15][1] + xor_out[88][15][1] + xor_out[89][15][1];
assign sum_out[18][15][1] = xor_out[90][15][1] + xor_out[91][15][1] + xor_out[92][15][1] + xor_out[93][15][1] + xor_out[94][15][1];
assign sum_out[19][15][1] = xor_out[95][15][1] + xor_out[96][15][1] + xor_out[97][15][1] + xor_out[98][15][1] + xor_out[99][15][1];

assign sum_out[0][15][2] = xor_out[0][15][2] + xor_out[1][15][2] + xor_out[2][15][2] + xor_out[3][15][2] + xor_out[4][15][2];
assign sum_out[1][15][2] = xor_out[5][15][2] + xor_out[6][15][2] + xor_out[7][15][2] + xor_out[8][15][2] + xor_out[9][15][2];
assign sum_out[2][15][2] = xor_out[10][15][2] + xor_out[11][15][2] + xor_out[12][15][2] + xor_out[13][15][2] + xor_out[14][15][2];
assign sum_out[3][15][2] = xor_out[15][15][2] + xor_out[16][15][2] + xor_out[17][15][2] + xor_out[18][15][2] + xor_out[19][15][2];
assign sum_out[4][15][2] = xor_out[20][15][2] + xor_out[21][15][2] + xor_out[22][15][2] + xor_out[23][15][2] + xor_out[24][15][2];
assign sum_out[5][15][2] = xor_out[25][15][2] + xor_out[26][15][2] + xor_out[27][15][2] + xor_out[28][15][2] + xor_out[29][15][2];
assign sum_out[6][15][2] = xor_out[30][15][2] + xor_out[31][15][2] + xor_out[32][15][2] + xor_out[33][15][2] + xor_out[34][15][2];
assign sum_out[7][15][2] = xor_out[35][15][2] + xor_out[36][15][2] + xor_out[37][15][2] + xor_out[38][15][2] + xor_out[39][15][2];
assign sum_out[8][15][2] = xor_out[40][15][2] + xor_out[41][15][2] + xor_out[42][15][2] + xor_out[43][15][2] + xor_out[44][15][2];
assign sum_out[9][15][2] = xor_out[45][15][2] + xor_out[46][15][2] + xor_out[47][15][2] + xor_out[48][15][2] + xor_out[49][15][2];
assign sum_out[10][15][2] = xor_out[50][15][2] + xor_out[51][15][2] + xor_out[52][15][2] + xor_out[53][15][2] + xor_out[54][15][2];
assign sum_out[11][15][2] = xor_out[55][15][2] + xor_out[56][15][2] + xor_out[57][15][2] + xor_out[58][15][2] + xor_out[59][15][2];
assign sum_out[12][15][2] = xor_out[60][15][2] + xor_out[61][15][2] + xor_out[62][15][2] + xor_out[63][15][2] + xor_out[64][15][2];
assign sum_out[13][15][2] = xor_out[65][15][2] + xor_out[66][15][2] + xor_out[67][15][2] + xor_out[68][15][2] + xor_out[69][15][2];
assign sum_out[14][15][2] = xor_out[70][15][2] + xor_out[71][15][2] + xor_out[72][15][2] + xor_out[73][15][2] + xor_out[74][15][2];
assign sum_out[15][15][2] = xor_out[75][15][2] + xor_out[76][15][2] + xor_out[77][15][2] + xor_out[78][15][2] + xor_out[79][15][2];
assign sum_out[16][15][2] = xor_out[80][15][2] + xor_out[81][15][2] + xor_out[82][15][2] + xor_out[83][15][2] + xor_out[84][15][2];
assign sum_out[17][15][2] = xor_out[85][15][2] + xor_out[86][15][2] + xor_out[87][15][2] + xor_out[88][15][2] + xor_out[89][15][2];
assign sum_out[18][15][2] = xor_out[90][15][2] + xor_out[91][15][2] + xor_out[92][15][2] + xor_out[93][15][2] + xor_out[94][15][2];
assign sum_out[19][15][2] = xor_out[95][15][2] + xor_out[96][15][2] + xor_out[97][15][2] + xor_out[98][15][2] + xor_out[99][15][2];

assign sum_out[0][15][3] = xor_out[0][15][3] + xor_out[1][15][3] + xor_out[2][15][3] + xor_out[3][15][3] + xor_out[4][15][3];
assign sum_out[1][15][3] = xor_out[5][15][3] + xor_out[6][15][3] + xor_out[7][15][3] + xor_out[8][15][3] + xor_out[9][15][3];
assign sum_out[2][15][3] = xor_out[10][15][3] + xor_out[11][15][3] + xor_out[12][15][3] + xor_out[13][15][3] + xor_out[14][15][3];
assign sum_out[3][15][3] = xor_out[15][15][3] + xor_out[16][15][3] + xor_out[17][15][3] + xor_out[18][15][3] + xor_out[19][15][3];
assign sum_out[4][15][3] = xor_out[20][15][3] + xor_out[21][15][3] + xor_out[22][15][3] + xor_out[23][15][3] + xor_out[24][15][3];
assign sum_out[5][15][3] = xor_out[25][15][3] + xor_out[26][15][3] + xor_out[27][15][3] + xor_out[28][15][3] + xor_out[29][15][3];
assign sum_out[6][15][3] = xor_out[30][15][3] + xor_out[31][15][3] + xor_out[32][15][3] + xor_out[33][15][3] + xor_out[34][15][3];
assign sum_out[7][15][3] = xor_out[35][15][3] + xor_out[36][15][3] + xor_out[37][15][3] + xor_out[38][15][3] + xor_out[39][15][3];
assign sum_out[8][15][3] = xor_out[40][15][3] + xor_out[41][15][3] + xor_out[42][15][3] + xor_out[43][15][3] + xor_out[44][15][3];
assign sum_out[9][15][3] = xor_out[45][15][3] + xor_out[46][15][3] + xor_out[47][15][3] + xor_out[48][15][3] + xor_out[49][15][3];
assign sum_out[10][15][3] = xor_out[50][15][3] + xor_out[51][15][3] + xor_out[52][15][3] + xor_out[53][15][3] + xor_out[54][15][3];
assign sum_out[11][15][3] = xor_out[55][15][3] + xor_out[56][15][3] + xor_out[57][15][3] + xor_out[58][15][3] + xor_out[59][15][3];
assign sum_out[12][15][3] = xor_out[60][15][3] + xor_out[61][15][3] + xor_out[62][15][3] + xor_out[63][15][3] + xor_out[64][15][3];
assign sum_out[13][15][3] = xor_out[65][15][3] + xor_out[66][15][3] + xor_out[67][15][3] + xor_out[68][15][3] + xor_out[69][15][3];
assign sum_out[14][15][3] = xor_out[70][15][3] + xor_out[71][15][3] + xor_out[72][15][3] + xor_out[73][15][3] + xor_out[74][15][3];
assign sum_out[15][15][3] = xor_out[75][15][3] + xor_out[76][15][3] + xor_out[77][15][3] + xor_out[78][15][3] + xor_out[79][15][3];
assign sum_out[16][15][3] = xor_out[80][15][3] + xor_out[81][15][3] + xor_out[82][15][3] + xor_out[83][15][3] + xor_out[84][15][3];
assign sum_out[17][15][3] = xor_out[85][15][3] + xor_out[86][15][3] + xor_out[87][15][3] + xor_out[88][15][3] + xor_out[89][15][3];
assign sum_out[18][15][3] = xor_out[90][15][3] + xor_out[91][15][3] + xor_out[92][15][3] + xor_out[93][15][3] + xor_out[94][15][3];
assign sum_out[19][15][3] = xor_out[95][15][3] + xor_out[96][15][3] + xor_out[97][15][3] + xor_out[98][15][3] + xor_out[99][15][3];

assign sum_out[0][15][4] = xor_out[0][15][4] + xor_out[1][15][4] + xor_out[2][15][4] + xor_out[3][15][4] + xor_out[4][15][4];
assign sum_out[1][15][4] = xor_out[5][15][4] + xor_out[6][15][4] + xor_out[7][15][4] + xor_out[8][15][4] + xor_out[9][15][4];
assign sum_out[2][15][4] = xor_out[10][15][4] + xor_out[11][15][4] + xor_out[12][15][4] + xor_out[13][15][4] + xor_out[14][15][4];
assign sum_out[3][15][4] = xor_out[15][15][4] + xor_out[16][15][4] + xor_out[17][15][4] + xor_out[18][15][4] + xor_out[19][15][4];
assign sum_out[4][15][4] = xor_out[20][15][4] + xor_out[21][15][4] + xor_out[22][15][4] + xor_out[23][15][4] + xor_out[24][15][4];
assign sum_out[5][15][4] = xor_out[25][15][4] + xor_out[26][15][4] + xor_out[27][15][4] + xor_out[28][15][4] + xor_out[29][15][4];
assign sum_out[6][15][4] = xor_out[30][15][4] + xor_out[31][15][4] + xor_out[32][15][4] + xor_out[33][15][4] + xor_out[34][15][4];
assign sum_out[7][15][4] = xor_out[35][15][4] + xor_out[36][15][4] + xor_out[37][15][4] + xor_out[38][15][4] + xor_out[39][15][4];
assign sum_out[8][15][4] = xor_out[40][15][4] + xor_out[41][15][4] + xor_out[42][15][4] + xor_out[43][15][4] + xor_out[44][15][4];
assign sum_out[9][15][4] = xor_out[45][15][4] + xor_out[46][15][4] + xor_out[47][15][4] + xor_out[48][15][4] + xor_out[49][15][4];
assign sum_out[10][15][4] = xor_out[50][15][4] + xor_out[51][15][4] + xor_out[52][15][4] + xor_out[53][15][4] + xor_out[54][15][4];
assign sum_out[11][15][4] = xor_out[55][15][4] + xor_out[56][15][4] + xor_out[57][15][4] + xor_out[58][15][4] + xor_out[59][15][4];
assign sum_out[12][15][4] = xor_out[60][15][4] + xor_out[61][15][4] + xor_out[62][15][4] + xor_out[63][15][4] + xor_out[64][15][4];
assign sum_out[13][15][4] = xor_out[65][15][4] + xor_out[66][15][4] + xor_out[67][15][4] + xor_out[68][15][4] + xor_out[69][15][4];
assign sum_out[14][15][4] = xor_out[70][15][4] + xor_out[71][15][4] + xor_out[72][15][4] + xor_out[73][15][4] + xor_out[74][15][4];
assign sum_out[15][15][4] = xor_out[75][15][4] + xor_out[76][15][4] + xor_out[77][15][4] + xor_out[78][15][4] + xor_out[79][15][4];
assign sum_out[16][15][4] = xor_out[80][15][4] + xor_out[81][15][4] + xor_out[82][15][4] + xor_out[83][15][4] + xor_out[84][15][4];
assign sum_out[17][15][4] = xor_out[85][15][4] + xor_out[86][15][4] + xor_out[87][15][4] + xor_out[88][15][4] + xor_out[89][15][4];
assign sum_out[18][15][4] = xor_out[90][15][4] + xor_out[91][15][4] + xor_out[92][15][4] + xor_out[93][15][4] + xor_out[94][15][4];
assign sum_out[19][15][4] = xor_out[95][15][4] + xor_out[96][15][4] + xor_out[97][15][4] + xor_out[98][15][4] + xor_out[99][15][4];

assign sum_out[0][15][5] = xor_out[0][15][5] + xor_out[1][15][5] + xor_out[2][15][5] + xor_out[3][15][5] + xor_out[4][15][5];
assign sum_out[1][15][5] = xor_out[5][15][5] + xor_out[6][15][5] + xor_out[7][15][5] + xor_out[8][15][5] + xor_out[9][15][5];
assign sum_out[2][15][5] = xor_out[10][15][5] + xor_out[11][15][5] + xor_out[12][15][5] + xor_out[13][15][5] + xor_out[14][15][5];
assign sum_out[3][15][5] = xor_out[15][15][5] + xor_out[16][15][5] + xor_out[17][15][5] + xor_out[18][15][5] + xor_out[19][15][5];
assign sum_out[4][15][5] = xor_out[20][15][5] + xor_out[21][15][5] + xor_out[22][15][5] + xor_out[23][15][5] + xor_out[24][15][5];
assign sum_out[5][15][5] = xor_out[25][15][5] + xor_out[26][15][5] + xor_out[27][15][5] + xor_out[28][15][5] + xor_out[29][15][5];
assign sum_out[6][15][5] = xor_out[30][15][5] + xor_out[31][15][5] + xor_out[32][15][5] + xor_out[33][15][5] + xor_out[34][15][5];
assign sum_out[7][15][5] = xor_out[35][15][5] + xor_out[36][15][5] + xor_out[37][15][5] + xor_out[38][15][5] + xor_out[39][15][5];
assign sum_out[8][15][5] = xor_out[40][15][5] + xor_out[41][15][5] + xor_out[42][15][5] + xor_out[43][15][5] + xor_out[44][15][5];
assign sum_out[9][15][5] = xor_out[45][15][5] + xor_out[46][15][5] + xor_out[47][15][5] + xor_out[48][15][5] + xor_out[49][15][5];
assign sum_out[10][15][5] = xor_out[50][15][5] + xor_out[51][15][5] + xor_out[52][15][5] + xor_out[53][15][5] + xor_out[54][15][5];
assign sum_out[11][15][5] = xor_out[55][15][5] + xor_out[56][15][5] + xor_out[57][15][5] + xor_out[58][15][5] + xor_out[59][15][5];
assign sum_out[12][15][5] = xor_out[60][15][5] + xor_out[61][15][5] + xor_out[62][15][5] + xor_out[63][15][5] + xor_out[64][15][5];
assign sum_out[13][15][5] = xor_out[65][15][5] + xor_out[66][15][5] + xor_out[67][15][5] + xor_out[68][15][5] + xor_out[69][15][5];
assign sum_out[14][15][5] = xor_out[70][15][5] + xor_out[71][15][5] + xor_out[72][15][5] + xor_out[73][15][5] + xor_out[74][15][5];
assign sum_out[15][15][5] = xor_out[75][15][5] + xor_out[76][15][5] + xor_out[77][15][5] + xor_out[78][15][5] + xor_out[79][15][5];
assign sum_out[16][15][5] = xor_out[80][15][5] + xor_out[81][15][5] + xor_out[82][15][5] + xor_out[83][15][5] + xor_out[84][15][5];
assign sum_out[17][15][5] = xor_out[85][15][5] + xor_out[86][15][5] + xor_out[87][15][5] + xor_out[88][15][5] + xor_out[89][15][5];
assign sum_out[18][15][5] = xor_out[90][15][5] + xor_out[91][15][5] + xor_out[92][15][5] + xor_out[93][15][5] + xor_out[94][15][5];
assign sum_out[19][15][5] = xor_out[95][15][5] + xor_out[96][15][5] + xor_out[97][15][5] + xor_out[98][15][5] + xor_out[99][15][5];

assign sum_out[0][15][6] = xor_out[0][15][6] + xor_out[1][15][6] + xor_out[2][15][6] + xor_out[3][15][6] + xor_out[4][15][6];
assign sum_out[1][15][6] = xor_out[5][15][6] + xor_out[6][15][6] + xor_out[7][15][6] + xor_out[8][15][6] + xor_out[9][15][6];
assign sum_out[2][15][6] = xor_out[10][15][6] + xor_out[11][15][6] + xor_out[12][15][6] + xor_out[13][15][6] + xor_out[14][15][6];
assign sum_out[3][15][6] = xor_out[15][15][6] + xor_out[16][15][6] + xor_out[17][15][6] + xor_out[18][15][6] + xor_out[19][15][6];
assign sum_out[4][15][6] = xor_out[20][15][6] + xor_out[21][15][6] + xor_out[22][15][6] + xor_out[23][15][6] + xor_out[24][15][6];
assign sum_out[5][15][6] = xor_out[25][15][6] + xor_out[26][15][6] + xor_out[27][15][6] + xor_out[28][15][6] + xor_out[29][15][6];
assign sum_out[6][15][6] = xor_out[30][15][6] + xor_out[31][15][6] + xor_out[32][15][6] + xor_out[33][15][6] + xor_out[34][15][6];
assign sum_out[7][15][6] = xor_out[35][15][6] + xor_out[36][15][6] + xor_out[37][15][6] + xor_out[38][15][6] + xor_out[39][15][6];
assign sum_out[8][15][6] = xor_out[40][15][6] + xor_out[41][15][6] + xor_out[42][15][6] + xor_out[43][15][6] + xor_out[44][15][6];
assign sum_out[9][15][6] = xor_out[45][15][6] + xor_out[46][15][6] + xor_out[47][15][6] + xor_out[48][15][6] + xor_out[49][15][6];
assign sum_out[10][15][6] = xor_out[50][15][6] + xor_out[51][15][6] + xor_out[52][15][6] + xor_out[53][15][6] + xor_out[54][15][6];
assign sum_out[11][15][6] = xor_out[55][15][6] + xor_out[56][15][6] + xor_out[57][15][6] + xor_out[58][15][6] + xor_out[59][15][6];
assign sum_out[12][15][6] = xor_out[60][15][6] + xor_out[61][15][6] + xor_out[62][15][6] + xor_out[63][15][6] + xor_out[64][15][6];
assign sum_out[13][15][6] = xor_out[65][15][6] + xor_out[66][15][6] + xor_out[67][15][6] + xor_out[68][15][6] + xor_out[69][15][6];
assign sum_out[14][15][6] = xor_out[70][15][6] + xor_out[71][15][6] + xor_out[72][15][6] + xor_out[73][15][6] + xor_out[74][15][6];
assign sum_out[15][15][6] = xor_out[75][15][6] + xor_out[76][15][6] + xor_out[77][15][6] + xor_out[78][15][6] + xor_out[79][15][6];
assign sum_out[16][15][6] = xor_out[80][15][6] + xor_out[81][15][6] + xor_out[82][15][6] + xor_out[83][15][6] + xor_out[84][15][6];
assign sum_out[17][15][6] = xor_out[85][15][6] + xor_out[86][15][6] + xor_out[87][15][6] + xor_out[88][15][6] + xor_out[89][15][6];
assign sum_out[18][15][6] = xor_out[90][15][6] + xor_out[91][15][6] + xor_out[92][15][6] + xor_out[93][15][6] + xor_out[94][15][6];
assign sum_out[19][15][6] = xor_out[95][15][6] + xor_out[96][15][6] + xor_out[97][15][6] + xor_out[98][15][6] + xor_out[99][15][6];

assign sum_out[0][15][7] = xor_out[0][15][7] + xor_out[1][15][7] + xor_out[2][15][7] + xor_out[3][15][7] + xor_out[4][15][7];
assign sum_out[1][15][7] = xor_out[5][15][7] + xor_out[6][15][7] + xor_out[7][15][7] + xor_out[8][15][7] + xor_out[9][15][7];
assign sum_out[2][15][7] = xor_out[10][15][7] + xor_out[11][15][7] + xor_out[12][15][7] + xor_out[13][15][7] + xor_out[14][15][7];
assign sum_out[3][15][7] = xor_out[15][15][7] + xor_out[16][15][7] + xor_out[17][15][7] + xor_out[18][15][7] + xor_out[19][15][7];
assign sum_out[4][15][7] = xor_out[20][15][7] + xor_out[21][15][7] + xor_out[22][15][7] + xor_out[23][15][7] + xor_out[24][15][7];
assign sum_out[5][15][7] = xor_out[25][15][7] + xor_out[26][15][7] + xor_out[27][15][7] + xor_out[28][15][7] + xor_out[29][15][7];
assign sum_out[6][15][7] = xor_out[30][15][7] + xor_out[31][15][7] + xor_out[32][15][7] + xor_out[33][15][7] + xor_out[34][15][7];
assign sum_out[7][15][7] = xor_out[35][15][7] + xor_out[36][15][7] + xor_out[37][15][7] + xor_out[38][15][7] + xor_out[39][15][7];
assign sum_out[8][15][7] = xor_out[40][15][7] + xor_out[41][15][7] + xor_out[42][15][7] + xor_out[43][15][7] + xor_out[44][15][7];
assign sum_out[9][15][7] = xor_out[45][15][7] + xor_out[46][15][7] + xor_out[47][15][7] + xor_out[48][15][7] + xor_out[49][15][7];
assign sum_out[10][15][7] = xor_out[50][15][7] + xor_out[51][15][7] + xor_out[52][15][7] + xor_out[53][15][7] + xor_out[54][15][7];
assign sum_out[11][15][7] = xor_out[55][15][7] + xor_out[56][15][7] + xor_out[57][15][7] + xor_out[58][15][7] + xor_out[59][15][7];
assign sum_out[12][15][7] = xor_out[60][15][7] + xor_out[61][15][7] + xor_out[62][15][7] + xor_out[63][15][7] + xor_out[64][15][7];
assign sum_out[13][15][7] = xor_out[65][15][7] + xor_out[66][15][7] + xor_out[67][15][7] + xor_out[68][15][7] + xor_out[69][15][7];
assign sum_out[14][15][7] = xor_out[70][15][7] + xor_out[71][15][7] + xor_out[72][15][7] + xor_out[73][15][7] + xor_out[74][15][7];
assign sum_out[15][15][7] = xor_out[75][15][7] + xor_out[76][15][7] + xor_out[77][15][7] + xor_out[78][15][7] + xor_out[79][15][7];
assign sum_out[16][15][7] = xor_out[80][15][7] + xor_out[81][15][7] + xor_out[82][15][7] + xor_out[83][15][7] + xor_out[84][15][7];
assign sum_out[17][15][7] = xor_out[85][15][7] + xor_out[86][15][7] + xor_out[87][15][7] + xor_out[88][15][7] + xor_out[89][15][7];
assign sum_out[18][15][7] = xor_out[90][15][7] + xor_out[91][15][7] + xor_out[92][15][7] + xor_out[93][15][7] + xor_out[94][15][7];
assign sum_out[19][15][7] = xor_out[95][15][7] + xor_out[96][15][7] + xor_out[97][15][7] + xor_out[98][15][7] + xor_out[99][15][7];

assign sum_out[0][15][8] = xor_out[0][15][8] + xor_out[1][15][8] + xor_out[2][15][8] + xor_out[3][15][8] + xor_out[4][15][8];
assign sum_out[1][15][8] = xor_out[5][15][8] + xor_out[6][15][8] + xor_out[7][15][8] + xor_out[8][15][8] + xor_out[9][15][8];
assign sum_out[2][15][8] = xor_out[10][15][8] + xor_out[11][15][8] + xor_out[12][15][8] + xor_out[13][15][8] + xor_out[14][15][8];
assign sum_out[3][15][8] = xor_out[15][15][8] + xor_out[16][15][8] + xor_out[17][15][8] + xor_out[18][15][8] + xor_out[19][15][8];
assign sum_out[4][15][8] = xor_out[20][15][8] + xor_out[21][15][8] + xor_out[22][15][8] + xor_out[23][15][8] + xor_out[24][15][8];
assign sum_out[5][15][8] = xor_out[25][15][8] + xor_out[26][15][8] + xor_out[27][15][8] + xor_out[28][15][8] + xor_out[29][15][8];
assign sum_out[6][15][8] = xor_out[30][15][8] + xor_out[31][15][8] + xor_out[32][15][8] + xor_out[33][15][8] + xor_out[34][15][8];
assign sum_out[7][15][8] = xor_out[35][15][8] + xor_out[36][15][8] + xor_out[37][15][8] + xor_out[38][15][8] + xor_out[39][15][8];
assign sum_out[8][15][8] = xor_out[40][15][8] + xor_out[41][15][8] + xor_out[42][15][8] + xor_out[43][15][8] + xor_out[44][15][8];
assign sum_out[9][15][8] = xor_out[45][15][8] + xor_out[46][15][8] + xor_out[47][15][8] + xor_out[48][15][8] + xor_out[49][15][8];
assign sum_out[10][15][8] = xor_out[50][15][8] + xor_out[51][15][8] + xor_out[52][15][8] + xor_out[53][15][8] + xor_out[54][15][8];
assign sum_out[11][15][8] = xor_out[55][15][8] + xor_out[56][15][8] + xor_out[57][15][8] + xor_out[58][15][8] + xor_out[59][15][8];
assign sum_out[12][15][8] = xor_out[60][15][8] + xor_out[61][15][8] + xor_out[62][15][8] + xor_out[63][15][8] + xor_out[64][15][8];
assign sum_out[13][15][8] = xor_out[65][15][8] + xor_out[66][15][8] + xor_out[67][15][8] + xor_out[68][15][8] + xor_out[69][15][8];
assign sum_out[14][15][8] = xor_out[70][15][8] + xor_out[71][15][8] + xor_out[72][15][8] + xor_out[73][15][8] + xor_out[74][15][8];
assign sum_out[15][15][8] = xor_out[75][15][8] + xor_out[76][15][8] + xor_out[77][15][8] + xor_out[78][15][8] + xor_out[79][15][8];
assign sum_out[16][15][8] = xor_out[80][15][8] + xor_out[81][15][8] + xor_out[82][15][8] + xor_out[83][15][8] + xor_out[84][15][8];
assign sum_out[17][15][8] = xor_out[85][15][8] + xor_out[86][15][8] + xor_out[87][15][8] + xor_out[88][15][8] + xor_out[89][15][8];
assign sum_out[18][15][8] = xor_out[90][15][8] + xor_out[91][15][8] + xor_out[92][15][8] + xor_out[93][15][8] + xor_out[94][15][8];
assign sum_out[19][15][8] = xor_out[95][15][8] + xor_out[96][15][8] + xor_out[97][15][8] + xor_out[98][15][8] + xor_out[99][15][8];

assign sum_out[0][15][9] = xor_out[0][15][9] + xor_out[1][15][9] + xor_out[2][15][9] + xor_out[3][15][9] + xor_out[4][15][9];
assign sum_out[1][15][9] = xor_out[5][15][9] + xor_out[6][15][9] + xor_out[7][15][9] + xor_out[8][15][9] + xor_out[9][15][9];
assign sum_out[2][15][9] = xor_out[10][15][9] + xor_out[11][15][9] + xor_out[12][15][9] + xor_out[13][15][9] + xor_out[14][15][9];
assign sum_out[3][15][9] = xor_out[15][15][9] + xor_out[16][15][9] + xor_out[17][15][9] + xor_out[18][15][9] + xor_out[19][15][9];
assign sum_out[4][15][9] = xor_out[20][15][9] + xor_out[21][15][9] + xor_out[22][15][9] + xor_out[23][15][9] + xor_out[24][15][9];
assign sum_out[5][15][9] = xor_out[25][15][9] + xor_out[26][15][9] + xor_out[27][15][9] + xor_out[28][15][9] + xor_out[29][15][9];
assign sum_out[6][15][9] = xor_out[30][15][9] + xor_out[31][15][9] + xor_out[32][15][9] + xor_out[33][15][9] + xor_out[34][15][9];
assign sum_out[7][15][9] = xor_out[35][15][9] + xor_out[36][15][9] + xor_out[37][15][9] + xor_out[38][15][9] + xor_out[39][15][9];
assign sum_out[8][15][9] = xor_out[40][15][9] + xor_out[41][15][9] + xor_out[42][15][9] + xor_out[43][15][9] + xor_out[44][15][9];
assign sum_out[9][15][9] = xor_out[45][15][9] + xor_out[46][15][9] + xor_out[47][15][9] + xor_out[48][15][9] + xor_out[49][15][9];
assign sum_out[10][15][9] = xor_out[50][15][9] + xor_out[51][15][9] + xor_out[52][15][9] + xor_out[53][15][9] + xor_out[54][15][9];
assign sum_out[11][15][9] = xor_out[55][15][9] + xor_out[56][15][9] + xor_out[57][15][9] + xor_out[58][15][9] + xor_out[59][15][9];
assign sum_out[12][15][9] = xor_out[60][15][9] + xor_out[61][15][9] + xor_out[62][15][9] + xor_out[63][15][9] + xor_out[64][15][9];
assign sum_out[13][15][9] = xor_out[65][15][9] + xor_out[66][15][9] + xor_out[67][15][9] + xor_out[68][15][9] + xor_out[69][15][9];
assign sum_out[14][15][9] = xor_out[70][15][9] + xor_out[71][15][9] + xor_out[72][15][9] + xor_out[73][15][9] + xor_out[74][15][9];
assign sum_out[15][15][9] = xor_out[75][15][9] + xor_out[76][15][9] + xor_out[77][15][9] + xor_out[78][15][9] + xor_out[79][15][9];
assign sum_out[16][15][9] = xor_out[80][15][9] + xor_out[81][15][9] + xor_out[82][15][9] + xor_out[83][15][9] + xor_out[84][15][9];
assign sum_out[17][15][9] = xor_out[85][15][9] + xor_out[86][15][9] + xor_out[87][15][9] + xor_out[88][15][9] + xor_out[89][15][9];
assign sum_out[18][15][9] = xor_out[90][15][9] + xor_out[91][15][9] + xor_out[92][15][9] + xor_out[93][15][9] + xor_out[94][15][9];
assign sum_out[19][15][9] = xor_out[95][15][9] + xor_out[96][15][9] + xor_out[97][15][9] + xor_out[98][15][9] + xor_out[99][15][9];

assign sum_out[0][15][10] = xor_out[0][15][10] + xor_out[1][15][10] + xor_out[2][15][10] + xor_out[3][15][10] + xor_out[4][15][10];
assign sum_out[1][15][10] = xor_out[5][15][10] + xor_out[6][15][10] + xor_out[7][15][10] + xor_out[8][15][10] + xor_out[9][15][10];
assign sum_out[2][15][10] = xor_out[10][15][10] + xor_out[11][15][10] + xor_out[12][15][10] + xor_out[13][15][10] + xor_out[14][15][10];
assign sum_out[3][15][10] = xor_out[15][15][10] + xor_out[16][15][10] + xor_out[17][15][10] + xor_out[18][15][10] + xor_out[19][15][10];
assign sum_out[4][15][10] = xor_out[20][15][10] + xor_out[21][15][10] + xor_out[22][15][10] + xor_out[23][15][10] + xor_out[24][15][10];
assign sum_out[5][15][10] = xor_out[25][15][10] + xor_out[26][15][10] + xor_out[27][15][10] + xor_out[28][15][10] + xor_out[29][15][10];
assign sum_out[6][15][10] = xor_out[30][15][10] + xor_out[31][15][10] + xor_out[32][15][10] + xor_out[33][15][10] + xor_out[34][15][10];
assign sum_out[7][15][10] = xor_out[35][15][10] + xor_out[36][15][10] + xor_out[37][15][10] + xor_out[38][15][10] + xor_out[39][15][10];
assign sum_out[8][15][10] = xor_out[40][15][10] + xor_out[41][15][10] + xor_out[42][15][10] + xor_out[43][15][10] + xor_out[44][15][10];
assign sum_out[9][15][10] = xor_out[45][15][10] + xor_out[46][15][10] + xor_out[47][15][10] + xor_out[48][15][10] + xor_out[49][15][10];
assign sum_out[10][15][10] = xor_out[50][15][10] + xor_out[51][15][10] + xor_out[52][15][10] + xor_out[53][15][10] + xor_out[54][15][10];
assign sum_out[11][15][10] = xor_out[55][15][10] + xor_out[56][15][10] + xor_out[57][15][10] + xor_out[58][15][10] + xor_out[59][15][10];
assign sum_out[12][15][10] = xor_out[60][15][10] + xor_out[61][15][10] + xor_out[62][15][10] + xor_out[63][15][10] + xor_out[64][15][10];
assign sum_out[13][15][10] = xor_out[65][15][10] + xor_out[66][15][10] + xor_out[67][15][10] + xor_out[68][15][10] + xor_out[69][15][10];
assign sum_out[14][15][10] = xor_out[70][15][10] + xor_out[71][15][10] + xor_out[72][15][10] + xor_out[73][15][10] + xor_out[74][15][10];
assign sum_out[15][15][10] = xor_out[75][15][10] + xor_out[76][15][10] + xor_out[77][15][10] + xor_out[78][15][10] + xor_out[79][15][10];
assign sum_out[16][15][10] = xor_out[80][15][10] + xor_out[81][15][10] + xor_out[82][15][10] + xor_out[83][15][10] + xor_out[84][15][10];
assign sum_out[17][15][10] = xor_out[85][15][10] + xor_out[86][15][10] + xor_out[87][15][10] + xor_out[88][15][10] + xor_out[89][15][10];
assign sum_out[18][15][10] = xor_out[90][15][10] + xor_out[91][15][10] + xor_out[92][15][10] + xor_out[93][15][10] + xor_out[94][15][10];
assign sum_out[19][15][10] = xor_out[95][15][10] + xor_out[96][15][10] + xor_out[97][15][10] + xor_out[98][15][10] + xor_out[99][15][10];

assign sum_out[0][15][11] = xor_out[0][15][11] + xor_out[1][15][11] + xor_out[2][15][11] + xor_out[3][15][11] + xor_out[4][15][11];
assign sum_out[1][15][11] = xor_out[5][15][11] + xor_out[6][15][11] + xor_out[7][15][11] + xor_out[8][15][11] + xor_out[9][15][11];
assign sum_out[2][15][11] = xor_out[10][15][11] + xor_out[11][15][11] + xor_out[12][15][11] + xor_out[13][15][11] + xor_out[14][15][11];
assign sum_out[3][15][11] = xor_out[15][15][11] + xor_out[16][15][11] + xor_out[17][15][11] + xor_out[18][15][11] + xor_out[19][15][11];
assign sum_out[4][15][11] = xor_out[20][15][11] + xor_out[21][15][11] + xor_out[22][15][11] + xor_out[23][15][11] + xor_out[24][15][11];
assign sum_out[5][15][11] = xor_out[25][15][11] + xor_out[26][15][11] + xor_out[27][15][11] + xor_out[28][15][11] + xor_out[29][15][11];
assign sum_out[6][15][11] = xor_out[30][15][11] + xor_out[31][15][11] + xor_out[32][15][11] + xor_out[33][15][11] + xor_out[34][15][11];
assign sum_out[7][15][11] = xor_out[35][15][11] + xor_out[36][15][11] + xor_out[37][15][11] + xor_out[38][15][11] + xor_out[39][15][11];
assign sum_out[8][15][11] = xor_out[40][15][11] + xor_out[41][15][11] + xor_out[42][15][11] + xor_out[43][15][11] + xor_out[44][15][11];
assign sum_out[9][15][11] = xor_out[45][15][11] + xor_out[46][15][11] + xor_out[47][15][11] + xor_out[48][15][11] + xor_out[49][15][11];
assign sum_out[10][15][11] = xor_out[50][15][11] + xor_out[51][15][11] + xor_out[52][15][11] + xor_out[53][15][11] + xor_out[54][15][11];
assign sum_out[11][15][11] = xor_out[55][15][11] + xor_out[56][15][11] + xor_out[57][15][11] + xor_out[58][15][11] + xor_out[59][15][11];
assign sum_out[12][15][11] = xor_out[60][15][11] + xor_out[61][15][11] + xor_out[62][15][11] + xor_out[63][15][11] + xor_out[64][15][11];
assign sum_out[13][15][11] = xor_out[65][15][11] + xor_out[66][15][11] + xor_out[67][15][11] + xor_out[68][15][11] + xor_out[69][15][11];
assign sum_out[14][15][11] = xor_out[70][15][11] + xor_out[71][15][11] + xor_out[72][15][11] + xor_out[73][15][11] + xor_out[74][15][11];
assign sum_out[15][15][11] = xor_out[75][15][11] + xor_out[76][15][11] + xor_out[77][15][11] + xor_out[78][15][11] + xor_out[79][15][11];
assign sum_out[16][15][11] = xor_out[80][15][11] + xor_out[81][15][11] + xor_out[82][15][11] + xor_out[83][15][11] + xor_out[84][15][11];
assign sum_out[17][15][11] = xor_out[85][15][11] + xor_out[86][15][11] + xor_out[87][15][11] + xor_out[88][15][11] + xor_out[89][15][11];
assign sum_out[18][15][11] = xor_out[90][15][11] + xor_out[91][15][11] + xor_out[92][15][11] + xor_out[93][15][11] + xor_out[94][15][11];
assign sum_out[19][15][11] = xor_out[95][15][11] + xor_out[96][15][11] + xor_out[97][15][11] + xor_out[98][15][11] + xor_out[99][15][11];

assign sum_out[0][15][12] = xor_out[0][15][12] + xor_out[1][15][12] + xor_out[2][15][12] + xor_out[3][15][12] + xor_out[4][15][12];
assign sum_out[1][15][12] = xor_out[5][15][12] + xor_out[6][15][12] + xor_out[7][15][12] + xor_out[8][15][12] + xor_out[9][15][12];
assign sum_out[2][15][12] = xor_out[10][15][12] + xor_out[11][15][12] + xor_out[12][15][12] + xor_out[13][15][12] + xor_out[14][15][12];
assign sum_out[3][15][12] = xor_out[15][15][12] + xor_out[16][15][12] + xor_out[17][15][12] + xor_out[18][15][12] + xor_out[19][15][12];
assign sum_out[4][15][12] = xor_out[20][15][12] + xor_out[21][15][12] + xor_out[22][15][12] + xor_out[23][15][12] + xor_out[24][15][12];
assign sum_out[5][15][12] = xor_out[25][15][12] + xor_out[26][15][12] + xor_out[27][15][12] + xor_out[28][15][12] + xor_out[29][15][12];
assign sum_out[6][15][12] = xor_out[30][15][12] + xor_out[31][15][12] + xor_out[32][15][12] + xor_out[33][15][12] + xor_out[34][15][12];
assign sum_out[7][15][12] = xor_out[35][15][12] + xor_out[36][15][12] + xor_out[37][15][12] + xor_out[38][15][12] + xor_out[39][15][12];
assign sum_out[8][15][12] = xor_out[40][15][12] + xor_out[41][15][12] + xor_out[42][15][12] + xor_out[43][15][12] + xor_out[44][15][12];
assign sum_out[9][15][12] = xor_out[45][15][12] + xor_out[46][15][12] + xor_out[47][15][12] + xor_out[48][15][12] + xor_out[49][15][12];
assign sum_out[10][15][12] = xor_out[50][15][12] + xor_out[51][15][12] + xor_out[52][15][12] + xor_out[53][15][12] + xor_out[54][15][12];
assign sum_out[11][15][12] = xor_out[55][15][12] + xor_out[56][15][12] + xor_out[57][15][12] + xor_out[58][15][12] + xor_out[59][15][12];
assign sum_out[12][15][12] = xor_out[60][15][12] + xor_out[61][15][12] + xor_out[62][15][12] + xor_out[63][15][12] + xor_out[64][15][12];
assign sum_out[13][15][12] = xor_out[65][15][12] + xor_out[66][15][12] + xor_out[67][15][12] + xor_out[68][15][12] + xor_out[69][15][12];
assign sum_out[14][15][12] = xor_out[70][15][12] + xor_out[71][15][12] + xor_out[72][15][12] + xor_out[73][15][12] + xor_out[74][15][12];
assign sum_out[15][15][12] = xor_out[75][15][12] + xor_out[76][15][12] + xor_out[77][15][12] + xor_out[78][15][12] + xor_out[79][15][12];
assign sum_out[16][15][12] = xor_out[80][15][12] + xor_out[81][15][12] + xor_out[82][15][12] + xor_out[83][15][12] + xor_out[84][15][12];
assign sum_out[17][15][12] = xor_out[85][15][12] + xor_out[86][15][12] + xor_out[87][15][12] + xor_out[88][15][12] + xor_out[89][15][12];
assign sum_out[18][15][12] = xor_out[90][15][12] + xor_out[91][15][12] + xor_out[92][15][12] + xor_out[93][15][12] + xor_out[94][15][12];
assign sum_out[19][15][12] = xor_out[95][15][12] + xor_out[96][15][12] + xor_out[97][15][12] + xor_out[98][15][12] + xor_out[99][15][12];

assign sum_out[0][15][13] = xor_out[0][15][13] + xor_out[1][15][13] + xor_out[2][15][13] + xor_out[3][15][13] + xor_out[4][15][13];
assign sum_out[1][15][13] = xor_out[5][15][13] + xor_out[6][15][13] + xor_out[7][15][13] + xor_out[8][15][13] + xor_out[9][15][13];
assign sum_out[2][15][13] = xor_out[10][15][13] + xor_out[11][15][13] + xor_out[12][15][13] + xor_out[13][15][13] + xor_out[14][15][13];
assign sum_out[3][15][13] = xor_out[15][15][13] + xor_out[16][15][13] + xor_out[17][15][13] + xor_out[18][15][13] + xor_out[19][15][13];
assign sum_out[4][15][13] = xor_out[20][15][13] + xor_out[21][15][13] + xor_out[22][15][13] + xor_out[23][15][13] + xor_out[24][15][13];
assign sum_out[5][15][13] = xor_out[25][15][13] + xor_out[26][15][13] + xor_out[27][15][13] + xor_out[28][15][13] + xor_out[29][15][13];
assign sum_out[6][15][13] = xor_out[30][15][13] + xor_out[31][15][13] + xor_out[32][15][13] + xor_out[33][15][13] + xor_out[34][15][13];
assign sum_out[7][15][13] = xor_out[35][15][13] + xor_out[36][15][13] + xor_out[37][15][13] + xor_out[38][15][13] + xor_out[39][15][13];
assign sum_out[8][15][13] = xor_out[40][15][13] + xor_out[41][15][13] + xor_out[42][15][13] + xor_out[43][15][13] + xor_out[44][15][13];
assign sum_out[9][15][13] = xor_out[45][15][13] + xor_out[46][15][13] + xor_out[47][15][13] + xor_out[48][15][13] + xor_out[49][15][13];
assign sum_out[10][15][13] = xor_out[50][15][13] + xor_out[51][15][13] + xor_out[52][15][13] + xor_out[53][15][13] + xor_out[54][15][13];
assign sum_out[11][15][13] = xor_out[55][15][13] + xor_out[56][15][13] + xor_out[57][15][13] + xor_out[58][15][13] + xor_out[59][15][13];
assign sum_out[12][15][13] = xor_out[60][15][13] + xor_out[61][15][13] + xor_out[62][15][13] + xor_out[63][15][13] + xor_out[64][15][13];
assign sum_out[13][15][13] = xor_out[65][15][13] + xor_out[66][15][13] + xor_out[67][15][13] + xor_out[68][15][13] + xor_out[69][15][13];
assign sum_out[14][15][13] = xor_out[70][15][13] + xor_out[71][15][13] + xor_out[72][15][13] + xor_out[73][15][13] + xor_out[74][15][13];
assign sum_out[15][15][13] = xor_out[75][15][13] + xor_out[76][15][13] + xor_out[77][15][13] + xor_out[78][15][13] + xor_out[79][15][13];
assign sum_out[16][15][13] = xor_out[80][15][13] + xor_out[81][15][13] + xor_out[82][15][13] + xor_out[83][15][13] + xor_out[84][15][13];
assign sum_out[17][15][13] = xor_out[85][15][13] + xor_out[86][15][13] + xor_out[87][15][13] + xor_out[88][15][13] + xor_out[89][15][13];
assign sum_out[18][15][13] = xor_out[90][15][13] + xor_out[91][15][13] + xor_out[92][15][13] + xor_out[93][15][13] + xor_out[94][15][13];
assign sum_out[19][15][13] = xor_out[95][15][13] + xor_out[96][15][13] + xor_out[97][15][13] + xor_out[98][15][13] + xor_out[99][15][13];

assign sum_out[0][15][14] = xor_out[0][15][14] + xor_out[1][15][14] + xor_out[2][15][14] + xor_out[3][15][14] + xor_out[4][15][14];
assign sum_out[1][15][14] = xor_out[5][15][14] + xor_out[6][15][14] + xor_out[7][15][14] + xor_out[8][15][14] + xor_out[9][15][14];
assign sum_out[2][15][14] = xor_out[10][15][14] + xor_out[11][15][14] + xor_out[12][15][14] + xor_out[13][15][14] + xor_out[14][15][14];
assign sum_out[3][15][14] = xor_out[15][15][14] + xor_out[16][15][14] + xor_out[17][15][14] + xor_out[18][15][14] + xor_out[19][15][14];
assign sum_out[4][15][14] = xor_out[20][15][14] + xor_out[21][15][14] + xor_out[22][15][14] + xor_out[23][15][14] + xor_out[24][15][14];
assign sum_out[5][15][14] = xor_out[25][15][14] + xor_out[26][15][14] + xor_out[27][15][14] + xor_out[28][15][14] + xor_out[29][15][14];
assign sum_out[6][15][14] = xor_out[30][15][14] + xor_out[31][15][14] + xor_out[32][15][14] + xor_out[33][15][14] + xor_out[34][15][14];
assign sum_out[7][15][14] = xor_out[35][15][14] + xor_out[36][15][14] + xor_out[37][15][14] + xor_out[38][15][14] + xor_out[39][15][14];
assign sum_out[8][15][14] = xor_out[40][15][14] + xor_out[41][15][14] + xor_out[42][15][14] + xor_out[43][15][14] + xor_out[44][15][14];
assign sum_out[9][15][14] = xor_out[45][15][14] + xor_out[46][15][14] + xor_out[47][15][14] + xor_out[48][15][14] + xor_out[49][15][14];
assign sum_out[10][15][14] = xor_out[50][15][14] + xor_out[51][15][14] + xor_out[52][15][14] + xor_out[53][15][14] + xor_out[54][15][14];
assign sum_out[11][15][14] = xor_out[55][15][14] + xor_out[56][15][14] + xor_out[57][15][14] + xor_out[58][15][14] + xor_out[59][15][14];
assign sum_out[12][15][14] = xor_out[60][15][14] + xor_out[61][15][14] + xor_out[62][15][14] + xor_out[63][15][14] + xor_out[64][15][14];
assign sum_out[13][15][14] = xor_out[65][15][14] + xor_out[66][15][14] + xor_out[67][15][14] + xor_out[68][15][14] + xor_out[69][15][14];
assign sum_out[14][15][14] = xor_out[70][15][14] + xor_out[71][15][14] + xor_out[72][15][14] + xor_out[73][15][14] + xor_out[74][15][14];
assign sum_out[15][15][14] = xor_out[75][15][14] + xor_out[76][15][14] + xor_out[77][15][14] + xor_out[78][15][14] + xor_out[79][15][14];
assign sum_out[16][15][14] = xor_out[80][15][14] + xor_out[81][15][14] + xor_out[82][15][14] + xor_out[83][15][14] + xor_out[84][15][14];
assign sum_out[17][15][14] = xor_out[85][15][14] + xor_out[86][15][14] + xor_out[87][15][14] + xor_out[88][15][14] + xor_out[89][15][14];
assign sum_out[18][15][14] = xor_out[90][15][14] + xor_out[91][15][14] + xor_out[92][15][14] + xor_out[93][15][14] + xor_out[94][15][14];
assign sum_out[19][15][14] = xor_out[95][15][14] + xor_out[96][15][14] + xor_out[97][15][14] + xor_out[98][15][14] + xor_out[99][15][14];

assign sum_out[0][15][15] = xor_out[0][15][15] + xor_out[1][15][15] + xor_out[2][15][15] + xor_out[3][15][15] + xor_out[4][15][15];
assign sum_out[1][15][15] = xor_out[5][15][15] + xor_out[6][15][15] + xor_out[7][15][15] + xor_out[8][15][15] + xor_out[9][15][15];
assign sum_out[2][15][15] = xor_out[10][15][15] + xor_out[11][15][15] + xor_out[12][15][15] + xor_out[13][15][15] + xor_out[14][15][15];
assign sum_out[3][15][15] = xor_out[15][15][15] + xor_out[16][15][15] + xor_out[17][15][15] + xor_out[18][15][15] + xor_out[19][15][15];
assign sum_out[4][15][15] = xor_out[20][15][15] + xor_out[21][15][15] + xor_out[22][15][15] + xor_out[23][15][15] + xor_out[24][15][15];
assign sum_out[5][15][15] = xor_out[25][15][15] + xor_out[26][15][15] + xor_out[27][15][15] + xor_out[28][15][15] + xor_out[29][15][15];
assign sum_out[6][15][15] = xor_out[30][15][15] + xor_out[31][15][15] + xor_out[32][15][15] + xor_out[33][15][15] + xor_out[34][15][15];
assign sum_out[7][15][15] = xor_out[35][15][15] + xor_out[36][15][15] + xor_out[37][15][15] + xor_out[38][15][15] + xor_out[39][15][15];
assign sum_out[8][15][15] = xor_out[40][15][15] + xor_out[41][15][15] + xor_out[42][15][15] + xor_out[43][15][15] + xor_out[44][15][15];
assign sum_out[9][15][15] = xor_out[45][15][15] + xor_out[46][15][15] + xor_out[47][15][15] + xor_out[48][15][15] + xor_out[49][15][15];
assign sum_out[10][15][15] = xor_out[50][15][15] + xor_out[51][15][15] + xor_out[52][15][15] + xor_out[53][15][15] + xor_out[54][15][15];
assign sum_out[11][15][15] = xor_out[55][15][15] + xor_out[56][15][15] + xor_out[57][15][15] + xor_out[58][15][15] + xor_out[59][15][15];
assign sum_out[12][15][15] = xor_out[60][15][15] + xor_out[61][15][15] + xor_out[62][15][15] + xor_out[63][15][15] + xor_out[64][15][15];
assign sum_out[13][15][15] = xor_out[65][15][15] + xor_out[66][15][15] + xor_out[67][15][15] + xor_out[68][15][15] + xor_out[69][15][15];
assign sum_out[14][15][15] = xor_out[70][15][15] + xor_out[71][15][15] + xor_out[72][15][15] + xor_out[73][15][15] + xor_out[74][15][15];
assign sum_out[15][15][15] = xor_out[75][15][15] + xor_out[76][15][15] + xor_out[77][15][15] + xor_out[78][15][15] + xor_out[79][15][15];
assign sum_out[16][15][15] = xor_out[80][15][15] + xor_out[81][15][15] + xor_out[82][15][15] + xor_out[83][15][15] + xor_out[84][15][15];
assign sum_out[17][15][15] = xor_out[85][15][15] + xor_out[86][15][15] + xor_out[87][15][15] + xor_out[88][15][15] + xor_out[89][15][15];
assign sum_out[18][15][15] = xor_out[90][15][15] + xor_out[91][15][15] + xor_out[92][15][15] + xor_out[93][15][15] + xor_out[94][15][15];
assign sum_out[19][15][15] = xor_out[95][15][15] + xor_out[96][15][15] + xor_out[97][15][15] + xor_out[98][15][15] + xor_out[99][15][15];

assign sum_out[0][15][16] = xor_out[0][15][16] + xor_out[1][15][16] + xor_out[2][15][16] + xor_out[3][15][16] + xor_out[4][15][16];
assign sum_out[1][15][16] = xor_out[5][15][16] + xor_out[6][15][16] + xor_out[7][15][16] + xor_out[8][15][16] + xor_out[9][15][16];
assign sum_out[2][15][16] = xor_out[10][15][16] + xor_out[11][15][16] + xor_out[12][15][16] + xor_out[13][15][16] + xor_out[14][15][16];
assign sum_out[3][15][16] = xor_out[15][15][16] + xor_out[16][15][16] + xor_out[17][15][16] + xor_out[18][15][16] + xor_out[19][15][16];
assign sum_out[4][15][16] = xor_out[20][15][16] + xor_out[21][15][16] + xor_out[22][15][16] + xor_out[23][15][16] + xor_out[24][15][16];
assign sum_out[5][15][16] = xor_out[25][15][16] + xor_out[26][15][16] + xor_out[27][15][16] + xor_out[28][15][16] + xor_out[29][15][16];
assign sum_out[6][15][16] = xor_out[30][15][16] + xor_out[31][15][16] + xor_out[32][15][16] + xor_out[33][15][16] + xor_out[34][15][16];
assign sum_out[7][15][16] = xor_out[35][15][16] + xor_out[36][15][16] + xor_out[37][15][16] + xor_out[38][15][16] + xor_out[39][15][16];
assign sum_out[8][15][16] = xor_out[40][15][16] + xor_out[41][15][16] + xor_out[42][15][16] + xor_out[43][15][16] + xor_out[44][15][16];
assign sum_out[9][15][16] = xor_out[45][15][16] + xor_out[46][15][16] + xor_out[47][15][16] + xor_out[48][15][16] + xor_out[49][15][16];
assign sum_out[10][15][16] = xor_out[50][15][16] + xor_out[51][15][16] + xor_out[52][15][16] + xor_out[53][15][16] + xor_out[54][15][16];
assign sum_out[11][15][16] = xor_out[55][15][16] + xor_out[56][15][16] + xor_out[57][15][16] + xor_out[58][15][16] + xor_out[59][15][16];
assign sum_out[12][15][16] = xor_out[60][15][16] + xor_out[61][15][16] + xor_out[62][15][16] + xor_out[63][15][16] + xor_out[64][15][16];
assign sum_out[13][15][16] = xor_out[65][15][16] + xor_out[66][15][16] + xor_out[67][15][16] + xor_out[68][15][16] + xor_out[69][15][16];
assign sum_out[14][15][16] = xor_out[70][15][16] + xor_out[71][15][16] + xor_out[72][15][16] + xor_out[73][15][16] + xor_out[74][15][16];
assign sum_out[15][15][16] = xor_out[75][15][16] + xor_out[76][15][16] + xor_out[77][15][16] + xor_out[78][15][16] + xor_out[79][15][16];
assign sum_out[16][15][16] = xor_out[80][15][16] + xor_out[81][15][16] + xor_out[82][15][16] + xor_out[83][15][16] + xor_out[84][15][16];
assign sum_out[17][15][16] = xor_out[85][15][16] + xor_out[86][15][16] + xor_out[87][15][16] + xor_out[88][15][16] + xor_out[89][15][16];
assign sum_out[18][15][16] = xor_out[90][15][16] + xor_out[91][15][16] + xor_out[92][15][16] + xor_out[93][15][16] + xor_out[94][15][16];
assign sum_out[19][15][16] = xor_out[95][15][16] + xor_out[96][15][16] + xor_out[97][15][16] + xor_out[98][15][16] + xor_out[99][15][16];

assign sum_out[0][15][17] = xor_out[0][15][17] + xor_out[1][15][17] + xor_out[2][15][17] + xor_out[3][15][17] + xor_out[4][15][17];
assign sum_out[1][15][17] = xor_out[5][15][17] + xor_out[6][15][17] + xor_out[7][15][17] + xor_out[8][15][17] + xor_out[9][15][17];
assign sum_out[2][15][17] = xor_out[10][15][17] + xor_out[11][15][17] + xor_out[12][15][17] + xor_out[13][15][17] + xor_out[14][15][17];
assign sum_out[3][15][17] = xor_out[15][15][17] + xor_out[16][15][17] + xor_out[17][15][17] + xor_out[18][15][17] + xor_out[19][15][17];
assign sum_out[4][15][17] = xor_out[20][15][17] + xor_out[21][15][17] + xor_out[22][15][17] + xor_out[23][15][17] + xor_out[24][15][17];
assign sum_out[5][15][17] = xor_out[25][15][17] + xor_out[26][15][17] + xor_out[27][15][17] + xor_out[28][15][17] + xor_out[29][15][17];
assign sum_out[6][15][17] = xor_out[30][15][17] + xor_out[31][15][17] + xor_out[32][15][17] + xor_out[33][15][17] + xor_out[34][15][17];
assign sum_out[7][15][17] = xor_out[35][15][17] + xor_out[36][15][17] + xor_out[37][15][17] + xor_out[38][15][17] + xor_out[39][15][17];
assign sum_out[8][15][17] = xor_out[40][15][17] + xor_out[41][15][17] + xor_out[42][15][17] + xor_out[43][15][17] + xor_out[44][15][17];
assign sum_out[9][15][17] = xor_out[45][15][17] + xor_out[46][15][17] + xor_out[47][15][17] + xor_out[48][15][17] + xor_out[49][15][17];
assign sum_out[10][15][17] = xor_out[50][15][17] + xor_out[51][15][17] + xor_out[52][15][17] + xor_out[53][15][17] + xor_out[54][15][17];
assign sum_out[11][15][17] = xor_out[55][15][17] + xor_out[56][15][17] + xor_out[57][15][17] + xor_out[58][15][17] + xor_out[59][15][17];
assign sum_out[12][15][17] = xor_out[60][15][17] + xor_out[61][15][17] + xor_out[62][15][17] + xor_out[63][15][17] + xor_out[64][15][17];
assign sum_out[13][15][17] = xor_out[65][15][17] + xor_out[66][15][17] + xor_out[67][15][17] + xor_out[68][15][17] + xor_out[69][15][17];
assign sum_out[14][15][17] = xor_out[70][15][17] + xor_out[71][15][17] + xor_out[72][15][17] + xor_out[73][15][17] + xor_out[74][15][17];
assign sum_out[15][15][17] = xor_out[75][15][17] + xor_out[76][15][17] + xor_out[77][15][17] + xor_out[78][15][17] + xor_out[79][15][17];
assign sum_out[16][15][17] = xor_out[80][15][17] + xor_out[81][15][17] + xor_out[82][15][17] + xor_out[83][15][17] + xor_out[84][15][17];
assign sum_out[17][15][17] = xor_out[85][15][17] + xor_out[86][15][17] + xor_out[87][15][17] + xor_out[88][15][17] + xor_out[89][15][17];
assign sum_out[18][15][17] = xor_out[90][15][17] + xor_out[91][15][17] + xor_out[92][15][17] + xor_out[93][15][17] + xor_out[94][15][17];
assign sum_out[19][15][17] = xor_out[95][15][17] + xor_out[96][15][17] + xor_out[97][15][17] + xor_out[98][15][17] + xor_out[99][15][17];

assign sum_out[0][15][18] = xor_out[0][15][18] + xor_out[1][15][18] + xor_out[2][15][18] + xor_out[3][15][18] + xor_out[4][15][18];
assign sum_out[1][15][18] = xor_out[5][15][18] + xor_out[6][15][18] + xor_out[7][15][18] + xor_out[8][15][18] + xor_out[9][15][18];
assign sum_out[2][15][18] = xor_out[10][15][18] + xor_out[11][15][18] + xor_out[12][15][18] + xor_out[13][15][18] + xor_out[14][15][18];
assign sum_out[3][15][18] = xor_out[15][15][18] + xor_out[16][15][18] + xor_out[17][15][18] + xor_out[18][15][18] + xor_out[19][15][18];
assign sum_out[4][15][18] = xor_out[20][15][18] + xor_out[21][15][18] + xor_out[22][15][18] + xor_out[23][15][18] + xor_out[24][15][18];
assign sum_out[5][15][18] = xor_out[25][15][18] + xor_out[26][15][18] + xor_out[27][15][18] + xor_out[28][15][18] + xor_out[29][15][18];
assign sum_out[6][15][18] = xor_out[30][15][18] + xor_out[31][15][18] + xor_out[32][15][18] + xor_out[33][15][18] + xor_out[34][15][18];
assign sum_out[7][15][18] = xor_out[35][15][18] + xor_out[36][15][18] + xor_out[37][15][18] + xor_out[38][15][18] + xor_out[39][15][18];
assign sum_out[8][15][18] = xor_out[40][15][18] + xor_out[41][15][18] + xor_out[42][15][18] + xor_out[43][15][18] + xor_out[44][15][18];
assign sum_out[9][15][18] = xor_out[45][15][18] + xor_out[46][15][18] + xor_out[47][15][18] + xor_out[48][15][18] + xor_out[49][15][18];
assign sum_out[10][15][18] = xor_out[50][15][18] + xor_out[51][15][18] + xor_out[52][15][18] + xor_out[53][15][18] + xor_out[54][15][18];
assign sum_out[11][15][18] = xor_out[55][15][18] + xor_out[56][15][18] + xor_out[57][15][18] + xor_out[58][15][18] + xor_out[59][15][18];
assign sum_out[12][15][18] = xor_out[60][15][18] + xor_out[61][15][18] + xor_out[62][15][18] + xor_out[63][15][18] + xor_out[64][15][18];
assign sum_out[13][15][18] = xor_out[65][15][18] + xor_out[66][15][18] + xor_out[67][15][18] + xor_out[68][15][18] + xor_out[69][15][18];
assign sum_out[14][15][18] = xor_out[70][15][18] + xor_out[71][15][18] + xor_out[72][15][18] + xor_out[73][15][18] + xor_out[74][15][18];
assign sum_out[15][15][18] = xor_out[75][15][18] + xor_out[76][15][18] + xor_out[77][15][18] + xor_out[78][15][18] + xor_out[79][15][18];
assign sum_out[16][15][18] = xor_out[80][15][18] + xor_out[81][15][18] + xor_out[82][15][18] + xor_out[83][15][18] + xor_out[84][15][18];
assign sum_out[17][15][18] = xor_out[85][15][18] + xor_out[86][15][18] + xor_out[87][15][18] + xor_out[88][15][18] + xor_out[89][15][18];
assign sum_out[18][15][18] = xor_out[90][15][18] + xor_out[91][15][18] + xor_out[92][15][18] + xor_out[93][15][18] + xor_out[94][15][18];
assign sum_out[19][15][18] = xor_out[95][15][18] + xor_out[96][15][18] + xor_out[97][15][18] + xor_out[98][15][18] + xor_out[99][15][18];

assign sum_out[0][15][19] = xor_out[0][15][19] + xor_out[1][15][19] + xor_out[2][15][19] + xor_out[3][15][19] + xor_out[4][15][19];
assign sum_out[1][15][19] = xor_out[5][15][19] + xor_out[6][15][19] + xor_out[7][15][19] + xor_out[8][15][19] + xor_out[9][15][19];
assign sum_out[2][15][19] = xor_out[10][15][19] + xor_out[11][15][19] + xor_out[12][15][19] + xor_out[13][15][19] + xor_out[14][15][19];
assign sum_out[3][15][19] = xor_out[15][15][19] + xor_out[16][15][19] + xor_out[17][15][19] + xor_out[18][15][19] + xor_out[19][15][19];
assign sum_out[4][15][19] = xor_out[20][15][19] + xor_out[21][15][19] + xor_out[22][15][19] + xor_out[23][15][19] + xor_out[24][15][19];
assign sum_out[5][15][19] = xor_out[25][15][19] + xor_out[26][15][19] + xor_out[27][15][19] + xor_out[28][15][19] + xor_out[29][15][19];
assign sum_out[6][15][19] = xor_out[30][15][19] + xor_out[31][15][19] + xor_out[32][15][19] + xor_out[33][15][19] + xor_out[34][15][19];
assign sum_out[7][15][19] = xor_out[35][15][19] + xor_out[36][15][19] + xor_out[37][15][19] + xor_out[38][15][19] + xor_out[39][15][19];
assign sum_out[8][15][19] = xor_out[40][15][19] + xor_out[41][15][19] + xor_out[42][15][19] + xor_out[43][15][19] + xor_out[44][15][19];
assign sum_out[9][15][19] = xor_out[45][15][19] + xor_out[46][15][19] + xor_out[47][15][19] + xor_out[48][15][19] + xor_out[49][15][19];
assign sum_out[10][15][19] = xor_out[50][15][19] + xor_out[51][15][19] + xor_out[52][15][19] + xor_out[53][15][19] + xor_out[54][15][19];
assign sum_out[11][15][19] = xor_out[55][15][19] + xor_out[56][15][19] + xor_out[57][15][19] + xor_out[58][15][19] + xor_out[59][15][19];
assign sum_out[12][15][19] = xor_out[60][15][19] + xor_out[61][15][19] + xor_out[62][15][19] + xor_out[63][15][19] + xor_out[64][15][19];
assign sum_out[13][15][19] = xor_out[65][15][19] + xor_out[66][15][19] + xor_out[67][15][19] + xor_out[68][15][19] + xor_out[69][15][19];
assign sum_out[14][15][19] = xor_out[70][15][19] + xor_out[71][15][19] + xor_out[72][15][19] + xor_out[73][15][19] + xor_out[74][15][19];
assign sum_out[15][15][19] = xor_out[75][15][19] + xor_out[76][15][19] + xor_out[77][15][19] + xor_out[78][15][19] + xor_out[79][15][19];
assign sum_out[16][15][19] = xor_out[80][15][19] + xor_out[81][15][19] + xor_out[82][15][19] + xor_out[83][15][19] + xor_out[84][15][19];
assign sum_out[17][15][19] = xor_out[85][15][19] + xor_out[86][15][19] + xor_out[87][15][19] + xor_out[88][15][19] + xor_out[89][15][19];
assign sum_out[18][15][19] = xor_out[90][15][19] + xor_out[91][15][19] + xor_out[92][15][19] + xor_out[93][15][19] + xor_out[94][15][19];
assign sum_out[19][15][19] = xor_out[95][15][19] + xor_out[96][15][19] + xor_out[97][15][19] + xor_out[98][15][19] + xor_out[99][15][19];

assign sum_out[0][15][20] = xor_out[0][15][20] + xor_out[1][15][20] + xor_out[2][15][20] + xor_out[3][15][20] + xor_out[4][15][20];
assign sum_out[1][15][20] = xor_out[5][15][20] + xor_out[6][15][20] + xor_out[7][15][20] + xor_out[8][15][20] + xor_out[9][15][20];
assign sum_out[2][15][20] = xor_out[10][15][20] + xor_out[11][15][20] + xor_out[12][15][20] + xor_out[13][15][20] + xor_out[14][15][20];
assign sum_out[3][15][20] = xor_out[15][15][20] + xor_out[16][15][20] + xor_out[17][15][20] + xor_out[18][15][20] + xor_out[19][15][20];
assign sum_out[4][15][20] = xor_out[20][15][20] + xor_out[21][15][20] + xor_out[22][15][20] + xor_out[23][15][20] + xor_out[24][15][20];
assign sum_out[5][15][20] = xor_out[25][15][20] + xor_out[26][15][20] + xor_out[27][15][20] + xor_out[28][15][20] + xor_out[29][15][20];
assign sum_out[6][15][20] = xor_out[30][15][20] + xor_out[31][15][20] + xor_out[32][15][20] + xor_out[33][15][20] + xor_out[34][15][20];
assign sum_out[7][15][20] = xor_out[35][15][20] + xor_out[36][15][20] + xor_out[37][15][20] + xor_out[38][15][20] + xor_out[39][15][20];
assign sum_out[8][15][20] = xor_out[40][15][20] + xor_out[41][15][20] + xor_out[42][15][20] + xor_out[43][15][20] + xor_out[44][15][20];
assign sum_out[9][15][20] = xor_out[45][15][20] + xor_out[46][15][20] + xor_out[47][15][20] + xor_out[48][15][20] + xor_out[49][15][20];
assign sum_out[10][15][20] = xor_out[50][15][20] + xor_out[51][15][20] + xor_out[52][15][20] + xor_out[53][15][20] + xor_out[54][15][20];
assign sum_out[11][15][20] = xor_out[55][15][20] + xor_out[56][15][20] + xor_out[57][15][20] + xor_out[58][15][20] + xor_out[59][15][20];
assign sum_out[12][15][20] = xor_out[60][15][20] + xor_out[61][15][20] + xor_out[62][15][20] + xor_out[63][15][20] + xor_out[64][15][20];
assign sum_out[13][15][20] = xor_out[65][15][20] + xor_out[66][15][20] + xor_out[67][15][20] + xor_out[68][15][20] + xor_out[69][15][20];
assign sum_out[14][15][20] = xor_out[70][15][20] + xor_out[71][15][20] + xor_out[72][15][20] + xor_out[73][15][20] + xor_out[74][15][20];
assign sum_out[15][15][20] = xor_out[75][15][20] + xor_out[76][15][20] + xor_out[77][15][20] + xor_out[78][15][20] + xor_out[79][15][20];
assign sum_out[16][15][20] = xor_out[80][15][20] + xor_out[81][15][20] + xor_out[82][15][20] + xor_out[83][15][20] + xor_out[84][15][20];
assign sum_out[17][15][20] = xor_out[85][15][20] + xor_out[86][15][20] + xor_out[87][15][20] + xor_out[88][15][20] + xor_out[89][15][20];
assign sum_out[18][15][20] = xor_out[90][15][20] + xor_out[91][15][20] + xor_out[92][15][20] + xor_out[93][15][20] + xor_out[94][15][20];
assign sum_out[19][15][20] = xor_out[95][15][20] + xor_out[96][15][20] + xor_out[97][15][20] + xor_out[98][15][20] + xor_out[99][15][20];

assign sum_out[0][15][21] = xor_out[0][15][21] + xor_out[1][15][21] + xor_out[2][15][21] + xor_out[3][15][21] + xor_out[4][15][21];
assign sum_out[1][15][21] = xor_out[5][15][21] + xor_out[6][15][21] + xor_out[7][15][21] + xor_out[8][15][21] + xor_out[9][15][21];
assign sum_out[2][15][21] = xor_out[10][15][21] + xor_out[11][15][21] + xor_out[12][15][21] + xor_out[13][15][21] + xor_out[14][15][21];
assign sum_out[3][15][21] = xor_out[15][15][21] + xor_out[16][15][21] + xor_out[17][15][21] + xor_out[18][15][21] + xor_out[19][15][21];
assign sum_out[4][15][21] = xor_out[20][15][21] + xor_out[21][15][21] + xor_out[22][15][21] + xor_out[23][15][21] + xor_out[24][15][21];
assign sum_out[5][15][21] = xor_out[25][15][21] + xor_out[26][15][21] + xor_out[27][15][21] + xor_out[28][15][21] + xor_out[29][15][21];
assign sum_out[6][15][21] = xor_out[30][15][21] + xor_out[31][15][21] + xor_out[32][15][21] + xor_out[33][15][21] + xor_out[34][15][21];
assign sum_out[7][15][21] = xor_out[35][15][21] + xor_out[36][15][21] + xor_out[37][15][21] + xor_out[38][15][21] + xor_out[39][15][21];
assign sum_out[8][15][21] = xor_out[40][15][21] + xor_out[41][15][21] + xor_out[42][15][21] + xor_out[43][15][21] + xor_out[44][15][21];
assign sum_out[9][15][21] = xor_out[45][15][21] + xor_out[46][15][21] + xor_out[47][15][21] + xor_out[48][15][21] + xor_out[49][15][21];
assign sum_out[10][15][21] = xor_out[50][15][21] + xor_out[51][15][21] + xor_out[52][15][21] + xor_out[53][15][21] + xor_out[54][15][21];
assign sum_out[11][15][21] = xor_out[55][15][21] + xor_out[56][15][21] + xor_out[57][15][21] + xor_out[58][15][21] + xor_out[59][15][21];
assign sum_out[12][15][21] = xor_out[60][15][21] + xor_out[61][15][21] + xor_out[62][15][21] + xor_out[63][15][21] + xor_out[64][15][21];
assign sum_out[13][15][21] = xor_out[65][15][21] + xor_out[66][15][21] + xor_out[67][15][21] + xor_out[68][15][21] + xor_out[69][15][21];
assign sum_out[14][15][21] = xor_out[70][15][21] + xor_out[71][15][21] + xor_out[72][15][21] + xor_out[73][15][21] + xor_out[74][15][21];
assign sum_out[15][15][21] = xor_out[75][15][21] + xor_out[76][15][21] + xor_out[77][15][21] + xor_out[78][15][21] + xor_out[79][15][21];
assign sum_out[16][15][21] = xor_out[80][15][21] + xor_out[81][15][21] + xor_out[82][15][21] + xor_out[83][15][21] + xor_out[84][15][21];
assign sum_out[17][15][21] = xor_out[85][15][21] + xor_out[86][15][21] + xor_out[87][15][21] + xor_out[88][15][21] + xor_out[89][15][21];
assign sum_out[18][15][21] = xor_out[90][15][21] + xor_out[91][15][21] + xor_out[92][15][21] + xor_out[93][15][21] + xor_out[94][15][21];
assign sum_out[19][15][21] = xor_out[95][15][21] + xor_out[96][15][21] + xor_out[97][15][21] + xor_out[98][15][21] + xor_out[99][15][21];

assign sum_out[0][15][22] = xor_out[0][15][22] + xor_out[1][15][22] + xor_out[2][15][22] + xor_out[3][15][22] + xor_out[4][15][22];
assign sum_out[1][15][22] = xor_out[5][15][22] + xor_out[6][15][22] + xor_out[7][15][22] + xor_out[8][15][22] + xor_out[9][15][22];
assign sum_out[2][15][22] = xor_out[10][15][22] + xor_out[11][15][22] + xor_out[12][15][22] + xor_out[13][15][22] + xor_out[14][15][22];
assign sum_out[3][15][22] = xor_out[15][15][22] + xor_out[16][15][22] + xor_out[17][15][22] + xor_out[18][15][22] + xor_out[19][15][22];
assign sum_out[4][15][22] = xor_out[20][15][22] + xor_out[21][15][22] + xor_out[22][15][22] + xor_out[23][15][22] + xor_out[24][15][22];
assign sum_out[5][15][22] = xor_out[25][15][22] + xor_out[26][15][22] + xor_out[27][15][22] + xor_out[28][15][22] + xor_out[29][15][22];
assign sum_out[6][15][22] = xor_out[30][15][22] + xor_out[31][15][22] + xor_out[32][15][22] + xor_out[33][15][22] + xor_out[34][15][22];
assign sum_out[7][15][22] = xor_out[35][15][22] + xor_out[36][15][22] + xor_out[37][15][22] + xor_out[38][15][22] + xor_out[39][15][22];
assign sum_out[8][15][22] = xor_out[40][15][22] + xor_out[41][15][22] + xor_out[42][15][22] + xor_out[43][15][22] + xor_out[44][15][22];
assign sum_out[9][15][22] = xor_out[45][15][22] + xor_out[46][15][22] + xor_out[47][15][22] + xor_out[48][15][22] + xor_out[49][15][22];
assign sum_out[10][15][22] = xor_out[50][15][22] + xor_out[51][15][22] + xor_out[52][15][22] + xor_out[53][15][22] + xor_out[54][15][22];
assign sum_out[11][15][22] = xor_out[55][15][22] + xor_out[56][15][22] + xor_out[57][15][22] + xor_out[58][15][22] + xor_out[59][15][22];
assign sum_out[12][15][22] = xor_out[60][15][22] + xor_out[61][15][22] + xor_out[62][15][22] + xor_out[63][15][22] + xor_out[64][15][22];
assign sum_out[13][15][22] = xor_out[65][15][22] + xor_out[66][15][22] + xor_out[67][15][22] + xor_out[68][15][22] + xor_out[69][15][22];
assign sum_out[14][15][22] = xor_out[70][15][22] + xor_out[71][15][22] + xor_out[72][15][22] + xor_out[73][15][22] + xor_out[74][15][22];
assign sum_out[15][15][22] = xor_out[75][15][22] + xor_out[76][15][22] + xor_out[77][15][22] + xor_out[78][15][22] + xor_out[79][15][22];
assign sum_out[16][15][22] = xor_out[80][15][22] + xor_out[81][15][22] + xor_out[82][15][22] + xor_out[83][15][22] + xor_out[84][15][22];
assign sum_out[17][15][22] = xor_out[85][15][22] + xor_out[86][15][22] + xor_out[87][15][22] + xor_out[88][15][22] + xor_out[89][15][22];
assign sum_out[18][15][22] = xor_out[90][15][22] + xor_out[91][15][22] + xor_out[92][15][22] + xor_out[93][15][22] + xor_out[94][15][22];
assign sum_out[19][15][22] = xor_out[95][15][22] + xor_out[96][15][22] + xor_out[97][15][22] + xor_out[98][15][22] + xor_out[99][15][22];

assign sum_out[0][15][23] = xor_out[0][15][23] + xor_out[1][15][23] + xor_out[2][15][23] + xor_out[3][15][23] + xor_out[4][15][23];
assign sum_out[1][15][23] = xor_out[5][15][23] + xor_out[6][15][23] + xor_out[7][15][23] + xor_out[8][15][23] + xor_out[9][15][23];
assign sum_out[2][15][23] = xor_out[10][15][23] + xor_out[11][15][23] + xor_out[12][15][23] + xor_out[13][15][23] + xor_out[14][15][23];
assign sum_out[3][15][23] = xor_out[15][15][23] + xor_out[16][15][23] + xor_out[17][15][23] + xor_out[18][15][23] + xor_out[19][15][23];
assign sum_out[4][15][23] = xor_out[20][15][23] + xor_out[21][15][23] + xor_out[22][15][23] + xor_out[23][15][23] + xor_out[24][15][23];
assign sum_out[5][15][23] = xor_out[25][15][23] + xor_out[26][15][23] + xor_out[27][15][23] + xor_out[28][15][23] + xor_out[29][15][23];
assign sum_out[6][15][23] = xor_out[30][15][23] + xor_out[31][15][23] + xor_out[32][15][23] + xor_out[33][15][23] + xor_out[34][15][23];
assign sum_out[7][15][23] = xor_out[35][15][23] + xor_out[36][15][23] + xor_out[37][15][23] + xor_out[38][15][23] + xor_out[39][15][23];
assign sum_out[8][15][23] = xor_out[40][15][23] + xor_out[41][15][23] + xor_out[42][15][23] + xor_out[43][15][23] + xor_out[44][15][23];
assign sum_out[9][15][23] = xor_out[45][15][23] + xor_out[46][15][23] + xor_out[47][15][23] + xor_out[48][15][23] + xor_out[49][15][23];
assign sum_out[10][15][23] = xor_out[50][15][23] + xor_out[51][15][23] + xor_out[52][15][23] + xor_out[53][15][23] + xor_out[54][15][23];
assign sum_out[11][15][23] = xor_out[55][15][23] + xor_out[56][15][23] + xor_out[57][15][23] + xor_out[58][15][23] + xor_out[59][15][23];
assign sum_out[12][15][23] = xor_out[60][15][23] + xor_out[61][15][23] + xor_out[62][15][23] + xor_out[63][15][23] + xor_out[64][15][23];
assign sum_out[13][15][23] = xor_out[65][15][23] + xor_out[66][15][23] + xor_out[67][15][23] + xor_out[68][15][23] + xor_out[69][15][23];
assign sum_out[14][15][23] = xor_out[70][15][23] + xor_out[71][15][23] + xor_out[72][15][23] + xor_out[73][15][23] + xor_out[74][15][23];
assign sum_out[15][15][23] = xor_out[75][15][23] + xor_out[76][15][23] + xor_out[77][15][23] + xor_out[78][15][23] + xor_out[79][15][23];
assign sum_out[16][15][23] = xor_out[80][15][23] + xor_out[81][15][23] + xor_out[82][15][23] + xor_out[83][15][23] + xor_out[84][15][23];
assign sum_out[17][15][23] = xor_out[85][15][23] + xor_out[86][15][23] + xor_out[87][15][23] + xor_out[88][15][23] + xor_out[89][15][23];
assign sum_out[18][15][23] = xor_out[90][15][23] + xor_out[91][15][23] + xor_out[92][15][23] + xor_out[93][15][23] + xor_out[94][15][23];
assign sum_out[19][15][23] = xor_out[95][15][23] + xor_out[96][15][23] + xor_out[97][15][23] + xor_out[98][15][23] + xor_out[99][15][23];

assign sum_out[0][16][0] = xor_out[0][16][0] + xor_out[1][16][0] + xor_out[2][16][0] + xor_out[3][16][0] + xor_out[4][16][0];
assign sum_out[1][16][0] = xor_out[5][16][0] + xor_out[6][16][0] + xor_out[7][16][0] + xor_out[8][16][0] + xor_out[9][16][0];
assign sum_out[2][16][0] = xor_out[10][16][0] + xor_out[11][16][0] + xor_out[12][16][0] + xor_out[13][16][0] + xor_out[14][16][0];
assign sum_out[3][16][0] = xor_out[15][16][0] + xor_out[16][16][0] + xor_out[17][16][0] + xor_out[18][16][0] + xor_out[19][16][0];
assign sum_out[4][16][0] = xor_out[20][16][0] + xor_out[21][16][0] + xor_out[22][16][0] + xor_out[23][16][0] + xor_out[24][16][0];
assign sum_out[5][16][0] = xor_out[25][16][0] + xor_out[26][16][0] + xor_out[27][16][0] + xor_out[28][16][0] + xor_out[29][16][0];
assign sum_out[6][16][0] = xor_out[30][16][0] + xor_out[31][16][0] + xor_out[32][16][0] + xor_out[33][16][0] + xor_out[34][16][0];
assign sum_out[7][16][0] = xor_out[35][16][0] + xor_out[36][16][0] + xor_out[37][16][0] + xor_out[38][16][0] + xor_out[39][16][0];
assign sum_out[8][16][0] = xor_out[40][16][0] + xor_out[41][16][0] + xor_out[42][16][0] + xor_out[43][16][0] + xor_out[44][16][0];
assign sum_out[9][16][0] = xor_out[45][16][0] + xor_out[46][16][0] + xor_out[47][16][0] + xor_out[48][16][0] + xor_out[49][16][0];
assign sum_out[10][16][0] = xor_out[50][16][0] + xor_out[51][16][0] + xor_out[52][16][0] + xor_out[53][16][0] + xor_out[54][16][0];
assign sum_out[11][16][0] = xor_out[55][16][0] + xor_out[56][16][0] + xor_out[57][16][0] + xor_out[58][16][0] + xor_out[59][16][0];
assign sum_out[12][16][0] = xor_out[60][16][0] + xor_out[61][16][0] + xor_out[62][16][0] + xor_out[63][16][0] + xor_out[64][16][0];
assign sum_out[13][16][0] = xor_out[65][16][0] + xor_out[66][16][0] + xor_out[67][16][0] + xor_out[68][16][0] + xor_out[69][16][0];
assign sum_out[14][16][0] = xor_out[70][16][0] + xor_out[71][16][0] + xor_out[72][16][0] + xor_out[73][16][0] + xor_out[74][16][0];
assign sum_out[15][16][0] = xor_out[75][16][0] + xor_out[76][16][0] + xor_out[77][16][0] + xor_out[78][16][0] + xor_out[79][16][0];
assign sum_out[16][16][0] = xor_out[80][16][0] + xor_out[81][16][0] + xor_out[82][16][0] + xor_out[83][16][0] + xor_out[84][16][0];
assign sum_out[17][16][0] = xor_out[85][16][0] + xor_out[86][16][0] + xor_out[87][16][0] + xor_out[88][16][0] + xor_out[89][16][0];
assign sum_out[18][16][0] = xor_out[90][16][0] + xor_out[91][16][0] + xor_out[92][16][0] + xor_out[93][16][0] + xor_out[94][16][0];
assign sum_out[19][16][0] = xor_out[95][16][0] + xor_out[96][16][0] + xor_out[97][16][0] + xor_out[98][16][0] + xor_out[99][16][0];

assign sum_out[0][16][1] = xor_out[0][16][1] + xor_out[1][16][1] + xor_out[2][16][1] + xor_out[3][16][1] + xor_out[4][16][1];
assign sum_out[1][16][1] = xor_out[5][16][1] + xor_out[6][16][1] + xor_out[7][16][1] + xor_out[8][16][1] + xor_out[9][16][1];
assign sum_out[2][16][1] = xor_out[10][16][1] + xor_out[11][16][1] + xor_out[12][16][1] + xor_out[13][16][1] + xor_out[14][16][1];
assign sum_out[3][16][1] = xor_out[15][16][1] + xor_out[16][16][1] + xor_out[17][16][1] + xor_out[18][16][1] + xor_out[19][16][1];
assign sum_out[4][16][1] = xor_out[20][16][1] + xor_out[21][16][1] + xor_out[22][16][1] + xor_out[23][16][1] + xor_out[24][16][1];
assign sum_out[5][16][1] = xor_out[25][16][1] + xor_out[26][16][1] + xor_out[27][16][1] + xor_out[28][16][1] + xor_out[29][16][1];
assign sum_out[6][16][1] = xor_out[30][16][1] + xor_out[31][16][1] + xor_out[32][16][1] + xor_out[33][16][1] + xor_out[34][16][1];
assign sum_out[7][16][1] = xor_out[35][16][1] + xor_out[36][16][1] + xor_out[37][16][1] + xor_out[38][16][1] + xor_out[39][16][1];
assign sum_out[8][16][1] = xor_out[40][16][1] + xor_out[41][16][1] + xor_out[42][16][1] + xor_out[43][16][1] + xor_out[44][16][1];
assign sum_out[9][16][1] = xor_out[45][16][1] + xor_out[46][16][1] + xor_out[47][16][1] + xor_out[48][16][1] + xor_out[49][16][1];
assign sum_out[10][16][1] = xor_out[50][16][1] + xor_out[51][16][1] + xor_out[52][16][1] + xor_out[53][16][1] + xor_out[54][16][1];
assign sum_out[11][16][1] = xor_out[55][16][1] + xor_out[56][16][1] + xor_out[57][16][1] + xor_out[58][16][1] + xor_out[59][16][1];
assign sum_out[12][16][1] = xor_out[60][16][1] + xor_out[61][16][1] + xor_out[62][16][1] + xor_out[63][16][1] + xor_out[64][16][1];
assign sum_out[13][16][1] = xor_out[65][16][1] + xor_out[66][16][1] + xor_out[67][16][1] + xor_out[68][16][1] + xor_out[69][16][1];
assign sum_out[14][16][1] = xor_out[70][16][1] + xor_out[71][16][1] + xor_out[72][16][1] + xor_out[73][16][1] + xor_out[74][16][1];
assign sum_out[15][16][1] = xor_out[75][16][1] + xor_out[76][16][1] + xor_out[77][16][1] + xor_out[78][16][1] + xor_out[79][16][1];
assign sum_out[16][16][1] = xor_out[80][16][1] + xor_out[81][16][1] + xor_out[82][16][1] + xor_out[83][16][1] + xor_out[84][16][1];
assign sum_out[17][16][1] = xor_out[85][16][1] + xor_out[86][16][1] + xor_out[87][16][1] + xor_out[88][16][1] + xor_out[89][16][1];
assign sum_out[18][16][1] = xor_out[90][16][1] + xor_out[91][16][1] + xor_out[92][16][1] + xor_out[93][16][1] + xor_out[94][16][1];
assign sum_out[19][16][1] = xor_out[95][16][1] + xor_out[96][16][1] + xor_out[97][16][1] + xor_out[98][16][1] + xor_out[99][16][1];

assign sum_out[0][16][2] = xor_out[0][16][2] + xor_out[1][16][2] + xor_out[2][16][2] + xor_out[3][16][2] + xor_out[4][16][2];
assign sum_out[1][16][2] = xor_out[5][16][2] + xor_out[6][16][2] + xor_out[7][16][2] + xor_out[8][16][2] + xor_out[9][16][2];
assign sum_out[2][16][2] = xor_out[10][16][2] + xor_out[11][16][2] + xor_out[12][16][2] + xor_out[13][16][2] + xor_out[14][16][2];
assign sum_out[3][16][2] = xor_out[15][16][2] + xor_out[16][16][2] + xor_out[17][16][2] + xor_out[18][16][2] + xor_out[19][16][2];
assign sum_out[4][16][2] = xor_out[20][16][2] + xor_out[21][16][2] + xor_out[22][16][2] + xor_out[23][16][2] + xor_out[24][16][2];
assign sum_out[5][16][2] = xor_out[25][16][2] + xor_out[26][16][2] + xor_out[27][16][2] + xor_out[28][16][2] + xor_out[29][16][2];
assign sum_out[6][16][2] = xor_out[30][16][2] + xor_out[31][16][2] + xor_out[32][16][2] + xor_out[33][16][2] + xor_out[34][16][2];
assign sum_out[7][16][2] = xor_out[35][16][2] + xor_out[36][16][2] + xor_out[37][16][2] + xor_out[38][16][2] + xor_out[39][16][2];
assign sum_out[8][16][2] = xor_out[40][16][2] + xor_out[41][16][2] + xor_out[42][16][2] + xor_out[43][16][2] + xor_out[44][16][2];
assign sum_out[9][16][2] = xor_out[45][16][2] + xor_out[46][16][2] + xor_out[47][16][2] + xor_out[48][16][2] + xor_out[49][16][2];
assign sum_out[10][16][2] = xor_out[50][16][2] + xor_out[51][16][2] + xor_out[52][16][2] + xor_out[53][16][2] + xor_out[54][16][2];
assign sum_out[11][16][2] = xor_out[55][16][2] + xor_out[56][16][2] + xor_out[57][16][2] + xor_out[58][16][2] + xor_out[59][16][2];
assign sum_out[12][16][2] = xor_out[60][16][2] + xor_out[61][16][2] + xor_out[62][16][2] + xor_out[63][16][2] + xor_out[64][16][2];
assign sum_out[13][16][2] = xor_out[65][16][2] + xor_out[66][16][2] + xor_out[67][16][2] + xor_out[68][16][2] + xor_out[69][16][2];
assign sum_out[14][16][2] = xor_out[70][16][2] + xor_out[71][16][2] + xor_out[72][16][2] + xor_out[73][16][2] + xor_out[74][16][2];
assign sum_out[15][16][2] = xor_out[75][16][2] + xor_out[76][16][2] + xor_out[77][16][2] + xor_out[78][16][2] + xor_out[79][16][2];
assign sum_out[16][16][2] = xor_out[80][16][2] + xor_out[81][16][2] + xor_out[82][16][2] + xor_out[83][16][2] + xor_out[84][16][2];
assign sum_out[17][16][2] = xor_out[85][16][2] + xor_out[86][16][2] + xor_out[87][16][2] + xor_out[88][16][2] + xor_out[89][16][2];
assign sum_out[18][16][2] = xor_out[90][16][2] + xor_out[91][16][2] + xor_out[92][16][2] + xor_out[93][16][2] + xor_out[94][16][2];
assign sum_out[19][16][2] = xor_out[95][16][2] + xor_out[96][16][2] + xor_out[97][16][2] + xor_out[98][16][2] + xor_out[99][16][2];

assign sum_out[0][16][3] = xor_out[0][16][3] + xor_out[1][16][3] + xor_out[2][16][3] + xor_out[3][16][3] + xor_out[4][16][3];
assign sum_out[1][16][3] = xor_out[5][16][3] + xor_out[6][16][3] + xor_out[7][16][3] + xor_out[8][16][3] + xor_out[9][16][3];
assign sum_out[2][16][3] = xor_out[10][16][3] + xor_out[11][16][3] + xor_out[12][16][3] + xor_out[13][16][3] + xor_out[14][16][3];
assign sum_out[3][16][3] = xor_out[15][16][3] + xor_out[16][16][3] + xor_out[17][16][3] + xor_out[18][16][3] + xor_out[19][16][3];
assign sum_out[4][16][3] = xor_out[20][16][3] + xor_out[21][16][3] + xor_out[22][16][3] + xor_out[23][16][3] + xor_out[24][16][3];
assign sum_out[5][16][3] = xor_out[25][16][3] + xor_out[26][16][3] + xor_out[27][16][3] + xor_out[28][16][3] + xor_out[29][16][3];
assign sum_out[6][16][3] = xor_out[30][16][3] + xor_out[31][16][3] + xor_out[32][16][3] + xor_out[33][16][3] + xor_out[34][16][3];
assign sum_out[7][16][3] = xor_out[35][16][3] + xor_out[36][16][3] + xor_out[37][16][3] + xor_out[38][16][3] + xor_out[39][16][3];
assign sum_out[8][16][3] = xor_out[40][16][3] + xor_out[41][16][3] + xor_out[42][16][3] + xor_out[43][16][3] + xor_out[44][16][3];
assign sum_out[9][16][3] = xor_out[45][16][3] + xor_out[46][16][3] + xor_out[47][16][3] + xor_out[48][16][3] + xor_out[49][16][3];
assign sum_out[10][16][3] = xor_out[50][16][3] + xor_out[51][16][3] + xor_out[52][16][3] + xor_out[53][16][3] + xor_out[54][16][3];
assign sum_out[11][16][3] = xor_out[55][16][3] + xor_out[56][16][3] + xor_out[57][16][3] + xor_out[58][16][3] + xor_out[59][16][3];
assign sum_out[12][16][3] = xor_out[60][16][3] + xor_out[61][16][3] + xor_out[62][16][3] + xor_out[63][16][3] + xor_out[64][16][3];
assign sum_out[13][16][3] = xor_out[65][16][3] + xor_out[66][16][3] + xor_out[67][16][3] + xor_out[68][16][3] + xor_out[69][16][3];
assign sum_out[14][16][3] = xor_out[70][16][3] + xor_out[71][16][3] + xor_out[72][16][3] + xor_out[73][16][3] + xor_out[74][16][3];
assign sum_out[15][16][3] = xor_out[75][16][3] + xor_out[76][16][3] + xor_out[77][16][3] + xor_out[78][16][3] + xor_out[79][16][3];
assign sum_out[16][16][3] = xor_out[80][16][3] + xor_out[81][16][3] + xor_out[82][16][3] + xor_out[83][16][3] + xor_out[84][16][3];
assign sum_out[17][16][3] = xor_out[85][16][3] + xor_out[86][16][3] + xor_out[87][16][3] + xor_out[88][16][3] + xor_out[89][16][3];
assign sum_out[18][16][3] = xor_out[90][16][3] + xor_out[91][16][3] + xor_out[92][16][3] + xor_out[93][16][3] + xor_out[94][16][3];
assign sum_out[19][16][3] = xor_out[95][16][3] + xor_out[96][16][3] + xor_out[97][16][3] + xor_out[98][16][3] + xor_out[99][16][3];

assign sum_out[0][16][4] = xor_out[0][16][4] + xor_out[1][16][4] + xor_out[2][16][4] + xor_out[3][16][4] + xor_out[4][16][4];
assign sum_out[1][16][4] = xor_out[5][16][4] + xor_out[6][16][4] + xor_out[7][16][4] + xor_out[8][16][4] + xor_out[9][16][4];
assign sum_out[2][16][4] = xor_out[10][16][4] + xor_out[11][16][4] + xor_out[12][16][4] + xor_out[13][16][4] + xor_out[14][16][4];
assign sum_out[3][16][4] = xor_out[15][16][4] + xor_out[16][16][4] + xor_out[17][16][4] + xor_out[18][16][4] + xor_out[19][16][4];
assign sum_out[4][16][4] = xor_out[20][16][4] + xor_out[21][16][4] + xor_out[22][16][4] + xor_out[23][16][4] + xor_out[24][16][4];
assign sum_out[5][16][4] = xor_out[25][16][4] + xor_out[26][16][4] + xor_out[27][16][4] + xor_out[28][16][4] + xor_out[29][16][4];
assign sum_out[6][16][4] = xor_out[30][16][4] + xor_out[31][16][4] + xor_out[32][16][4] + xor_out[33][16][4] + xor_out[34][16][4];
assign sum_out[7][16][4] = xor_out[35][16][4] + xor_out[36][16][4] + xor_out[37][16][4] + xor_out[38][16][4] + xor_out[39][16][4];
assign sum_out[8][16][4] = xor_out[40][16][4] + xor_out[41][16][4] + xor_out[42][16][4] + xor_out[43][16][4] + xor_out[44][16][4];
assign sum_out[9][16][4] = xor_out[45][16][4] + xor_out[46][16][4] + xor_out[47][16][4] + xor_out[48][16][4] + xor_out[49][16][4];
assign sum_out[10][16][4] = xor_out[50][16][4] + xor_out[51][16][4] + xor_out[52][16][4] + xor_out[53][16][4] + xor_out[54][16][4];
assign sum_out[11][16][4] = xor_out[55][16][4] + xor_out[56][16][4] + xor_out[57][16][4] + xor_out[58][16][4] + xor_out[59][16][4];
assign sum_out[12][16][4] = xor_out[60][16][4] + xor_out[61][16][4] + xor_out[62][16][4] + xor_out[63][16][4] + xor_out[64][16][4];
assign sum_out[13][16][4] = xor_out[65][16][4] + xor_out[66][16][4] + xor_out[67][16][4] + xor_out[68][16][4] + xor_out[69][16][4];
assign sum_out[14][16][4] = xor_out[70][16][4] + xor_out[71][16][4] + xor_out[72][16][4] + xor_out[73][16][4] + xor_out[74][16][4];
assign sum_out[15][16][4] = xor_out[75][16][4] + xor_out[76][16][4] + xor_out[77][16][4] + xor_out[78][16][4] + xor_out[79][16][4];
assign sum_out[16][16][4] = xor_out[80][16][4] + xor_out[81][16][4] + xor_out[82][16][4] + xor_out[83][16][4] + xor_out[84][16][4];
assign sum_out[17][16][4] = xor_out[85][16][4] + xor_out[86][16][4] + xor_out[87][16][4] + xor_out[88][16][4] + xor_out[89][16][4];
assign sum_out[18][16][4] = xor_out[90][16][4] + xor_out[91][16][4] + xor_out[92][16][4] + xor_out[93][16][4] + xor_out[94][16][4];
assign sum_out[19][16][4] = xor_out[95][16][4] + xor_out[96][16][4] + xor_out[97][16][4] + xor_out[98][16][4] + xor_out[99][16][4];

assign sum_out[0][16][5] = xor_out[0][16][5] + xor_out[1][16][5] + xor_out[2][16][5] + xor_out[3][16][5] + xor_out[4][16][5];
assign sum_out[1][16][5] = xor_out[5][16][5] + xor_out[6][16][5] + xor_out[7][16][5] + xor_out[8][16][5] + xor_out[9][16][5];
assign sum_out[2][16][5] = xor_out[10][16][5] + xor_out[11][16][5] + xor_out[12][16][5] + xor_out[13][16][5] + xor_out[14][16][5];
assign sum_out[3][16][5] = xor_out[15][16][5] + xor_out[16][16][5] + xor_out[17][16][5] + xor_out[18][16][5] + xor_out[19][16][5];
assign sum_out[4][16][5] = xor_out[20][16][5] + xor_out[21][16][5] + xor_out[22][16][5] + xor_out[23][16][5] + xor_out[24][16][5];
assign sum_out[5][16][5] = xor_out[25][16][5] + xor_out[26][16][5] + xor_out[27][16][5] + xor_out[28][16][5] + xor_out[29][16][5];
assign sum_out[6][16][5] = xor_out[30][16][5] + xor_out[31][16][5] + xor_out[32][16][5] + xor_out[33][16][5] + xor_out[34][16][5];
assign sum_out[7][16][5] = xor_out[35][16][5] + xor_out[36][16][5] + xor_out[37][16][5] + xor_out[38][16][5] + xor_out[39][16][5];
assign sum_out[8][16][5] = xor_out[40][16][5] + xor_out[41][16][5] + xor_out[42][16][5] + xor_out[43][16][5] + xor_out[44][16][5];
assign sum_out[9][16][5] = xor_out[45][16][5] + xor_out[46][16][5] + xor_out[47][16][5] + xor_out[48][16][5] + xor_out[49][16][5];
assign sum_out[10][16][5] = xor_out[50][16][5] + xor_out[51][16][5] + xor_out[52][16][5] + xor_out[53][16][5] + xor_out[54][16][5];
assign sum_out[11][16][5] = xor_out[55][16][5] + xor_out[56][16][5] + xor_out[57][16][5] + xor_out[58][16][5] + xor_out[59][16][5];
assign sum_out[12][16][5] = xor_out[60][16][5] + xor_out[61][16][5] + xor_out[62][16][5] + xor_out[63][16][5] + xor_out[64][16][5];
assign sum_out[13][16][5] = xor_out[65][16][5] + xor_out[66][16][5] + xor_out[67][16][5] + xor_out[68][16][5] + xor_out[69][16][5];
assign sum_out[14][16][5] = xor_out[70][16][5] + xor_out[71][16][5] + xor_out[72][16][5] + xor_out[73][16][5] + xor_out[74][16][5];
assign sum_out[15][16][5] = xor_out[75][16][5] + xor_out[76][16][5] + xor_out[77][16][5] + xor_out[78][16][5] + xor_out[79][16][5];
assign sum_out[16][16][5] = xor_out[80][16][5] + xor_out[81][16][5] + xor_out[82][16][5] + xor_out[83][16][5] + xor_out[84][16][5];
assign sum_out[17][16][5] = xor_out[85][16][5] + xor_out[86][16][5] + xor_out[87][16][5] + xor_out[88][16][5] + xor_out[89][16][5];
assign sum_out[18][16][5] = xor_out[90][16][5] + xor_out[91][16][5] + xor_out[92][16][5] + xor_out[93][16][5] + xor_out[94][16][5];
assign sum_out[19][16][5] = xor_out[95][16][5] + xor_out[96][16][5] + xor_out[97][16][5] + xor_out[98][16][5] + xor_out[99][16][5];

assign sum_out[0][16][6] = xor_out[0][16][6] + xor_out[1][16][6] + xor_out[2][16][6] + xor_out[3][16][6] + xor_out[4][16][6];
assign sum_out[1][16][6] = xor_out[5][16][6] + xor_out[6][16][6] + xor_out[7][16][6] + xor_out[8][16][6] + xor_out[9][16][6];
assign sum_out[2][16][6] = xor_out[10][16][6] + xor_out[11][16][6] + xor_out[12][16][6] + xor_out[13][16][6] + xor_out[14][16][6];
assign sum_out[3][16][6] = xor_out[15][16][6] + xor_out[16][16][6] + xor_out[17][16][6] + xor_out[18][16][6] + xor_out[19][16][6];
assign sum_out[4][16][6] = xor_out[20][16][6] + xor_out[21][16][6] + xor_out[22][16][6] + xor_out[23][16][6] + xor_out[24][16][6];
assign sum_out[5][16][6] = xor_out[25][16][6] + xor_out[26][16][6] + xor_out[27][16][6] + xor_out[28][16][6] + xor_out[29][16][6];
assign sum_out[6][16][6] = xor_out[30][16][6] + xor_out[31][16][6] + xor_out[32][16][6] + xor_out[33][16][6] + xor_out[34][16][6];
assign sum_out[7][16][6] = xor_out[35][16][6] + xor_out[36][16][6] + xor_out[37][16][6] + xor_out[38][16][6] + xor_out[39][16][6];
assign sum_out[8][16][6] = xor_out[40][16][6] + xor_out[41][16][6] + xor_out[42][16][6] + xor_out[43][16][6] + xor_out[44][16][6];
assign sum_out[9][16][6] = xor_out[45][16][6] + xor_out[46][16][6] + xor_out[47][16][6] + xor_out[48][16][6] + xor_out[49][16][6];
assign sum_out[10][16][6] = xor_out[50][16][6] + xor_out[51][16][6] + xor_out[52][16][6] + xor_out[53][16][6] + xor_out[54][16][6];
assign sum_out[11][16][6] = xor_out[55][16][6] + xor_out[56][16][6] + xor_out[57][16][6] + xor_out[58][16][6] + xor_out[59][16][6];
assign sum_out[12][16][6] = xor_out[60][16][6] + xor_out[61][16][6] + xor_out[62][16][6] + xor_out[63][16][6] + xor_out[64][16][6];
assign sum_out[13][16][6] = xor_out[65][16][6] + xor_out[66][16][6] + xor_out[67][16][6] + xor_out[68][16][6] + xor_out[69][16][6];
assign sum_out[14][16][6] = xor_out[70][16][6] + xor_out[71][16][6] + xor_out[72][16][6] + xor_out[73][16][6] + xor_out[74][16][6];
assign sum_out[15][16][6] = xor_out[75][16][6] + xor_out[76][16][6] + xor_out[77][16][6] + xor_out[78][16][6] + xor_out[79][16][6];
assign sum_out[16][16][6] = xor_out[80][16][6] + xor_out[81][16][6] + xor_out[82][16][6] + xor_out[83][16][6] + xor_out[84][16][6];
assign sum_out[17][16][6] = xor_out[85][16][6] + xor_out[86][16][6] + xor_out[87][16][6] + xor_out[88][16][6] + xor_out[89][16][6];
assign sum_out[18][16][6] = xor_out[90][16][6] + xor_out[91][16][6] + xor_out[92][16][6] + xor_out[93][16][6] + xor_out[94][16][6];
assign sum_out[19][16][6] = xor_out[95][16][6] + xor_out[96][16][6] + xor_out[97][16][6] + xor_out[98][16][6] + xor_out[99][16][6];

assign sum_out[0][16][7] = xor_out[0][16][7] + xor_out[1][16][7] + xor_out[2][16][7] + xor_out[3][16][7] + xor_out[4][16][7];
assign sum_out[1][16][7] = xor_out[5][16][7] + xor_out[6][16][7] + xor_out[7][16][7] + xor_out[8][16][7] + xor_out[9][16][7];
assign sum_out[2][16][7] = xor_out[10][16][7] + xor_out[11][16][7] + xor_out[12][16][7] + xor_out[13][16][7] + xor_out[14][16][7];
assign sum_out[3][16][7] = xor_out[15][16][7] + xor_out[16][16][7] + xor_out[17][16][7] + xor_out[18][16][7] + xor_out[19][16][7];
assign sum_out[4][16][7] = xor_out[20][16][7] + xor_out[21][16][7] + xor_out[22][16][7] + xor_out[23][16][7] + xor_out[24][16][7];
assign sum_out[5][16][7] = xor_out[25][16][7] + xor_out[26][16][7] + xor_out[27][16][7] + xor_out[28][16][7] + xor_out[29][16][7];
assign sum_out[6][16][7] = xor_out[30][16][7] + xor_out[31][16][7] + xor_out[32][16][7] + xor_out[33][16][7] + xor_out[34][16][7];
assign sum_out[7][16][7] = xor_out[35][16][7] + xor_out[36][16][7] + xor_out[37][16][7] + xor_out[38][16][7] + xor_out[39][16][7];
assign sum_out[8][16][7] = xor_out[40][16][7] + xor_out[41][16][7] + xor_out[42][16][7] + xor_out[43][16][7] + xor_out[44][16][7];
assign sum_out[9][16][7] = xor_out[45][16][7] + xor_out[46][16][7] + xor_out[47][16][7] + xor_out[48][16][7] + xor_out[49][16][7];
assign sum_out[10][16][7] = xor_out[50][16][7] + xor_out[51][16][7] + xor_out[52][16][7] + xor_out[53][16][7] + xor_out[54][16][7];
assign sum_out[11][16][7] = xor_out[55][16][7] + xor_out[56][16][7] + xor_out[57][16][7] + xor_out[58][16][7] + xor_out[59][16][7];
assign sum_out[12][16][7] = xor_out[60][16][7] + xor_out[61][16][7] + xor_out[62][16][7] + xor_out[63][16][7] + xor_out[64][16][7];
assign sum_out[13][16][7] = xor_out[65][16][7] + xor_out[66][16][7] + xor_out[67][16][7] + xor_out[68][16][7] + xor_out[69][16][7];
assign sum_out[14][16][7] = xor_out[70][16][7] + xor_out[71][16][7] + xor_out[72][16][7] + xor_out[73][16][7] + xor_out[74][16][7];
assign sum_out[15][16][7] = xor_out[75][16][7] + xor_out[76][16][7] + xor_out[77][16][7] + xor_out[78][16][7] + xor_out[79][16][7];
assign sum_out[16][16][7] = xor_out[80][16][7] + xor_out[81][16][7] + xor_out[82][16][7] + xor_out[83][16][7] + xor_out[84][16][7];
assign sum_out[17][16][7] = xor_out[85][16][7] + xor_out[86][16][7] + xor_out[87][16][7] + xor_out[88][16][7] + xor_out[89][16][7];
assign sum_out[18][16][7] = xor_out[90][16][7] + xor_out[91][16][7] + xor_out[92][16][7] + xor_out[93][16][7] + xor_out[94][16][7];
assign sum_out[19][16][7] = xor_out[95][16][7] + xor_out[96][16][7] + xor_out[97][16][7] + xor_out[98][16][7] + xor_out[99][16][7];

assign sum_out[0][16][8] = xor_out[0][16][8] + xor_out[1][16][8] + xor_out[2][16][8] + xor_out[3][16][8] + xor_out[4][16][8];
assign sum_out[1][16][8] = xor_out[5][16][8] + xor_out[6][16][8] + xor_out[7][16][8] + xor_out[8][16][8] + xor_out[9][16][8];
assign sum_out[2][16][8] = xor_out[10][16][8] + xor_out[11][16][8] + xor_out[12][16][8] + xor_out[13][16][8] + xor_out[14][16][8];
assign sum_out[3][16][8] = xor_out[15][16][8] + xor_out[16][16][8] + xor_out[17][16][8] + xor_out[18][16][8] + xor_out[19][16][8];
assign sum_out[4][16][8] = xor_out[20][16][8] + xor_out[21][16][8] + xor_out[22][16][8] + xor_out[23][16][8] + xor_out[24][16][8];
assign sum_out[5][16][8] = xor_out[25][16][8] + xor_out[26][16][8] + xor_out[27][16][8] + xor_out[28][16][8] + xor_out[29][16][8];
assign sum_out[6][16][8] = xor_out[30][16][8] + xor_out[31][16][8] + xor_out[32][16][8] + xor_out[33][16][8] + xor_out[34][16][8];
assign sum_out[7][16][8] = xor_out[35][16][8] + xor_out[36][16][8] + xor_out[37][16][8] + xor_out[38][16][8] + xor_out[39][16][8];
assign sum_out[8][16][8] = xor_out[40][16][8] + xor_out[41][16][8] + xor_out[42][16][8] + xor_out[43][16][8] + xor_out[44][16][8];
assign sum_out[9][16][8] = xor_out[45][16][8] + xor_out[46][16][8] + xor_out[47][16][8] + xor_out[48][16][8] + xor_out[49][16][8];
assign sum_out[10][16][8] = xor_out[50][16][8] + xor_out[51][16][8] + xor_out[52][16][8] + xor_out[53][16][8] + xor_out[54][16][8];
assign sum_out[11][16][8] = xor_out[55][16][8] + xor_out[56][16][8] + xor_out[57][16][8] + xor_out[58][16][8] + xor_out[59][16][8];
assign sum_out[12][16][8] = xor_out[60][16][8] + xor_out[61][16][8] + xor_out[62][16][8] + xor_out[63][16][8] + xor_out[64][16][8];
assign sum_out[13][16][8] = xor_out[65][16][8] + xor_out[66][16][8] + xor_out[67][16][8] + xor_out[68][16][8] + xor_out[69][16][8];
assign sum_out[14][16][8] = xor_out[70][16][8] + xor_out[71][16][8] + xor_out[72][16][8] + xor_out[73][16][8] + xor_out[74][16][8];
assign sum_out[15][16][8] = xor_out[75][16][8] + xor_out[76][16][8] + xor_out[77][16][8] + xor_out[78][16][8] + xor_out[79][16][8];
assign sum_out[16][16][8] = xor_out[80][16][8] + xor_out[81][16][8] + xor_out[82][16][8] + xor_out[83][16][8] + xor_out[84][16][8];
assign sum_out[17][16][8] = xor_out[85][16][8] + xor_out[86][16][8] + xor_out[87][16][8] + xor_out[88][16][8] + xor_out[89][16][8];
assign sum_out[18][16][8] = xor_out[90][16][8] + xor_out[91][16][8] + xor_out[92][16][8] + xor_out[93][16][8] + xor_out[94][16][8];
assign sum_out[19][16][8] = xor_out[95][16][8] + xor_out[96][16][8] + xor_out[97][16][8] + xor_out[98][16][8] + xor_out[99][16][8];

assign sum_out[0][16][9] = xor_out[0][16][9] + xor_out[1][16][9] + xor_out[2][16][9] + xor_out[3][16][9] + xor_out[4][16][9];
assign sum_out[1][16][9] = xor_out[5][16][9] + xor_out[6][16][9] + xor_out[7][16][9] + xor_out[8][16][9] + xor_out[9][16][9];
assign sum_out[2][16][9] = xor_out[10][16][9] + xor_out[11][16][9] + xor_out[12][16][9] + xor_out[13][16][9] + xor_out[14][16][9];
assign sum_out[3][16][9] = xor_out[15][16][9] + xor_out[16][16][9] + xor_out[17][16][9] + xor_out[18][16][9] + xor_out[19][16][9];
assign sum_out[4][16][9] = xor_out[20][16][9] + xor_out[21][16][9] + xor_out[22][16][9] + xor_out[23][16][9] + xor_out[24][16][9];
assign sum_out[5][16][9] = xor_out[25][16][9] + xor_out[26][16][9] + xor_out[27][16][9] + xor_out[28][16][9] + xor_out[29][16][9];
assign sum_out[6][16][9] = xor_out[30][16][9] + xor_out[31][16][9] + xor_out[32][16][9] + xor_out[33][16][9] + xor_out[34][16][9];
assign sum_out[7][16][9] = xor_out[35][16][9] + xor_out[36][16][9] + xor_out[37][16][9] + xor_out[38][16][9] + xor_out[39][16][9];
assign sum_out[8][16][9] = xor_out[40][16][9] + xor_out[41][16][9] + xor_out[42][16][9] + xor_out[43][16][9] + xor_out[44][16][9];
assign sum_out[9][16][9] = xor_out[45][16][9] + xor_out[46][16][9] + xor_out[47][16][9] + xor_out[48][16][9] + xor_out[49][16][9];
assign sum_out[10][16][9] = xor_out[50][16][9] + xor_out[51][16][9] + xor_out[52][16][9] + xor_out[53][16][9] + xor_out[54][16][9];
assign sum_out[11][16][9] = xor_out[55][16][9] + xor_out[56][16][9] + xor_out[57][16][9] + xor_out[58][16][9] + xor_out[59][16][9];
assign sum_out[12][16][9] = xor_out[60][16][9] + xor_out[61][16][9] + xor_out[62][16][9] + xor_out[63][16][9] + xor_out[64][16][9];
assign sum_out[13][16][9] = xor_out[65][16][9] + xor_out[66][16][9] + xor_out[67][16][9] + xor_out[68][16][9] + xor_out[69][16][9];
assign sum_out[14][16][9] = xor_out[70][16][9] + xor_out[71][16][9] + xor_out[72][16][9] + xor_out[73][16][9] + xor_out[74][16][9];
assign sum_out[15][16][9] = xor_out[75][16][9] + xor_out[76][16][9] + xor_out[77][16][9] + xor_out[78][16][9] + xor_out[79][16][9];
assign sum_out[16][16][9] = xor_out[80][16][9] + xor_out[81][16][9] + xor_out[82][16][9] + xor_out[83][16][9] + xor_out[84][16][9];
assign sum_out[17][16][9] = xor_out[85][16][9] + xor_out[86][16][9] + xor_out[87][16][9] + xor_out[88][16][9] + xor_out[89][16][9];
assign sum_out[18][16][9] = xor_out[90][16][9] + xor_out[91][16][9] + xor_out[92][16][9] + xor_out[93][16][9] + xor_out[94][16][9];
assign sum_out[19][16][9] = xor_out[95][16][9] + xor_out[96][16][9] + xor_out[97][16][9] + xor_out[98][16][9] + xor_out[99][16][9];

assign sum_out[0][16][10] = xor_out[0][16][10] + xor_out[1][16][10] + xor_out[2][16][10] + xor_out[3][16][10] + xor_out[4][16][10];
assign sum_out[1][16][10] = xor_out[5][16][10] + xor_out[6][16][10] + xor_out[7][16][10] + xor_out[8][16][10] + xor_out[9][16][10];
assign sum_out[2][16][10] = xor_out[10][16][10] + xor_out[11][16][10] + xor_out[12][16][10] + xor_out[13][16][10] + xor_out[14][16][10];
assign sum_out[3][16][10] = xor_out[15][16][10] + xor_out[16][16][10] + xor_out[17][16][10] + xor_out[18][16][10] + xor_out[19][16][10];
assign sum_out[4][16][10] = xor_out[20][16][10] + xor_out[21][16][10] + xor_out[22][16][10] + xor_out[23][16][10] + xor_out[24][16][10];
assign sum_out[5][16][10] = xor_out[25][16][10] + xor_out[26][16][10] + xor_out[27][16][10] + xor_out[28][16][10] + xor_out[29][16][10];
assign sum_out[6][16][10] = xor_out[30][16][10] + xor_out[31][16][10] + xor_out[32][16][10] + xor_out[33][16][10] + xor_out[34][16][10];
assign sum_out[7][16][10] = xor_out[35][16][10] + xor_out[36][16][10] + xor_out[37][16][10] + xor_out[38][16][10] + xor_out[39][16][10];
assign sum_out[8][16][10] = xor_out[40][16][10] + xor_out[41][16][10] + xor_out[42][16][10] + xor_out[43][16][10] + xor_out[44][16][10];
assign sum_out[9][16][10] = xor_out[45][16][10] + xor_out[46][16][10] + xor_out[47][16][10] + xor_out[48][16][10] + xor_out[49][16][10];
assign sum_out[10][16][10] = xor_out[50][16][10] + xor_out[51][16][10] + xor_out[52][16][10] + xor_out[53][16][10] + xor_out[54][16][10];
assign sum_out[11][16][10] = xor_out[55][16][10] + xor_out[56][16][10] + xor_out[57][16][10] + xor_out[58][16][10] + xor_out[59][16][10];
assign sum_out[12][16][10] = xor_out[60][16][10] + xor_out[61][16][10] + xor_out[62][16][10] + xor_out[63][16][10] + xor_out[64][16][10];
assign sum_out[13][16][10] = xor_out[65][16][10] + xor_out[66][16][10] + xor_out[67][16][10] + xor_out[68][16][10] + xor_out[69][16][10];
assign sum_out[14][16][10] = xor_out[70][16][10] + xor_out[71][16][10] + xor_out[72][16][10] + xor_out[73][16][10] + xor_out[74][16][10];
assign sum_out[15][16][10] = xor_out[75][16][10] + xor_out[76][16][10] + xor_out[77][16][10] + xor_out[78][16][10] + xor_out[79][16][10];
assign sum_out[16][16][10] = xor_out[80][16][10] + xor_out[81][16][10] + xor_out[82][16][10] + xor_out[83][16][10] + xor_out[84][16][10];
assign sum_out[17][16][10] = xor_out[85][16][10] + xor_out[86][16][10] + xor_out[87][16][10] + xor_out[88][16][10] + xor_out[89][16][10];
assign sum_out[18][16][10] = xor_out[90][16][10] + xor_out[91][16][10] + xor_out[92][16][10] + xor_out[93][16][10] + xor_out[94][16][10];
assign sum_out[19][16][10] = xor_out[95][16][10] + xor_out[96][16][10] + xor_out[97][16][10] + xor_out[98][16][10] + xor_out[99][16][10];

assign sum_out[0][16][11] = xor_out[0][16][11] + xor_out[1][16][11] + xor_out[2][16][11] + xor_out[3][16][11] + xor_out[4][16][11];
assign sum_out[1][16][11] = xor_out[5][16][11] + xor_out[6][16][11] + xor_out[7][16][11] + xor_out[8][16][11] + xor_out[9][16][11];
assign sum_out[2][16][11] = xor_out[10][16][11] + xor_out[11][16][11] + xor_out[12][16][11] + xor_out[13][16][11] + xor_out[14][16][11];
assign sum_out[3][16][11] = xor_out[15][16][11] + xor_out[16][16][11] + xor_out[17][16][11] + xor_out[18][16][11] + xor_out[19][16][11];
assign sum_out[4][16][11] = xor_out[20][16][11] + xor_out[21][16][11] + xor_out[22][16][11] + xor_out[23][16][11] + xor_out[24][16][11];
assign sum_out[5][16][11] = xor_out[25][16][11] + xor_out[26][16][11] + xor_out[27][16][11] + xor_out[28][16][11] + xor_out[29][16][11];
assign sum_out[6][16][11] = xor_out[30][16][11] + xor_out[31][16][11] + xor_out[32][16][11] + xor_out[33][16][11] + xor_out[34][16][11];
assign sum_out[7][16][11] = xor_out[35][16][11] + xor_out[36][16][11] + xor_out[37][16][11] + xor_out[38][16][11] + xor_out[39][16][11];
assign sum_out[8][16][11] = xor_out[40][16][11] + xor_out[41][16][11] + xor_out[42][16][11] + xor_out[43][16][11] + xor_out[44][16][11];
assign sum_out[9][16][11] = xor_out[45][16][11] + xor_out[46][16][11] + xor_out[47][16][11] + xor_out[48][16][11] + xor_out[49][16][11];
assign sum_out[10][16][11] = xor_out[50][16][11] + xor_out[51][16][11] + xor_out[52][16][11] + xor_out[53][16][11] + xor_out[54][16][11];
assign sum_out[11][16][11] = xor_out[55][16][11] + xor_out[56][16][11] + xor_out[57][16][11] + xor_out[58][16][11] + xor_out[59][16][11];
assign sum_out[12][16][11] = xor_out[60][16][11] + xor_out[61][16][11] + xor_out[62][16][11] + xor_out[63][16][11] + xor_out[64][16][11];
assign sum_out[13][16][11] = xor_out[65][16][11] + xor_out[66][16][11] + xor_out[67][16][11] + xor_out[68][16][11] + xor_out[69][16][11];
assign sum_out[14][16][11] = xor_out[70][16][11] + xor_out[71][16][11] + xor_out[72][16][11] + xor_out[73][16][11] + xor_out[74][16][11];
assign sum_out[15][16][11] = xor_out[75][16][11] + xor_out[76][16][11] + xor_out[77][16][11] + xor_out[78][16][11] + xor_out[79][16][11];
assign sum_out[16][16][11] = xor_out[80][16][11] + xor_out[81][16][11] + xor_out[82][16][11] + xor_out[83][16][11] + xor_out[84][16][11];
assign sum_out[17][16][11] = xor_out[85][16][11] + xor_out[86][16][11] + xor_out[87][16][11] + xor_out[88][16][11] + xor_out[89][16][11];
assign sum_out[18][16][11] = xor_out[90][16][11] + xor_out[91][16][11] + xor_out[92][16][11] + xor_out[93][16][11] + xor_out[94][16][11];
assign sum_out[19][16][11] = xor_out[95][16][11] + xor_out[96][16][11] + xor_out[97][16][11] + xor_out[98][16][11] + xor_out[99][16][11];

assign sum_out[0][16][12] = xor_out[0][16][12] + xor_out[1][16][12] + xor_out[2][16][12] + xor_out[3][16][12] + xor_out[4][16][12];
assign sum_out[1][16][12] = xor_out[5][16][12] + xor_out[6][16][12] + xor_out[7][16][12] + xor_out[8][16][12] + xor_out[9][16][12];
assign sum_out[2][16][12] = xor_out[10][16][12] + xor_out[11][16][12] + xor_out[12][16][12] + xor_out[13][16][12] + xor_out[14][16][12];
assign sum_out[3][16][12] = xor_out[15][16][12] + xor_out[16][16][12] + xor_out[17][16][12] + xor_out[18][16][12] + xor_out[19][16][12];
assign sum_out[4][16][12] = xor_out[20][16][12] + xor_out[21][16][12] + xor_out[22][16][12] + xor_out[23][16][12] + xor_out[24][16][12];
assign sum_out[5][16][12] = xor_out[25][16][12] + xor_out[26][16][12] + xor_out[27][16][12] + xor_out[28][16][12] + xor_out[29][16][12];
assign sum_out[6][16][12] = xor_out[30][16][12] + xor_out[31][16][12] + xor_out[32][16][12] + xor_out[33][16][12] + xor_out[34][16][12];
assign sum_out[7][16][12] = xor_out[35][16][12] + xor_out[36][16][12] + xor_out[37][16][12] + xor_out[38][16][12] + xor_out[39][16][12];
assign sum_out[8][16][12] = xor_out[40][16][12] + xor_out[41][16][12] + xor_out[42][16][12] + xor_out[43][16][12] + xor_out[44][16][12];
assign sum_out[9][16][12] = xor_out[45][16][12] + xor_out[46][16][12] + xor_out[47][16][12] + xor_out[48][16][12] + xor_out[49][16][12];
assign sum_out[10][16][12] = xor_out[50][16][12] + xor_out[51][16][12] + xor_out[52][16][12] + xor_out[53][16][12] + xor_out[54][16][12];
assign sum_out[11][16][12] = xor_out[55][16][12] + xor_out[56][16][12] + xor_out[57][16][12] + xor_out[58][16][12] + xor_out[59][16][12];
assign sum_out[12][16][12] = xor_out[60][16][12] + xor_out[61][16][12] + xor_out[62][16][12] + xor_out[63][16][12] + xor_out[64][16][12];
assign sum_out[13][16][12] = xor_out[65][16][12] + xor_out[66][16][12] + xor_out[67][16][12] + xor_out[68][16][12] + xor_out[69][16][12];
assign sum_out[14][16][12] = xor_out[70][16][12] + xor_out[71][16][12] + xor_out[72][16][12] + xor_out[73][16][12] + xor_out[74][16][12];
assign sum_out[15][16][12] = xor_out[75][16][12] + xor_out[76][16][12] + xor_out[77][16][12] + xor_out[78][16][12] + xor_out[79][16][12];
assign sum_out[16][16][12] = xor_out[80][16][12] + xor_out[81][16][12] + xor_out[82][16][12] + xor_out[83][16][12] + xor_out[84][16][12];
assign sum_out[17][16][12] = xor_out[85][16][12] + xor_out[86][16][12] + xor_out[87][16][12] + xor_out[88][16][12] + xor_out[89][16][12];
assign sum_out[18][16][12] = xor_out[90][16][12] + xor_out[91][16][12] + xor_out[92][16][12] + xor_out[93][16][12] + xor_out[94][16][12];
assign sum_out[19][16][12] = xor_out[95][16][12] + xor_out[96][16][12] + xor_out[97][16][12] + xor_out[98][16][12] + xor_out[99][16][12];

assign sum_out[0][16][13] = xor_out[0][16][13] + xor_out[1][16][13] + xor_out[2][16][13] + xor_out[3][16][13] + xor_out[4][16][13];
assign sum_out[1][16][13] = xor_out[5][16][13] + xor_out[6][16][13] + xor_out[7][16][13] + xor_out[8][16][13] + xor_out[9][16][13];
assign sum_out[2][16][13] = xor_out[10][16][13] + xor_out[11][16][13] + xor_out[12][16][13] + xor_out[13][16][13] + xor_out[14][16][13];
assign sum_out[3][16][13] = xor_out[15][16][13] + xor_out[16][16][13] + xor_out[17][16][13] + xor_out[18][16][13] + xor_out[19][16][13];
assign sum_out[4][16][13] = xor_out[20][16][13] + xor_out[21][16][13] + xor_out[22][16][13] + xor_out[23][16][13] + xor_out[24][16][13];
assign sum_out[5][16][13] = xor_out[25][16][13] + xor_out[26][16][13] + xor_out[27][16][13] + xor_out[28][16][13] + xor_out[29][16][13];
assign sum_out[6][16][13] = xor_out[30][16][13] + xor_out[31][16][13] + xor_out[32][16][13] + xor_out[33][16][13] + xor_out[34][16][13];
assign sum_out[7][16][13] = xor_out[35][16][13] + xor_out[36][16][13] + xor_out[37][16][13] + xor_out[38][16][13] + xor_out[39][16][13];
assign sum_out[8][16][13] = xor_out[40][16][13] + xor_out[41][16][13] + xor_out[42][16][13] + xor_out[43][16][13] + xor_out[44][16][13];
assign sum_out[9][16][13] = xor_out[45][16][13] + xor_out[46][16][13] + xor_out[47][16][13] + xor_out[48][16][13] + xor_out[49][16][13];
assign sum_out[10][16][13] = xor_out[50][16][13] + xor_out[51][16][13] + xor_out[52][16][13] + xor_out[53][16][13] + xor_out[54][16][13];
assign sum_out[11][16][13] = xor_out[55][16][13] + xor_out[56][16][13] + xor_out[57][16][13] + xor_out[58][16][13] + xor_out[59][16][13];
assign sum_out[12][16][13] = xor_out[60][16][13] + xor_out[61][16][13] + xor_out[62][16][13] + xor_out[63][16][13] + xor_out[64][16][13];
assign sum_out[13][16][13] = xor_out[65][16][13] + xor_out[66][16][13] + xor_out[67][16][13] + xor_out[68][16][13] + xor_out[69][16][13];
assign sum_out[14][16][13] = xor_out[70][16][13] + xor_out[71][16][13] + xor_out[72][16][13] + xor_out[73][16][13] + xor_out[74][16][13];
assign sum_out[15][16][13] = xor_out[75][16][13] + xor_out[76][16][13] + xor_out[77][16][13] + xor_out[78][16][13] + xor_out[79][16][13];
assign sum_out[16][16][13] = xor_out[80][16][13] + xor_out[81][16][13] + xor_out[82][16][13] + xor_out[83][16][13] + xor_out[84][16][13];
assign sum_out[17][16][13] = xor_out[85][16][13] + xor_out[86][16][13] + xor_out[87][16][13] + xor_out[88][16][13] + xor_out[89][16][13];
assign sum_out[18][16][13] = xor_out[90][16][13] + xor_out[91][16][13] + xor_out[92][16][13] + xor_out[93][16][13] + xor_out[94][16][13];
assign sum_out[19][16][13] = xor_out[95][16][13] + xor_out[96][16][13] + xor_out[97][16][13] + xor_out[98][16][13] + xor_out[99][16][13];

assign sum_out[0][16][14] = xor_out[0][16][14] + xor_out[1][16][14] + xor_out[2][16][14] + xor_out[3][16][14] + xor_out[4][16][14];
assign sum_out[1][16][14] = xor_out[5][16][14] + xor_out[6][16][14] + xor_out[7][16][14] + xor_out[8][16][14] + xor_out[9][16][14];
assign sum_out[2][16][14] = xor_out[10][16][14] + xor_out[11][16][14] + xor_out[12][16][14] + xor_out[13][16][14] + xor_out[14][16][14];
assign sum_out[3][16][14] = xor_out[15][16][14] + xor_out[16][16][14] + xor_out[17][16][14] + xor_out[18][16][14] + xor_out[19][16][14];
assign sum_out[4][16][14] = xor_out[20][16][14] + xor_out[21][16][14] + xor_out[22][16][14] + xor_out[23][16][14] + xor_out[24][16][14];
assign sum_out[5][16][14] = xor_out[25][16][14] + xor_out[26][16][14] + xor_out[27][16][14] + xor_out[28][16][14] + xor_out[29][16][14];
assign sum_out[6][16][14] = xor_out[30][16][14] + xor_out[31][16][14] + xor_out[32][16][14] + xor_out[33][16][14] + xor_out[34][16][14];
assign sum_out[7][16][14] = xor_out[35][16][14] + xor_out[36][16][14] + xor_out[37][16][14] + xor_out[38][16][14] + xor_out[39][16][14];
assign sum_out[8][16][14] = xor_out[40][16][14] + xor_out[41][16][14] + xor_out[42][16][14] + xor_out[43][16][14] + xor_out[44][16][14];
assign sum_out[9][16][14] = xor_out[45][16][14] + xor_out[46][16][14] + xor_out[47][16][14] + xor_out[48][16][14] + xor_out[49][16][14];
assign sum_out[10][16][14] = xor_out[50][16][14] + xor_out[51][16][14] + xor_out[52][16][14] + xor_out[53][16][14] + xor_out[54][16][14];
assign sum_out[11][16][14] = xor_out[55][16][14] + xor_out[56][16][14] + xor_out[57][16][14] + xor_out[58][16][14] + xor_out[59][16][14];
assign sum_out[12][16][14] = xor_out[60][16][14] + xor_out[61][16][14] + xor_out[62][16][14] + xor_out[63][16][14] + xor_out[64][16][14];
assign sum_out[13][16][14] = xor_out[65][16][14] + xor_out[66][16][14] + xor_out[67][16][14] + xor_out[68][16][14] + xor_out[69][16][14];
assign sum_out[14][16][14] = xor_out[70][16][14] + xor_out[71][16][14] + xor_out[72][16][14] + xor_out[73][16][14] + xor_out[74][16][14];
assign sum_out[15][16][14] = xor_out[75][16][14] + xor_out[76][16][14] + xor_out[77][16][14] + xor_out[78][16][14] + xor_out[79][16][14];
assign sum_out[16][16][14] = xor_out[80][16][14] + xor_out[81][16][14] + xor_out[82][16][14] + xor_out[83][16][14] + xor_out[84][16][14];
assign sum_out[17][16][14] = xor_out[85][16][14] + xor_out[86][16][14] + xor_out[87][16][14] + xor_out[88][16][14] + xor_out[89][16][14];
assign sum_out[18][16][14] = xor_out[90][16][14] + xor_out[91][16][14] + xor_out[92][16][14] + xor_out[93][16][14] + xor_out[94][16][14];
assign sum_out[19][16][14] = xor_out[95][16][14] + xor_out[96][16][14] + xor_out[97][16][14] + xor_out[98][16][14] + xor_out[99][16][14];

assign sum_out[0][16][15] = xor_out[0][16][15] + xor_out[1][16][15] + xor_out[2][16][15] + xor_out[3][16][15] + xor_out[4][16][15];
assign sum_out[1][16][15] = xor_out[5][16][15] + xor_out[6][16][15] + xor_out[7][16][15] + xor_out[8][16][15] + xor_out[9][16][15];
assign sum_out[2][16][15] = xor_out[10][16][15] + xor_out[11][16][15] + xor_out[12][16][15] + xor_out[13][16][15] + xor_out[14][16][15];
assign sum_out[3][16][15] = xor_out[15][16][15] + xor_out[16][16][15] + xor_out[17][16][15] + xor_out[18][16][15] + xor_out[19][16][15];
assign sum_out[4][16][15] = xor_out[20][16][15] + xor_out[21][16][15] + xor_out[22][16][15] + xor_out[23][16][15] + xor_out[24][16][15];
assign sum_out[5][16][15] = xor_out[25][16][15] + xor_out[26][16][15] + xor_out[27][16][15] + xor_out[28][16][15] + xor_out[29][16][15];
assign sum_out[6][16][15] = xor_out[30][16][15] + xor_out[31][16][15] + xor_out[32][16][15] + xor_out[33][16][15] + xor_out[34][16][15];
assign sum_out[7][16][15] = xor_out[35][16][15] + xor_out[36][16][15] + xor_out[37][16][15] + xor_out[38][16][15] + xor_out[39][16][15];
assign sum_out[8][16][15] = xor_out[40][16][15] + xor_out[41][16][15] + xor_out[42][16][15] + xor_out[43][16][15] + xor_out[44][16][15];
assign sum_out[9][16][15] = xor_out[45][16][15] + xor_out[46][16][15] + xor_out[47][16][15] + xor_out[48][16][15] + xor_out[49][16][15];
assign sum_out[10][16][15] = xor_out[50][16][15] + xor_out[51][16][15] + xor_out[52][16][15] + xor_out[53][16][15] + xor_out[54][16][15];
assign sum_out[11][16][15] = xor_out[55][16][15] + xor_out[56][16][15] + xor_out[57][16][15] + xor_out[58][16][15] + xor_out[59][16][15];
assign sum_out[12][16][15] = xor_out[60][16][15] + xor_out[61][16][15] + xor_out[62][16][15] + xor_out[63][16][15] + xor_out[64][16][15];
assign sum_out[13][16][15] = xor_out[65][16][15] + xor_out[66][16][15] + xor_out[67][16][15] + xor_out[68][16][15] + xor_out[69][16][15];
assign sum_out[14][16][15] = xor_out[70][16][15] + xor_out[71][16][15] + xor_out[72][16][15] + xor_out[73][16][15] + xor_out[74][16][15];
assign sum_out[15][16][15] = xor_out[75][16][15] + xor_out[76][16][15] + xor_out[77][16][15] + xor_out[78][16][15] + xor_out[79][16][15];
assign sum_out[16][16][15] = xor_out[80][16][15] + xor_out[81][16][15] + xor_out[82][16][15] + xor_out[83][16][15] + xor_out[84][16][15];
assign sum_out[17][16][15] = xor_out[85][16][15] + xor_out[86][16][15] + xor_out[87][16][15] + xor_out[88][16][15] + xor_out[89][16][15];
assign sum_out[18][16][15] = xor_out[90][16][15] + xor_out[91][16][15] + xor_out[92][16][15] + xor_out[93][16][15] + xor_out[94][16][15];
assign sum_out[19][16][15] = xor_out[95][16][15] + xor_out[96][16][15] + xor_out[97][16][15] + xor_out[98][16][15] + xor_out[99][16][15];

assign sum_out[0][16][16] = xor_out[0][16][16] + xor_out[1][16][16] + xor_out[2][16][16] + xor_out[3][16][16] + xor_out[4][16][16];
assign sum_out[1][16][16] = xor_out[5][16][16] + xor_out[6][16][16] + xor_out[7][16][16] + xor_out[8][16][16] + xor_out[9][16][16];
assign sum_out[2][16][16] = xor_out[10][16][16] + xor_out[11][16][16] + xor_out[12][16][16] + xor_out[13][16][16] + xor_out[14][16][16];
assign sum_out[3][16][16] = xor_out[15][16][16] + xor_out[16][16][16] + xor_out[17][16][16] + xor_out[18][16][16] + xor_out[19][16][16];
assign sum_out[4][16][16] = xor_out[20][16][16] + xor_out[21][16][16] + xor_out[22][16][16] + xor_out[23][16][16] + xor_out[24][16][16];
assign sum_out[5][16][16] = xor_out[25][16][16] + xor_out[26][16][16] + xor_out[27][16][16] + xor_out[28][16][16] + xor_out[29][16][16];
assign sum_out[6][16][16] = xor_out[30][16][16] + xor_out[31][16][16] + xor_out[32][16][16] + xor_out[33][16][16] + xor_out[34][16][16];
assign sum_out[7][16][16] = xor_out[35][16][16] + xor_out[36][16][16] + xor_out[37][16][16] + xor_out[38][16][16] + xor_out[39][16][16];
assign sum_out[8][16][16] = xor_out[40][16][16] + xor_out[41][16][16] + xor_out[42][16][16] + xor_out[43][16][16] + xor_out[44][16][16];
assign sum_out[9][16][16] = xor_out[45][16][16] + xor_out[46][16][16] + xor_out[47][16][16] + xor_out[48][16][16] + xor_out[49][16][16];
assign sum_out[10][16][16] = xor_out[50][16][16] + xor_out[51][16][16] + xor_out[52][16][16] + xor_out[53][16][16] + xor_out[54][16][16];
assign sum_out[11][16][16] = xor_out[55][16][16] + xor_out[56][16][16] + xor_out[57][16][16] + xor_out[58][16][16] + xor_out[59][16][16];
assign sum_out[12][16][16] = xor_out[60][16][16] + xor_out[61][16][16] + xor_out[62][16][16] + xor_out[63][16][16] + xor_out[64][16][16];
assign sum_out[13][16][16] = xor_out[65][16][16] + xor_out[66][16][16] + xor_out[67][16][16] + xor_out[68][16][16] + xor_out[69][16][16];
assign sum_out[14][16][16] = xor_out[70][16][16] + xor_out[71][16][16] + xor_out[72][16][16] + xor_out[73][16][16] + xor_out[74][16][16];
assign sum_out[15][16][16] = xor_out[75][16][16] + xor_out[76][16][16] + xor_out[77][16][16] + xor_out[78][16][16] + xor_out[79][16][16];
assign sum_out[16][16][16] = xor_out[80][16][16] + xor_out[81][16][16] + xor_out[82][16][16] + xor_out[83][16][16] + xor_out[84][16][16];
assign sum_out[17][16][16] = xor_out[85][16][16] + xor_out[86][16][16] + xor_out[87][16][16] + xor_out[88][16][16] + xor_out[89][16][16];
assign sum_out[18][16][16] = xor_out[90][16][16] + xor_out[91][16][16] + xor_out[92][16][16] + xor_out[93][16][16] + xor_out[94][16][16];
assign sum_out[19][16][16] = xor_out[95][16][16] + xor_out[96][16][16] + xor_out[97][16][16] + xor_out[98][16][16] + xor_out[99][16][16];

assign sum_out[0][16][17] = xor_out[0][16][17] + xor_out[1][16][17] + xor_out[2][16][17] + xor_out[3][16][17] + xor_out[4][16][17];
assign sum_out[1][16][17] = xor_out[5][16][17] + xor_out[6][16][17] + xor_out[7][16][17] + xor_out[8][16][17] + xor_out[9][16][17];
assign sum_out[2][16][17] = xor_out[10][16][17] + xor_out[11][16][17] + xor_out[12][16][17] + xor_out[13][16][17] + xor_out[14][16][17];
assign sum_out[3][16][17] = xor_out[15][16][17] + xor_out[16][16][17] + xor_out[17][16][17] + xor_out[18][16][17] + xor_out[19][16][17];
assign sum_out[4][16][17] = xor_out[20][16][17] + xor_out[21][16][17] + xor_out[22][16][17] + xor_out[23][16][17] + xor_out[24][16][17];
assign sum_out[5][16][17] = xor_out[25][16][17] + xor_out[26][16][17] + xor_out[27][16][17] + xor_out[28][16][17] + xor_out[29][16][17];
assign sum_out[6][16][17] = xor_out[30][16][17] + xor_out[31][16][17] + xor_out[32][16][17] + xor_out[33][16][17] + xor_out[34][16][17];
assign sum_out[7][16][17] = xor_out[35][16][17] + xor_out[36][16][17] + xor_out[37][16][17] + xor_out[38][16][17] + xor_out[39][16][17];
assign sum_out[8][16][17] = xor_out[40][16][17] + xor_out[41][16][17] + xor_out[42][16][17] + xor_out[43][16][17] + xor_out[44][16][17];
assign sum_out[9][16][17] = xor_out[45][16][17] + xor_out[46][16][17] + xor_out[47][16][17] + xor_out[48][16][17] + xor_out[49][16][17];
assign sum_out[10][16][17] = xor_out[50][16][17] + xor_out[51][16][17] + xor_out[52][16][17] + xor_out[53][16][17] + xor_out[54][16][17];
assign sum_out[11][16][17] = xor_out[55][16][17] + xor_out[56][16][17] + xor_out[57][16][17] + xor_out[58][16][17] + xor_out[59][16][17];
assign sum_out[12][16][17] = xor_out[60][16][17] + xor_out[61][16][17] + xor_out[62][16][17] + xor_out[63][16][17] + xor_out[64][16][17];
assign sum_out[13][16][17] = xor_out[65][16][17] + xor_out[66][16][17] + xor_out[67][16][17] + xor_out[68][16][17] + xor_out[69][16][17];
assign sum_out[14][16][17] = xor_out[70][16][17] + xor_out[71][16][17] + xor_out[72][16][17] + xor_out[73][16][17] + xor_out[74][16][17];
assign sum_out[15][16][17] = xor_out[75][16][17] + xor_out[76][16][17] + xor_out[77][16][17] + xor_out[78][16][17] + xor_out[79][16][17];
assign sum_out[16][16][17] = xor_out[80][16][17] + xor_out[81][16][17] + xor_out[82][16][17] + xor_out[83][16][17] + xor_out[84][16][17];
assign sum_out[17][16][17] = xor_out[85][16][17] + xor_out[86][16][17] + xor_out[87][16][17] + xor_out[88][16][17] + xor_out[89][16][17];
assign sum_out[18][16][17] = xor_out[90][16][17] + xor_out[91][16][17] + xor_out[92][16][17] + xor_out[93][16][17] + xor_out[94][16][17];
assign sum_out[19][16][17] = xor_out[95][16][17] + xor_out[96][16][17] + xor_out[97][16][17] + xor_out[98][16][17] + xor_out[99][16][17];

assign sum_out[0][16][18] = xor_out[0][16][18] + xor_out[1][16][18] + xor_out[2][16][18] + xor_out[3][16][18] + xor_out[4][16][18];
assign sum_out[1][16][18] = xor_out[5][16][18] + xor_out[6][16][18] + xor_out[7][16][18] + xor_out[8][16][18] + xor_out[9][16][18];
assign sum_out[2][16][18] = xor_out[10][16][18] + xor_out[11][16][18] + xor_out[12][16][18] + xor_out[13][16][18] + xor_out[14][16][18];
assign sum_out[3][16][18] = xor_out[15][16][18] + xor_out[16][16][18] + xor_out[17][16][18] + xor_out[18][16][18] + xor_out[19][16][18];
assign sum_out[4][16][18] = xor_out[20][16][18] + xor_out[21][16][18] + xor_out[22][16][18] + xor_out[23][16][18] + xor_out[24][16][18];
assign sum_out[5][16][18] = xor_out[25][16][18] + xor_out[26][16][18] + xor_out[27][16][18] + xor_out[28][16][18] + xor_out[29][16][18];
assign sum_out[6][16][18] = xor_out[30][16][18] + xor_out[31][16][18] + xor_out[32][16][18] + xor_out[33][16][18] + xor_out[34][16][18];
assign sum_out[7][16][18] = xor_out[35][16][18] + xor_out[36][16][18] + xor_out[37][16][18] + xor_out[38][16][18] + xor_out[39][16][18];
assign sum_out[8][16][18] = xor_out[40][16][18] + xor_out[41][16][18] + xor_out[42][16][18] + xor_out[43][16][18] + xor_out[44][16][18];
assign sum_out[9][16][18] = xor_out[45][16][18] + xor_out[46][16][18] + xor_out[47][16][18] + xor_out[48][16][18] + xor_out[49][16][18];
assign sum_out[10][16][18] = xor_out[50][16][18] + xor_out[51][16][18] + xor_out[52][16][18] + xor_out[53][16][18] + xor_out[54][16][18];
assign sum_out[11][16][18] = xor_out[55][16][18] + xor_out[56][16][18] + xor_out[57][16][18] + xor_out[58][16][18] + xor_out[59][16][18];
assign sum_out[12][16][18] = xor_out[60][16][18] + xor_out[61][16][18] + xor_out[62][16][18] + xor_out[63][16][18] + xor_out[64][16][18];
assign sum_out[13][16][18] = xor_out[65][16][18] + xor_out[66][16][18] + xor_out[67][16][18] + xor_out[68][16][18] + xor_out[69][16][18];
assign sum_out[14][16][18] = xor_out[70][16][18] + xor_out[71][16][18] + xor_out[72][16][18] + xor_out[73][16][18] + xor_out[74][16][18];
assign sum_out[15][16][18] = xor_out[75][16][18] + xor_out[76][16][18] + xor_out[77][16][18] + xor_out[78][16][18] + xor_out[79][16][18];
assign sum_out[16][16][18] = xor_out[80][16][18] + xor_out[81][16][18] + xor_out[82][16][18] + xor_out[83][16][18] + xor_out[84][16][18];
assign sum_out[17][16][18] = xor_out[85][16][18] + xor_out[86][16][18] + xor_out[87][16][18] + xor_out[88][16][18] + xor_out[89][16][18];
assign sum_out[18][16][18] = xor_out[90][16][18] + xor_out[91][16][18] + xor_out[92][16][18] + xor_out[93][16][18] + xor_out[94][16][18];
assign sum_out[19][16][18] = xor_out[95][16][18] + xor_out[96][16][18] + xor_out[97][16][18] + xor_out[98][16][18] + xor_out[99][16][18];

assign sum_out[0][16][19] = xor_out[0][16][19] + xor_out[1][16][19] + xor_out[2][16][19] + xor_out[3][16][19] + xor_out[4][16][19];
assign sum_out[1][16][19] = xor_out[5][16][19] + xor_out[6][16][19] + xor_out[7][16][19] + xor_out[8][16][19] + xor_out[9][16][19];
assign sum_out[2][16][19] = xor_out[10][16][19] + xor_out[11][16][19] + xor_out[12][16][19] + xor_out[13][16][19] + xor_out[14][16][19];
assign sum_out[3][16][19] = xor_out[15][16][19] + xor_out[16][16][19] + xor_out[17][16][19] + xor_out[18][16][19] + xor_out[19][16][19];
assign sum_out[4][16][19] = xor_out[20][16][19] + xor_out[21][16][19] + xor_out[22][16][19] + xor_out[23][16][19] + xor_out[24][16][19];
assign sum_out[5][16][19] = xor_out[25][16][19] + xor_out[26][16][19] + xor_out[27][16][19] + xor_out[28][16][19] + xor_out[29][16][19];
assign sum_out[6][16][19] = xor_out[30][16][19] + xor_out[31][16][19] + xor_out[32][16][19] + xor_out[33][16][19] + xor_out[34][16][19];
assign sum_out[7][16][19] = xor_out[35][16][19] + xor_out[36][16][19] + xor_out[37][16][19] + xor_out[38][16][19] + xor_out[39][16][19];
assign sum_out[8][16][19] = xor_out[40][16][19] + xor_out[41][16][19] + xor_out[42][16][19] + xor_out[43][16][19] + xor_out[44][16][19];
assign sum_out[9][16][19] = xor_out[45][16][19] + xor_out[46][16][19] + xor_out[47][16][19] + xor_out[48][16][19] + xor_out[49][16][19];
assign sum_out[10][16][19] = xor_out[50][16][19] + xor_out[51][16][19] + xor_out[52][16][19] + xor_out[53][16][19] + xor_out[54][16][19];
assign sum_out[11][16][19] = xor_out[55][16][19] + xor_out[56][16][19] + xor_out[57][16][19] + xor_out[58][16][19] + xor_out[59][16][19];
assign sum_out[12][16][19] = xor_out[60][16][19] + xor_out[61][16][19] + xor_out[62][16][19] + xor_out[63][16][19] + xor_out[64][16][19];
assign sum_out[13][16][19] = xor_out[65][16][19] + xor_out[66][16][19] + xor_out[67][16][19] + xor_out[68][16][19] + xor_out[69][16][19];
assign sum_out[14][16][19] = xor_out[70][16][19] + xor_out[71][16][19] + xor_out[72][16][19] + xor_out[73][16][19] + xor_out[74][16][19];
assign sum_out[15][16][19] = xor_out[75][16][19] + xor_out[76][16][19] + xor_out[77][16][19] + xor_out[78][16][19] + xor_out[79][16][19];
assign sum_out[16][16][19] = xor_out[80][16][19] + xor_out[81][16][19] + xor_out[82][16][19] + xor_out[83][16][19] + xor_out[84][16][19];
assign sum_out[17][16][19] = xor_out[85][16][19] + xor_out[86][16][19] + xor_out[87][16][19] + xor_out[88][16][19] + xor_out[89][16][19];
assign sum_out[18][16][19] = xor_out[90][16][19] + xor_out[91][16][19] + xor_out[92][16][19] + xor_out[93][16][19] + xor_out[94][16][19];
assign sum_out[19][16][19] = xor_out[95][16][19] + xor_out[96][16][19] + xor_out[97][16][19] + xor_out[98][16][19] + xor_out[99][16][19];

assign sum_out[0][16][20] = xor_out[0][16][20] + xor_out[1][16][20] + xor_out[2][16][20] + xor_out[3][16][20] + xor_out[4][16][20];
assign sum_out[1][16][20] = xor_out[5][16][20] + xor_out[6][16][20] + xor_out[7][16][20] + xor_out[8][16][20] + xor_out[9][16][20];
assign sum_out[2][16][20] = xor_out[10][16][20] + xor_out[11][16][20] + xor_out[12][16][20] + xor_out[13][16][20] + xor_out[14][16][20];
assign sum_out[3][16][20] = xor_out[15][16][20] + xor_out[16][16][20] + xor_out[17][16][20] + xor_out[18][16][20] + xor_out[19][16][20];
assign sum_out[4][16][20] = xor_out[20][16][20] + xor_out[21][16][20] + xor_out[22][16][20] + xor_out[23][16][20] + xor_out[24][16][20];
assign sum_out[5][16][20] = xor_out[25][16][20] + xor_out[26][16][20] + xor_out[27][16][20] + xor_out[28][16][20] + xor_out[29][16][20];
assign sum_out[6][16][20] = xor_out[30][16][20] + xor_out[31][16][20] + xor_out[32][16][20] + xor_out[33][16][20] + xor_out[34][16][20];
assign sum_out[7][16][20] = xor_out[35][16][20] + xor_out[36][16][20] + xor_out[37][16][20] + xor_out[38][16][20] + xor_out[39][16][20];
assign sum_out[8][16][20] = xor_out[40][16][20] + xor_out[41][16][20] + xor_out[42][16][20] + xor_out[43][16][20] + xor_out[44][16][20];
assign sum_out[9][16][20] = xor_out[45][16][20] + xor_out[46][16][20] + xor_out[47][16][20] + xor_out[48][16][20] + xor_out[49][16][20];
assign sum_out[10][16][20] = xor_out[50][16][20] + xor_out[51][16][20] + xor_out[52][16][20] + xor_out[53][16][20] + xor_out[54][16][20];
assign sum_out[11][16][20] = xor_out[55][16][20] + xor_out[56][16][20] + xor_out[57][16][20] + xor_out[58][16][20] + xor_out[59][16][20];
assign sum_out[12][16][20] = xor_out[60][16][20] + xor_out[61][16][20] + xor_out[62][16][20] + xor_out[63][16][20] + xor_out[64][16][20];
assign sum_out[13][16][20] = xor_out[65][16][20] + xor_out[66][16][20] + xor_out[67][16][20] + xor_out[68][16][20] + xor_out[69][16][20];
assign sum_out[14][16][20] = xor_out[70][16][20] + xor_out[71][16][20] + xor_out[72][16][20] + xor_out[73][16][20] + xor_out[74][16][20];
assign sum_out[15][16][20] = xor_out[75][16][20] + xor_out[76][16][20] + xor_out[77][16][20] + xor_out[78][16][20] + xor_out[79][16][20];
assign sum_out[16][16][20] = xor_out[80][16][20] + xor_out[81][16][20] + xor_out[82][16][20] + xor_out[83][16][20] + xor_out[84][16][20];
assign sum_out[17][16][20] = xor_out[85][16][20] + xor_out[86][16][20] + xor_out[87][16][20] + xor_out[88][16][20] + xor_out[89][16][20];
assign sum_out[18][16][20] = xor_out[90][16][20] + xor_out[91][16][20] + xor_out[92][16][20] + xor_out[93][16][20] + xor_out[94][16][20];
assign sum_out[19][16][20] = xor_out[95][16][20] + xor_out[96][16][20] + xor_out[97][16][20] + xor_out[98][16][20] + xor_out[99][16][20];

assign sum_out[0][16][21] = xor_out[0][16][21] + xor_out[1][16][21] + xor_out[2][16][21] + xor_out[3][16][21] + xor_out[4][16][21];
assign sum_out[1][16][21] = xor_out[5][16][21] + xor_out[6][16][21] + xor_out[7][16][21] + xor_out[8][16][21] + xor_out[9][16][21];
assign sum_out[2][16][21] = xor_out[10][16][21] + xor_out[11][16][21] + xor_out[12][16][21] + xor_out[13][16][21] + xor_out[14][16][21];
assign sum_out[3][16][21] = xor_out[15][16][21] + xor_out[16][16][21] + xor_out[17][16][21] + xor_out[18][16][21] + xor_out[19][16][21];
assign sum_out[4][16][21] = xor_out[20][16][21] + xor_out[21][16][21] + xor_out[22][16][21] + xor_out[23][16][21] + xor_out[24][16][21];
assign sum_out[5][16][21] = xor_out[25][16][21] + xor_out[26][16][21] + xor_out[27][16][21] + xor_out[28][16][21] + xor_out[29][16][21];
assign sum_out[6][16][21] = xor_out[30][16][21] + xor_out[31][16][21] + xor_out[32][16][21] + xor_out[33][16][21] + xor_out[34][16][21];
assign sum_out[7][16][21] = xor_out[35][16][21] + xor_out[36][16][21] + xor_out[37][16][21] + xor_out[38][16][21] + xor_out[39][16][21];
assign sum_out[8][16][21] = xor_out[40][16][21] + xor_out[41][16][21] + xor_out[42][16][21] + xor_out[43][16][21] + xor_out[44][16][21];
assign sum_out[9][16][21] = xor_out[45][16][21] + xor_out[46][16][21] + xor_out[47][16][21] + xor_out[48][16][21] + xor_out[49][16][21];
assign sum_out[10][16][21] = xor_out[50][16][21] + xor_out[51][16][21] + xor_out[52][16][21] + xor_out[53][16][21] + xor_out[54][16][21];
assign sum_out[11][16][21] = xor_out[55][16][21] + xor_out[56][16][21] + xor_out[57][16][21] + xor_out[58][16][21] + xor_out[59][16][21];
assign sum_out[12][16][21] = xor_out[60][16][21] + xor_out[61][16][21] + xor_out[62][16][21] + xor_out[63][16][21] + xor_out[64][16][21];
assign sum_out[13][16][21] = xor_out[65][16][21] + xor_out[66][16][21] + xor_out[67][16][21] + xor_out[68][16][21] + xor_out[69][16][21];
assign sum_out[14][16][21] = xor_out[70][16][21] + xor_out[71][16][21] + xor_out[72][16][21] + xor_out[73][16][21] + xor_out[74][16][21];
assign sum_out[15][16][21] = xor_out[75][16][21] + xor_out[76][16][21] + xor_out[77][16][21] + xor_out[78][16][21] + xor_out[79][16][21];
assign sum_out[16][16][21] = xor_out[80][16][21] + xor_out[81][16][21] + xor_out[82][16][21] + xor_out[83][16][21] + xor_out[84][16][21];
assign sum_out[17][16][21] = xor_out[85][16][21] + xor_out[86][16][21] + xor_out[87][16][21] + xor_out[88][16][21] + xor_out[89][16][21];
assign sum_out[18][16][21] = xor_out[90][16][21] + xor_out[91][16][21] + xor_out[92][16][21] + xor_out[93][16][21] + xor_out[94][16][21];
assign sum_out[19][16][21] = xor_out[95][16][21] + xor_out[96][16][21] + xor_out[97][16][21] + xor_out[98][16][21] + xor_out[99][16][21];

assign sum_out[0][16][22] = xor_out[0][16][22] + xor_out[1][16][22] + xor_out[2][16][22] + xor_out[3][16][22] + xor_out[4][16][22];
assign sum_out[1][16][22] = xor_out[5][16][22] + xor_out[6][16][22] + xor_out[7][16][22] + xor_out[8][16][22] + xor_out[9][16][22];
assign sum_out[2][16][22] = xor_out[10][16][22] + xor_out[11][16][22] + xor_out[12][16][22] + xor_out[13][16][22] + xor_out[14][16][22];
assign sum_out[3][16][22] = xor_out[15][16][22] + xor_out[16][16][22] + xor_out[17][16][22] + xor_out[18][16][22] + xor_out[19][16][22];
assign sum_out[4][16][22] = xor_out[20][16][22] + xor_out[21][16][22] + xor_out[22][16][22] + xor_out[23][16][22] + xor_out[24][16][22];
assign sum_out[5][16][22] = xor_out[25][16][22] + xor_out[26][16][22] + xor_out[27][16][22] + xor_out[28][16][22] + xor_out[29][16][22];
assign sum_out[6][16][22] = xor_out[30][16][22] + xor_out[31][16][22] + xor_out[32][16][22] + xor_out[33][16][22] + xor_out[34][16][22];
assign sum_out[7][16][22] = xor_out[35][16][22] + xor_out[36][16][22] + xor_out[37][16][22] + xor_out[38][16][22] + xor_out[39][16][22];
assign sum_out[8][16][22] = xor_out[40][16][22] + xor_out[41][16][22] + xor_out[42][16][22] + xor_out[43][16][22] + xor_out[44][16][22];
assign sum_out[9][16][22] = xor_out[45][16][22] + xor_out[46][16][22] + xor_out[47][16][22] + xor_out[48][16][22] + xor_out[49][16][22];
assign sum_out[10][16][22] = xor_out[50][16][22] + xor_out[51][16][22] + xor_out[52][16][22] + xor_out[53][16][22] + xor_out[54][16][22];
assign sum_out[11][16][22] = xor_out[55][16][22] + xor_out[56][16][22] + xor_out[57][16][22] + xor_out[58][16][22] + xor_out[59][16][22];
assign sum_out[12][16][22] = xor_out[60][16][22] + xor_out[61][16][22] + xor_out[62][16][22] + xor_out[63][16][22] + xor_out[64][16][22];
assign sum_out[13][16][22] = xor_out[65][16][22] + xor_out[66][16][22] + xor_out[67][16][22] + xor_out[68][16][22] + xor_out[69][16][22];
assign sum_out[14][16][22] = xor_out[70][16][22] + xor_out[71][16][22] + xor_out[72][16][22] + xor_out[73][16][22] + xor_out[74][16][22];
assign sum_out[15][16][22] = xor_out[75][16][22] + xor_out[76][16][22] + xor_out[77][16][22] + xor_out[78][16][22] + xor_out[79][16][22];
assign sum_out[16][16][22] = xor_out[80][16][22] + xor_out[81][16][22] + xor_out[82][16][22] + xor_out[83][16][22] + xor_out[84][16][22];
assign sum_out[17][16][22] = xor_out[85][16][22] + xor_out[86][16][22] + xor_out[87][16][22] + xor_out[88][16][22] + xor_out[89][16][22];
assign sum_out[18][16][22] = xor_out[90][16][22] + xor_out[91][16][22] + xor_out[92][16][22] + xor_out[93][16][22] + xor_out[94][16][22];
assign sum_out[19][16][22] = xor_out[95][16][22] + xor_out[96][16][22] + xor_out[97][16][22] + xor_out[98][16][22] + xor_out[99][16][22];

assign sum_out[0][16][23] = xor_out[0][16][23] + xor_out[1][16][23] + xor_out[2][16][23] + xor_out[3][16][23] + xor_out[4][16][23];
assign sum_out[1][16][23] = xor_out[5][16][23] + xor_out[6][16][23] + xor_out[7][16][23] + xor_out[8][16][23] + xor_out[9][16][23];
assign sum_out[2][16][23] = xor_out[10][16][23] + xor_out[11][16][23] + xor_out[12][16][23] + xor_out[13][16][23] + xor_out[14][16][23];
assign sum_out[3][16][23] = xor_out[15][16][23] + xor_out[16][16][23] + xor_out[17][16][23] + xor_out[18][16][23] + xor_out[19][16][23];
assign sum_out[4][16][23] = xor_out[20][16][23] + xor_out[21][16][23] + xor_out[22][16][23] + xor_out[23][16][23] + xor_out[24][16][23];
assign sum_out[5][16][23] = xor_out[25][16][23] + xor_out[26][16][23] + xor_out[27][16][23] + xor_out[28][16][23] + xor_out[29][16][23];
assign sum_out[6][16][23] = xor_out[30][16][23] + xor_out[31][16][23] + xor_out[32][16][23] + xor_out[33][16][23] + xor_out[34][16][23];
assign sum_out[7][16][23] = xor_out[35][16][23] + xor_out[36][16][23] + xor_out[37][16][23] + xor_out[38][16][23] + xor_out[39][16][23];
assign sum_out[8][16][23] = xor_out[40][16][23] + xor_out[41][16][23] + xor_out[42][16][23] + xor_out[43][16][23] + xor_out[44][16][23];
assign sum_out[9][16][23] = xor_out[45][16][23] + xor_out[46][16][23] + xor_out[47][16][23] + xor_out[48][16][23] + xor_out[49][16][23];
assign sum_out[10][16][23] = xor_out[50][16][23] + xor_out[51][16][23] + xor_out[52][16][23] + xor_out[53][16][23] + xor_out[54][16][23];
assign sum_out[11][16][23] = xor_out[55][16][23] + xor_out[56][16][23] + xor_out[57][16][23] + xor_out[58][16][23] + xor_out[59][16][23];
assign sum_out[12][16][23] = xor_out[60][16][23] + xor_out[61][16][23] + xor_out[62][16][23] + xor_out[63][16][23] + xor_out[64][16][23];
assign sum_out[13][16][23] = xor_out[65][16][23] + xor_out[66][16][23] + xor_out[67][16][23] + xor_out[68][16][23] + xor_out[69][16][23];
assign sum_out[14][16][23] = xor_out[70][16][23] + xor_out[71][16][23] + xor_out[72][16][23] + xor_out[73][16][23] + xor_out[74][16][23];
assign sum_out[15][16][23] = xor_out[75][16][23] + xor_out[76][16][23] + xor_out[77][16][23] + xor_out[78][16][23] + xor_out[79][16][23];
assign sum_out[16][16][23] = xor_out[80][16][23] + xor_out[81][16][23] + xor_out[82][16][23] + xor_out[83][16][23] + xor_out[84][16][23];
assign sum_out[17][16][23] = xor_out[85][16][23] + xor_out[86][16][23] + xor_out[87][16][23] + xor_out[88][16][23] + xor_out[89][16][23];
assign sum_out[18][16][23] = xor_out[90][16][23] + xor_out[91][16][23] + xor_out[92][16][23] + xor_out[93][16][23] + xor_out[94][16][23];
assign sum_out[19][16][23] = xor_out[95][16][23] + xor_out[96][16][23] + xor_out[97][16][23] + xor_out[98][16][23] + xor_out[99][16][23];

assign sum_out[0][17][0] = xor_out[0][17][0] + xor_out[1][17][0] + xor_out[2][17][0] + xor_out[3][17][0] + xor_out[4][17][0];
assign sum_out[1][17][0] = xor_out[5][17][0] + xor_out[6][17][0] + xor_out[7][17][0] + xor_out[8][17][0] + xor_out[9][17][0];
assign sum_out[2][17][0] = xor_out[10][17][0] + xor_out[11][17][0] + xor_out[12][17][0] + xor_out[13][17][0] + xor_out[14][17][0];
assign sum_out[3][17][0] = xor_out[15][17][0] + xor_out[16][17][0] + xor_out[17][17][0] + xor_out[18][17][0] + xor_out[19][17][0];
assign sum_out[4][17][0] = xor_out[20][17][0] + xor_out[21][17][0] + xor_out[22][17][0] + xor_out[23][17][0] + xor_out[24][17][0];
assign sum_out[5][17][0] = xor_out[25][17][0] + xor_out[26][17][0] + xor_out[27][17][0] + xor_out[28][17][0] + xor_out[29][17][0];
assign sum_out[6][17][0] = xor_out[30][17][0] + xor_out[31][17][0] + xor_out[32][17][0] + xor_out[33][17][0] + xor_out[34][17][0];
assign sum_out[7][17][0] = xor_out[35][17][0] + xor_out[36][17][0] + xor_out[37][17][0] + xor_out[38][17][0] + xor_out[39][17][0];
assign sum_out[8][17][0] = xor_out[40][17][0] + xor_out[41][17][0] + xor_out[42][17][0] + xor_out[43][17][0] + xor_out[44][17][0];
assign sum_out[9][17][0] = xor_out[45][17][0] + xor_out[46][17][0] + xor_out[47][17][0] + xor_out[48][17][0] + xor_out[49][17][0];
assign sum_out[10][17][0] = xor_out[50][17][0] + xor_out[51][17][0] + xor_out[52][17][0] + xor_out[53][17][0] + xor_out[54][17][0];
assign sum_out[11][17][0] = xor_out[55][17][0] + xor_out[56][17][0] + xor_out[57][17][0] + xor_out[58][17][0] + xor_out[59][17][0];
assign sum_out[12][17][0] = xor_out[60][17][0] + xor_out[61][17][0] + xor_out[62][17][0] + xor_out[63][17][0] + xor_out[64][17][0];
assign sum_out[13][17][0] = xor_out[65][17][0] + xor_out[66][17][0] + xor_out[67][17][0] + xor_out[68][17][0] + xor_out[69][17][0];
assign sum_out[14][17][0] = xor_out[70][17][0] + xor_out[71][17][0] + xor_out[72][17][0] + xor_out[73][17][0] + xor_out[74][17][0];
assign sum_out[15][17][0] = xor_out[75][17][0] + xor_out[76][17][0] + xor_out[77][17][0] + xor_out[78][17][0] + xor_out[79][17][0];
assign sum_out[16][17][0] = xor_out[80][17][0] + xor_out[81][17][0] + xor_out[82][17][0] + xor_out[83][17][0] + xor_out[84][17][0];
assign sum_out[17][17][0] = xor_out[85][17][0] + xor_out[86][17][0] + xor_out[87][17][0] + xor_out[88][17][0] + xor_out[89][17][0];
assign sum_out[18][17][0] = xor_out[90][17][0] + xor_out[91][17][0] + xor_out[92][17][0] + xor_out[93][17][0] + xor_out[94][17][0];
assign sum_out[19][17][0] = xor_out[95][17][0] + xor_out[96][17][0] + xor_out[97][17][0] + xor_out[98][17][0] + xor_out[99][17][0];

assign sum_out[0][17][1] = xor_out[0][17][1] + xor_out[1][17][1] + xor_out[2][17][1] + xor_out[3][17][1] + xor_out[4][17][1];
assign sum_out[1][17][1] = xor_out[5][17][1] + xor_out[6][17][1] + xor_out[7][17][1] + xor_out[8][17][1] + xor_out[9][17][1];
assign sum_out[2][17][1] = xor_out[10][17][1] + xor_out[11][17][1] + xor_out[12][17][1] + xor_out[13][17][1] + xor_out[14][17][1];
assign sum_out[3][17][1] = xor_out[15][17][1] + xor_out[16][17][1] + xor_out[17][17][1] + xor_out[18][17][1] + xor_out[19][17][1];
assign sum_out[4][17][1] = xor_out[20][17][1] + xor_out[21][17][1] + xor_out[22][17][1] + xor_out[23][17][1] + xor_out[24][17][1];
assign sum_out[5][17][1] = xor_out[25][17][1] + xor_out[26][17][1] + xor_out[27][17][1] + xor_out[28][17][1] + xor_out[29][17][1];
assign sum_out[6][17][1] = xor_out[30][17][1] + xor_out[31][17][1] + xor_out[32][17][1] + xor_out[33][17][1] + xor_out[34][17][1];
assign sum_out[7][17][1] = xor_out[35][17][1] + xor_out[36][17][1] + xor_out[37][17][1] + xor_out[38][17][1] + xor_out[39][17][1];
assign sum_out[8][17][1] = xor_out[40][17][1] + xor_out[41][17][1] + xor_out[42][17][1] + xor_out[43][17][1] + xor_out[44][17][1];
assign sum_out[9][17][1] = xor_out[45][17][1] + xor_out[46][17][1] + xor_out[47][17][1] + xor_out[48][17][1] + xor_out[49][17][1];
assign sum_out[10][17][1] = xor_out[50][17][1] + xor_out[51][17][1] + xor_out[52][17][1] + xor_out[53][17][1] + xor_out[54][17][1];
assign sum_out[11][17][1] = xor_out[55][17][1] + xor_out[56][17][1] + xor_out[57][17][1] + xor_out[58][17][1] + xor_out[59][17][1];
assign sum_out[12][17][1] = xor_out[60][17][1] + xor_out[61][17][1] + xor_out[62][17][1] + xor_out[63][17][1] + xor_out[64][17][1];
assign sum_out[13][17][1] = xor_out[65][17][1] + xor_out[66][17][1] + xor_out[67][17][1] + xor_out[68][17][1] + xor_out[69][17][1];
assign sum_out[14][17][1] = xor_out[70][17][1] + xor_out[71][17][1] + xor_out[72][17][1] + xor_out[73][17][1] + xor_out[74][17][1];
assign sum_out[15][17][1] = xor_out[75][17][1] + xor_out[76][17][1] + xor_out[77][17][1] + xor_out[78][17][1] + xor_out[79][17][1];
assign sum_out[16][17][1] = xor_out[80][17][1] + xor_out[81][17][1] + xor_out[82][17][1] + xor_out[83][17][1] + xor_out[84][17][1];
assign sum_out[17][17][1] = xor_out[85][17][1] + xor_out[86][17][1] + xor_out[87][17][1] + xor_out[88][17][1] + xor_out[89][17][1];
assign sum_out[18][17][1] = xor_out[90][17][1] + xor_out[91][17][1] + xor_out[92][17][1] + xor_out[93][17][1] + xor_out[94][17][1];
assign sum_out[19][17][1] = xor_out[95][17][1] + xor_out[96][17][1] + xor_out[97][17][1] + xor_out[98][17][1] + xor_out[99][17][1];

assign sum_out[0][17][2] = xor_out[0][17][2] + xor_out[1][17][2] + xor_out[2][17][2] + xor_out[3][17][2] + xor_out[4][17][2];
assign sum_out[1][17][2] = xor_out[5][17][2] + xor_out[6][17][2] + xor_out[7][17][2] + xor_out[8][17][2] + xor_out[9][17][2];
assign sum_out[2][17][2] = xor_out[10][17][2] + xor_out[11][17][2] + xor_out[12][17][2] + xor_out[13][17][2] + xor_out[14][17][2];
assign sum_out[3][17][2] = xor_out[15][17][2] + xor_out[16][17][2] + xor_out[17][17][2] + xor_out[18][17][2] + xor_out[19][17][2];
assign sum_out[4][17][2] = xor_out[20][17][2] + xor_out[21][17][2] + xor_out[22][17][2] + xor_out[23][17][2] + xor_out[24][17][2];
assign sum_out[5][17][2] = xor_out[25][17][2] + xor_out[26][17][2] + xor_out[27][17][2] + xor_out[28][17][2] + xor_out[29][17][2];
assign sum_out[6][17][2] = xor_out[30][17][2] + xor_out[31][17][2] + xor_out[32][17][2] + xor_out[33][17][2] + xor_out[34][17][2];
assign sum_out[7][17][2] = xor_out[35][17][2] + xor_out[36][17][2] + xor_out[37][17][2] + xor_out[38][17][2] + xor_out[39][17][2];
assign sum_out[8][17][2] = xor_out[40][17][2] + xor_out[41][17][2] + xor_out[42][17][2] + xor_out[43][17][2] + xor_out[44][17][2];
assign sum_out[9][17][2] = xor_out[45][17][2] + xor_out[46][17][2] + xor_out[47][17][2] + xor_out[48][17][2] + xor_out[49][17][2];
assign sum_out[10][17][2] = xor_out[50][17][2] + xor_out[51][17][2] + xor_out[52][17][2] + xor_out[53][17][2] + xor_out[54][17][2];
assign sum_out[11][17][2] = xor_out[55][17][2] + xor_out[56][17][2] + xor_out[57][17][2] + xor_out[58][17][2] + xor_out[59][17][2];
assign sum_out[12][17][2] = xor_out[60][17][2] + xor_out[61][17][2] + xor_out[62][17][2] + xor_out[63][17][2] + xor_out[64][17][2];
assign sum_out[13][17][2] = xor_out[65][17][2] + xor_out[66][17][2] + xor_out[67][17][2] + xor_out[68][17][2] + xor_out[69][17][2];
assign sum_out[14][17][2] = xor_out[70][17][2] + xor_out[71][17][2] + xor_out[72][17][2] + xor_out[73][17][2] + xor_out[74][17][2];
assign sum_out[15][17][2] = xor_out[75][17][2] + xor_out[76][17][2] + xor_out[77][17][2] + xor_out[78][17][2] + xor_out[79][17][2];
assign sum_out[16][17][2] = xor_out[80][17][2] + xor_out[81][17][2] + xor_out[82][17][2] + xor_out[83][17][2] + xor_out[84][17][2];
assign sum_out[17][17][2] = xor_out[85][17][2] + xor_out[86][17][2] + xor_out[87][17][2] + xor_out[88][17][2] + xor_out[89][17][2];
assign sum_out[18][17][2] = xor_out[90][17][2] + xor_out[91][17][2] + xor_out[92][17][2] + xor_out[93][17][2] + xor_out[94][17][2];
assign sum_out[19][17][2] = xor_out[95][17][2] + xor_out[96][17][2] + xor_out[97][17][2] + xor_out[98][17][2] + xor_out[99][17][2];

assign sum_out[0][17][3] = xor_out[0][17][3] + xor_out[1][17][3] + xor_out[2][17][3] + xor_out[3][17][3] + xor_out[4][17][3];
assign sum_out[1][17][3] = xor_out[5][17][3] + xor_out[6][17][3] + xor_out[7][17][3] + xor_out[8][17][3] + xor_out[9][17][3];
assign sum_out[2][17][3] = xor_out[10][17][3] + xor_out[11][17][3] + xor_out[12][17][3] + xor_out[13][17][3] + xor_out[14][17][3];
assign sum_out[3][17][3] = xor_out[15][17][3] + xor_out[16][17][3] + xor_out[17][17][3] + xor_out[18][17][3] + xor_out[19][17][3];
assign sum_out[4][17][3] = xor_out[20][17][3] + xor_out[21][17][3] + xor_out[22][17][3] + xor_out[23][17][3] + xor_out[24][17][3];
assign sum_out[5][17][3] = xor_out[25][17][3] + xor_out[26][17][3] + xor_out[27][17][3] + xor_out[28][17][3] + xor_out[29][17][3];
assign sum_out[6][17][3] = xor_out[30][17][3] + xor_out[31][17][3] + xor_out[32][17][3] + xor_out[33][17][3] + xor_out[34][17][3];
assign sum_out[7][17][3] = xor_out[35][17][3] + xor_out[36][17][3] + xor_out[37][17][3] + xor_out[38][17][3] + xor_out[39][17][3];
assign sum_out[8][17][3] = xor_out[40][17][3] + xor_out[41][17][3] + xor_out[42][17][3] + xor_out[43][17][3] + xor_out[44][17][3];
assign sum_out[9][17][3] = xor_out[45][17][3] + xor_out[46][17][3] + xor_out[47][17][3] + xor_out[48][17][3] + xor_out[49][17][3];
assign sum_out[10][17][3] = xor_out[50][17][3] + xor_out[51][17][3] + xor_out[52][17][3] + xor_out[53][17][3] + xor_out[54][17][3];
assign sum_out[11][17][3] = xor_out[55][17][3] + xor_out[56][17][3] + xor_out[57][17][3] + xor_out[58][17][3] + xor_out[59][17][3];
assign sum_out[12][17][3] = xor_out[60][17][3] + xor_out[61][17][3] + xor_out[62][17][3] + xor_out[63][17][3] + xor_out[64][17][3];
assign sum_out[13][17][3] = xor_out[65][17][3] + xor_out[66][17][3] + xor_out[67][17][3] + xor_out[68][17][3] + xor_out[69][17][3];
assign sum_out[14][17][3] = xor_out[70][17][3] + xor_out[71][17][3] + xor_out[72][17][3] + xor_out[73][17][3] + xor_out[74][17][3];
assign sum_out[15][17][3] = xor_out[75][17][3] + xor_out[76][17][3] + xor_out[77][17][3] + xor_out[78][17][3] + xor_out[79][17][3];
assign sum_out[16][17][3] = xor_out[80][17][3] + xor_out[81][17][3] + xor_out[82][17][3] + xor_out[83][17][3] + xor_out[84][17][3];
assign sum_out[17][17][3] = xor_out[85][17][3] + xor_out[86][17][3] + xor_out[87][17][3] + xor_out[88][17][3] + xor_out[89][17][3];
assign sum_out[18][17][3] = xor_out[90][17][3] + xor_out[91][17][3] + xor_out[92][17][3] + xor_out[93][17][3] + xor_out[94][17][3];
assign sum_out[19][17][3] = xor_out[95][17][3] + xor_out[96][17][3] + xor_out[97][17][3] + xor_out[98][17][3] + xor_out[99][17][3];

assign sum_out[0][17][4] = xor_out[0][17][4] + xor_out[1][17][4] + xor_out[2][17][4] + xor_out[3][17][4] + xor_out[4][17][4];
assign sum_out[1][17][4] = xor_out[5][17][4] + xor_out[6][17][4] + xor_out[7][17][4] + xor_out[8][17][4] + xor_out[9][17][4];
assign sum_out[2][17][4] = xor_out[10][17][4] + xor_out[11][17][4] + xor_out[12][17][4] + xor_out[13][17][4] + xor_out[14][17][4];
assign sum_out[3][17][4] = xor_out[15][17][4] + xor_out[16][17][4] + xor_out[17][17][4] + xor_out[18][17][4] + xor_out[19][17][4];
assign sum_out[4][17][4] = xor_out[20][17][4] + xor_out[21][17][4] + xor_out[22][17][4] + xor_out[23][17][4] + xor_out[24][17][4];
assign sum_out[5][17][4] = xor_out[25][17][4] + xor_out[26][17][4] + xor_out[27][17][4] + xor_out[28][17][4] + xor_out[29][17][4];
assign sum_out[6][17][4] = xor_out[30][17][4] + xor_out[31][17][4] + xor_out[32][17][4] + xor_out[33][17][4] + xor_out[34][17][4];
assign sum_out[7][17][4] = xor_out[35][17][4] + xor_out[36][17][4] + xor_out[37][17][4] + xor_out[38][17][4] + xor_out[39][17][4];
assign sum_out[8][17][4] = xor_out[40][17][4] + xor_out[41][17][4] + xor_out[42][17][4] + xor_out[43][17][4] + xor_out[44][17][4];
assign sum_out[9][17][4] = xor_out[45][17][4] + xor_out[46][17][4] + xor_out[47][17][4] + xor_out[48][17][4] + xor_out[49][17][4];
assign sum_out[10][17][4] = xor_out[50][17][4] + xor_out[51][17][4] + xor_out[52][17][4] + xor_out[53][17][4] + xor_out[54][17][4];
assign sum_out[11][17][4] = xor_out[55][17][4] + xor_out[56][17][4] + xor_out[57][17][4] + xor_out[58][17][4] + xor_out[59][17][4];
assign sum_out[12][17][4] = xor_out[60][17][4] + xor_out[61][17][4] + xor_out[62][17][4] + xor_out[63][17][4] + xor_out[64][17][4];
assign sum_out[13][17][4] = xor_out[65][17][4] + xor_out[66][17][4] + xor_out[67][17][4] + xor_out[68][17][4] + xor_out[69][17][4];
assign sum_out[14][17][4] = xor_out[70][17][4] + xor_out[71][17][4] + xor_out[72][17][4] + xor_out[73][17][4] + xor_out[74][17][4];
assign sum_out[15][17][4] = xor_out[75][17][4] + xor_out[76][17][4] + xor_out[77][17][4] + xor_out[78][17][4] + xor_out[79][17][4];
assign sum_out[16][17][4] = xor_out[80][17][4] + xor_out[81][17][4] + xor_out[82][17][4] + xor_out[83][17][4] + xor_out[84][17][4];
assign sum_out[17][17][4] = xor_out[85][17][4] + xor_out[86][17][4] + xor_out[87][17][4] + xor_out[88][17][4] + xor_out[89][17][4];
assign sum_out[18][17][4] = xor_out[90][17][4] + xor_out[91][17][4] + xor_out[92][17][4] + xor_out[93][17][4] + xor_out[94][17][4];
assign sum_out[19][17][4] = xor_out[95][17][4] + xor_out[96][17][4] + xor_out[97][17][4] + xor_out[98][17][4] + xor_out[99][17][4];

assign sum_out[0][17][5] = xor_out[0][17][5] + xor_out[1][17][5] + xor_out[2][17][5] + xor_out[3][17][5] + xor_out[4][17][5];
assign sum_out[1][17][5] = xor_out[5][17][5] + xor_out[6][17][5] + xor_out[7][17][5] + xor_out[8][17][5] + xor_out[9][17][5];
assign sum_out[2][17][5] = xor_out[10][17][5] + xor_out[11][17][5] + xor_out[12][17][5] + xor_out[13][17][5] + xor_out[14][17][5];
assign sum_out[3][17][5] = xor_out[15][17][5] + xor_out[16][17][5] + xor_out[17][17][5] + xor_out[18][17][5] + xor_out[19][17][5];
assign sum_out[4][17][5] = xor_out[20][17][5] + xor_out[21][17][5] + xor_out[22][17][5] + xor_out[23][17][5] + xor_out[24][17][5];
assign sum_out[5][17][5] = xor_out[25][17][5] + xor_out[26][17][5] + xor_out[27][17][5] + xor_out[28][17][5] + xor_out[29][17][5];
assign sum_out[6][17][5] = xor_out[30][17][5] + xor_out[31][17][5] + xor_out[32][17][5] + xor_out[33][17][5] + xor_out[34][17][5];
assign sum_out[7][17][5] = xor_out[35][17][5] + xor_out[36][17][5] + xor_out[37][17][5] + xor_out[38][17][5] + xor_out[39][17][5];
assign sum_out[8][17][5] = xor_out[40][17][5] + xor_out[41][17][5] + xor_out[42][17][5] + xor_out[43][17][5] + xor_out[44][17][5];
assign sum_out[9][17][5] = xor_out[45][17][5] + xor_out[46][17][5] + xor_out[47][17][5] + xor_out[48][17][5] + xor_out[49][17][5];
assign sum_out[10][17][5] = xor_out[50][17][5] + xor_out[51][17][5] + xor_out[52][17][5] + xor_out[53][17][5] + xor_out[54][17][5];
assign sum_out[11][17][5] = xor_out[55][17][5] + xor_out[56][17][5] + xor_out[57][17][5] + xor_out[58][17][5] + xor_out[59][17][5];
assign sum_out[12][17][5] = xor_out[60][17][5] + xor_out[61][17][5] + xor_out[62][17][5] + xor_out[63][17][5] + xor_out[64][17][5];
assign sum_out[13][17][5] = xor_out[65][17][5] + xor_out[66][17][5] + xor_out[67][17][5] + xor_out[68][17][5] + xor_out[69][17][5];
assign sum_out[14][17][5] = xor_out[70][17][5] + xor_out[71][17][5] + xor_out[72][17][5] + xor_out[73][17][5] + xor_out[74][17][5];
assign sum_out[15][17][5] = xor_out[75][17][5] + xor_out[76][17][5] + xor_out[77][17][5] + xor_out[78][17][5] + xor_out[79][17][5];
assign sum_out[16][17][5] = xor_out[80][17][5] + xor_out[81][17][5] + xor_out[82][17][5] + xor_out[83][17][5] + xor_out[84][17][5];
assign sum_out[17][17][5] = xor_out[85][17][5] + xor_out[86][17][5] + xor_out[87][17][5] + xor_out[88][17][5] + xor_out[89][17][5];
assign sum_out[18][17][5] = xor_out[90][17][5] + xor_out[91][17][5] + xor_out[92][17][5] + xor_out[93][17][5] + xor_out[94][17][5];
assign sum_out[19][17][5] = xor_out[95][17][5] + xor_out[96][17][5] + xor_out[97][17][5] + xor_out[98][17][5] + xor_out[99][17][5];

assign sum_out[0][17][6] = xor_out[0][17][6] + xor_out[1][17][6] + xor_out[2][17][6] + xor_out[3][17][6] + xor_out[4][17][6];
assign sum_out[1][17][6] = xor_out[5][17][6] + xor_out[6][17][6] + xor_out[7][17][6] + xor_out[8][17][6] + xor_out[9][17][6];
assign sum_out[2][17][6] = xor_out[10][17][6] + xor_out[11][17][6] + xor_out[12][17][6] + xor_out[13][17][6] + xor_out[14][17][6];
assign sum_out[3][17][6] = xor_out[15][17][6] + xor_out[16][17][6] + xor_out[17][17][6] + xor_out[18][17][6] + xor_out[19][17][6];
assign sum_out[4][17][6] = xor_out[20][17][6] + xor_out[21][17][6] + xor_out[22][17][6] + xor_out[23][17][6] + xor_out[24][17][6];
assign sum_out[5][17][6] = xor_out[25][17][6] + xor_out[26][17][6] + xor_out[27][17][6] + xor_out[28][17][6] + xor_out[29][17][6];
assign sum_out[6][17][6] = xor_out[30][17][6] + xor_out[31][17][6] + xor_out[32][17][6] + xor_out[33][17][6] + xor_out[34][17][6];
assign sum_out[7][17][6] = xor_out[35][17][6] + xor_out[36][17][6] + xor_out[37][17][6] + xor_out[38][17][6] + xor_out[39][17][6];
assign sum_out[8][17][6] = xor_out[40][17][6] + xor_out[41][17][6] + xor_out[42][17][6] + xor_out[43][17][6] + xor_out[44][17][6];
assign sum_out[9][17][6] = xor_out[45][17][6] + xor_out[46][17][6] + xor_out[47][17][6] + xor_out[48][17][6] + xor_out[49][17][6];
assign sum_out[10][17][6] = xor_out[50][17][6] + xor_out[51][17][6] + xor_out[52][17][6] + xor_out[53][17][6] + xor_out[54][17][6];
assign sum_out[11][17][6] = xor_out[55][17][6] + xor_out[56][17][6] + xor_out[57][17][6] + xor_out[58][17][6] + xor_out[59][17][6];
assign sum_out[12][17][6] = xor_out[60][17][6] + xor_out[61][17][6] + xor_out[62][17][6] + xor_out[63][17][6] + xor_out[64][17][6];
assign sum_out[13][17][6] = xor_out[65][17][6] + xor_out[66][17][6] + xor_out[67][17][6] + xor_out[68][17][6] + xor_out[69][17][6];
assign sum_out[14][17][6] = xor_out[70][17][6] + xor_out[71][17][6] + xor_out[72][17][6] + xor_out[73][17][6] + xor_out[74][17][6];
assign sum_out[15][17][6] = xor_out[75][17][6] + xor_out[76][17][6] + xor_out[77][17][6] + xor_out[78][17][6] + xor_out[79][17][6];
assign sum_out[16][17][6] = xor_out[80][17][6] + xor_out[81][17][6] + xor_out[82][17][6] + xor_out[83][17][6] + xor_out[84][17][6];
assign sum_out[17][17][6] = xor_out[85][17][6] + xor_out[86][17][6] + xor_out[87][17][6] + xor_out[88][17][6] + xor_out[89][17][6];
assign sum_out[18][17][6] = xor_out[90][17][6] + xor_out[91][17][6] + xor_out[92][17][6] + xor_out[93][17][6] + xor_out[94][17][6];
assign sum_out[19][17][6] = xor_out[95][17][6] + xor_out[96][17][6] + xor_out[97][17][6] + xor_out[98][17][6] + xor_out[99][17][6];

assign sum_out[0][17][7] = xor_out[0][17][7] + xor_out[1][17][7] + xor_out[2][17][7] + xor_out[3][17][7] + xor_out[4][17][7];
assign sum_out[1][17][7] = xor_out[5][17][7] + xor_out[6][17][7] + xor_out[7][17][7] + xor_out[8][17][7] + xor_out[9][17][7];
assign sum_out[2][17][7] = xor_out[10][17][7] + xor_out[11][17][7] + xor_out[12][17][7] + xor_out[13][17][7] + xor_out[14][17][7];
assign sum_out[3][17][7] = xor_out[15][17][7] + xor_out[16][17][7] + xor_out[17][17][7] + xor_out[18][17][7] + xor_out[19][17][7];
assign sum_out[4][17][7] = xor_out[20][17][7] + xor_out[21][17][7] + xor_out[22][17][7] + xor_out[23][17][7] + xor_out[24][17][7];
assign sum_out[5][17][7] = xor_out[25][17][7] + xor_out[26][17][7] + xor_out[27][17][7] + xor_out[28][17][7] + xor_out[29][17][7];
assign sum_out[6][17][7] = xor_out[30][17][7] + xor_out[31][17][7] + xor_out[32][17][7] + xor_out[33][17][7] + xor_out[34][17][7];
assign sum_out[7][17][7] = xor_out[35][17][7] + xor_out[36][17][7] + xor_out[37][17][7] + xor_out[38][17][7] + xor_out[39][17][7];
assign sum_out[8][17][7] = xor_out[40][17][7] + xor_out[41][17][7] + xor_out[42][17][7] + xor_out[43][17][7] + xor_out[44][17][7];
assign sum_out[9][17][7] = xor_out[45][17][7] + xor_out[46][17][7] + xor_out[47][17][7] + xor_out[48][17][7] + xor_out[49][17][7];
assign sum_out[10][17][7] = xor_out[50][17][7] + xor_out[51][17][7] + xor_out[52][17][7] + xor_out[53][17][7] + xor_out[54][17][7];
assign sum_out[11][17][7] = xor_out[55][17][7] + xor_out[56][17][7] + xor_out[57][17][7] + xor_out[58][17][7] + xor_out[59][17][7];
assign sum_out[12][17][7] = xor_out[60][17][7] + xor_out[61][17][7] + xor_out[62][17][7] + xor_out[63][17][7] + xor_out[64][17][7];
assign sum_out[13][17][7] = xor_out[65][17][7] + xor_out[66][17][7] + xor_out[67][17][7] + xor_out[68][17][7] + xor_out[69][17][7];
assign sum_out[14][17][7] = xor_out[70][17][7] + xor_out[71][17][7] + xor_out[72][17][7] + xor_out[73][17][7] + xor_out[74][17][7];
assign sum_out[15][17][7] = xor_out[75][17][7] + xor_out[76][17][7] + xor_out[77][17][7] + xor_out[78][17][7] + xor_out[79][17][7];
assign sum_out[16][17][7] = xor_out[80][17][7] + xor_out[81][17][7] + xor_out[82][17][7] + xor_out[83][17][7] + xor_out[84][17][7];
assign sum_out[17][17][7] = xor_out[85][17][7] + xor_out[86][17][7] + xor_out[87][17][7] + xor_out[88][17][7] + xor_out[89][17][7];
assign sum_out[18][17][7] = xor_out[90][17][7] + xor_out[91][17][7] + xor_out[92][17][7] + xor_out[93][17][7] + xor_out[94][17][7];
assign sum_out[19][17][7] = xor_out[95][17][7] + xor_out[96][17][7] + xor_out[97][17][7] + xor_out[98][17][7] + xor_out[99][17][7];

assign sum_out[0][17][8] = xor_out[0][17][8] + xor_out[1][17][8] + xor_out[2][17][8] + xor_out[3][17][8] + xor_out[4][17][8];
assign sum_out[1][17][8] = xor_out[5][17][8] + xor_out[6][17][8] + xor_out[7][17][8] + xor_out[8][17][8] + xor_out[9][17][8];
assign sum_out[2][17][8] = xor_out[10][17][8] + xor_out[11][17][8] + xor_out[12][17][8] + xor_out[13][17][8] + xor_out[14][17][8];
assign sum_out[3][17][8] = xor_out[15][17][8] + xor_out[16][17][8] + xor_out[17][17][8] + xor_out[18][17][8] + xor_out[19][17][8];
assign sum_out[4][17][8] = xor_out[20][17][8] + xor_out[21][17][8] + xor_out[22][17][8] + xor_out[23][17][8] + xor_out[24][17][8];
assign sum_out[5][17][8] = xor_out[25][17][8] + xor_out[26][17][8] + xor_out[27][17][8] + xor_out[28][17][8] + xor_out[29][17][8];
assign sum_out[6][17][8] = xor_out[30][17][8] + xor_out[31][17][8] + xor_out[32][17][8] + xor_out[33][17][8] + xor_out[34][17][8];
assign sum_out[7][17][8] = xor_out[35][17][8] + xor_out[36][17][8] + xor_out[37][17][8] + xor_out[38][17][8] + xor_out[39][17][8];
assign sum_out[8][17][8] = xor_out[40][17][8] + xor_out[41][17][8] + xor_out[42][17][8] + xor_out[43][17][8] + xor_out[44][17][8];
assign sum_out[9][17][8] = xor_out[45][17][8] + xor_out[46][17][8] + xor_out[47][17][8] + xor_out[48][17][8] + xor_out[49][17][8];
assign sum_out[10][17][8] = xor_out[50][17][8] + xor_out[51][17][8] + xor_out[52][17][8] + xor_out[53][17][8] + xor_out[54][17][8];
assign sum_out[11][17][8] = xor_out[55][17][8] + xor_out[56][17][8] + xor_out[57][17][8] + xor_out[58][17][8] + xor_out[59][17][8];
assign sum_out[12][17][8] = xor_out[60][17][8] + xor_out[61][17][8] + xor_out[62][17][8] + xor_out[63][17][8] + xor_out[64][17][8];
assign sum_out[13][17][8] = xor_out[65][17][8] + xor_out[66][17][8] + xor_out[67][17][8] + xor_out[68][17][8] + xor_out[69][17][8];
assign sum_out[14][17][8] = xor_out[70][17][8] + xor_out[71][17][8] + xor_out[72][17][8] + xor_out[73][17][8] + xor_out[74][17][8];
assign sum_out[15][17][8] = xor_out[75][17][8] + xor_out[76][17][8] + xor_out[77][17][8] + xor_out[78][17][8] + xor_out[79][17][8];
assign sum_out[16][17][8] = xor_out[80][17][8] + xor_out[81][17][8] + xor_out[82][17][8] + xor_out[83][17][8] + xor_out[84][17][8];
assign sum_out[17][17][8] = xor_out[85][17][8] + xor_out[86][17][8] + xor_out[87][17][8] + xor_out[88][17][8] + xor_out[89][17][8];
assign sum_out[18][17][8] = xor_out[90][17][8] + xor_out[91][17][8] + xor_out[92][17][8] + xor_out[93][17][8] + xor_out[94][17][8];
assign sum_out[19][17][8] = xor_out[95][17][8] + xor_out[96][17][8] + xor_out[97][17][8] + xor_out[98][17][8] + xor_out[99][17][8];

assign sum_out[0][17][9] = xor_out[0][17][9] + xor_out[1][17][9] + xor_out[2][17][9] + xor_out[3][17][9] + xor_out[4][17][9];
assign sum_out[1][17][9] = xor_out[5][17][9] + xor_out[6][17][9] + xor_out[7][17][9] + xor_out[8][17][9] + xor_out[9][17][9];
assign sum_out[2][17][9] = xor_out[10][17][9] + xor_out[11][17][9] + xor_out[12][17][9] + xor_out[13][17][9] + xor_out[14][17][9];
assign sum_out[3][17][9] = xor_out[15][17][9] + xor_out[16][17][9] + xor_out[17][17][9] + xor_out[18][17][9] + xor_out[19][17][9];
assign sum_out[4][17][9] = xor_out[20][17][9] + xor_out[21][17][9] + xor_out[22][17][9] + xor_out[23][17][9] + xor_out[24][17][9];
assign sum_out[5][17][9] = xor_out[25][17][9] + xor_out[26][17][9] + xor_out[27][17][9] + xor_out[28][17][9] + xor_out[29][17][9];
assign sum_out[6][17][9] = xor_out[30][17][9] + xor_out[31][17][9] + xor_out[32][17][9] + xor_out[33][17][9] + xor_out[34][17][9];
assign sum_out[7][17][9] = xor_out[35][17][9] + xor_out[36][17][9] + xor_out[37][17][9] + xor_out[38][17][9] + xor_out[39][17][9];
assign sum_out[8][17][9] = xor_out[40][17][9] + xor_out[41][17][9] + xor_out[42][17][9] + xor_out[43][17][9] + xor_out[44][17][9];
assign sum_out[9][17][9] = xor_out[45][17][9] + xor_out[46][17][9] + xor_out[47][17][9] + xor_out[48][17][9] + xor_out[49][17][9];
assign sum_out[10][17][9] = xor_out[50][17][9] + xor_out[51][17][9] + xor_out[52][17][9] + xor_out[53][17][9] + xor_out[54][17][9];
assign sum_out[11][17][9] = xor_out[55][17][9] + xor_out[56][17][9] + xor_out[57][17][9] + xor_out[58][17][9] + xor_out[59][17][9];
assign sum_out[12][17][9] = xor_out[60][17][9] + xor_out[61][17][9] + xor_out[62][17][9] + xor_out[63][17][9] + xor_out[64][17][9];
assign sum_out[13][17][9] = xor_out[65][17][9] + xor_out[66][17][9] + xor_out[67][17][9] + xor_out[68][17][9] + xor_out[69][17][9];
assign sum_out[14][17][9] = xor_out[70][17][9] + xor_out[71][17][9] + xor_out[72][17][9] + xor_out[73][17][9] + xor_out[74][17][9];
assign sum_out[15][17][9] = xor_out[75][17][9] + xor_out[76][17][9] + xor_out[77][17][9] + xor_out[78][17][9] + xor_out[79][17][9];
assign sum_out[16][17][9] = xor_out[80][17][9] + xor_out[81][17][9] + xor_out[82][17][9] + xor_out[83][17][9] + xor_out[84][17][9];
assign sum_out[17][17][9] = xor_out[85][17][9] + xor_out[86][17][9] + xor_out[87][17][9] + xor_out[88][17][9] + xor_out[89][17][9];
assign sum_out[18][17][9] = xor_out[90][17][9] + xor_out[91][17][9] + xor_out[92][17][9] + xor_out[93][17][9] + xor_out[94][17][9];
assign sum_out[19][17][9] = xor_out[95][17][9] + xor_out[96][17][9] + xor_out[97][17][9] + xor_out[98][17][9] + xor_out[99][17][9];

assign sum_out[0][17][10] = xor_out[0][17][10] + xor_out[1][17][10] + xor_out[2][17][10] + xor_out[3][17][10] + xor_out[4][17][10];
assign sum_out[1][17][10] = xor_out[5][17][10] + xor_out[6][17][10] + xor_out[7][17][10] + xor_out[8][17][10] + xor_out[9][17][10];
assign sum_out[2][17][10] = xor_out[10][17][10] + xor_out[11][17][10] + xor_out[12][17][10] + xor_out[13][17][10] + xor_out[14][17][10];
assign sum_out[3][17][10] = xor_out[15][17][10] + xor_out[16][17][10] + xor_out[17][17][10] + xor_out[18][17][10] + xor_out[19][17][10];
assign sum_out[4][17][10] = xor_out[20][17][10] + xor_out[21][17][10] + xor_out[22][17][10] + xor_out[23][17][10] + xor_out[24][17][10];
assign sum_out[5][17][10] = xor_out[25][17][10] + xor_out[26][17][10] + xor_out[27][17][10] + xor_out[28][17][10] + xor_out[29][17][10];
assign sum_out[6][17][10] = xor_out[30][17][10] + xor_out[31][17][10] + xor_out[32][17][10] + xor_out[33][17][10] + xor_out[34][17][10];
assign sum_out[7][17][10] = xor_out[35][17][10] + xor_out[36][17][10] + xor_out[37][17][10] + xor_out[38][17][10] + xor_out[39][17][10];
assign sum_out[8][17][10] = xor_out[40][17][10] + xor_out[41][17][10] + xor_out[42][17][10] + xor_out[43][17][10] + xor_out[44][17][10];
assign sum_out[9][17][10] = xor_out[45][17][10] + xor_out[46][17][10] + xor_out[47][17][10] + xor_out[48][17][10] + xor_out[49][17][10];
assign sum_out[10][17][10] = xor_out[50][17][10] + xor_out[51][17][10] + xor_out[52][17][10] + xor_out[53][17][10] + xor_out[54][17][10];
assign sum_out[11][17][10] = xor_out[55][17][10] + xor_out[56][17][10] + xor_out[57][17][10] + xor_out[58][17][10] + xor_out[59][17][10];
assign sum_out[12][17][10] = xor_out[60][17][10] + xor_out[61][17][10] + xor_out[62][17][10] + xor_out[63][17][10] + xor_out[64][17][10];
assign sum_out[13][17][10] = xor_out[65][17][10] + xor_out[66][17][10] + xor_out[67][17][10] + xor_out[68][17][10] + xor_out[69][17][10];
assign sum_out[14][17][10] = xor_out[70][17][10] + xor_out[71][17][10] + xor_out[72][17][10] + xor_out[73][17][10] + xor_out[74][17][10];
assign sum_out[15][17][10] = xor_out[75][17][10] + xor_out[76][17][10] + xor_out[77][17][10] + xor_out[78][17][10] + xor_out[79][17][10];
assign sum_out[16][17][10] = xor_out[80][17][10] + xor_out[81][17][10] + xor_out[82][17][10] + xor_out[83][17][10] + xor_out[84][17][10];
assign sum_out[17][17][10] = xor_out[85][17][10] + xor_out[86][17][10] + xor_out[87][17][10] + xor_out[88][17][10] + xor_out[89][17][10];
assign sum_out[18][17][10] = xor_out[90][17][10] + xor_out[91][17][10] + xor_out[92][17][10] + xor_out[93][17][10] + xor_out[94][17][10];
assign sum_out[19][17][10] = xor_out[95][17][10] + xor_out[96][17][10] + xor_out[97][17][10] + xor_out[98][17][10] + xor_out[99][17][10];

assign sum_out[0][17][11] = xor_out[0][17][11] + xor_out[1][17][11] + xor_out[2][17][11] + xor_out[3][17][11] + xor_out[4][17][11];
assign sum_out[1][17][11] = xor_out[5][17][11] + xor_out[6][17][11] + xor_out[7][17][11] + xor_out[8][17][11] + xor_out[9][17][11];
assign sum_out[2][17][11] = xor_out[10][17][11] + xor_out[11][17][11] + xor_out[12][17][11] + xor_out[13][17][11] + xor_out[14][17][11];
assign sum_out[3][17][11] = xor_out[15][17][11] + xor_out[16][17][11] + xor_out[17][17][11] + xor_out[18][17][11] + xor_out[19][17][11];
assign sum_out[4][17][11] = xor_out[20][17][11] + xor_out[21][17][11] + xor_out[22][17][11] + xor_out[23][17][11] + xor_out[24][17][11];
assign sum_out[5][17][11] = xor_out[25][17][11] + xor_out[26][17][11] + xor_out[27][17][11] + xor_out[28][17][11] + xor_out[29][17][11];
assign sum_out[6][17][11] = xor_out[30][17][11] + xor_out[31][17][11] + xor_out[32][17][11] + xor_out[33][17][11] + xor_out[34][17][11];
assign sum_out[7][17][11] = xor_out[35][17][11] + xor_out[36][17][11] + xor_out[37][17][11] + xor_out[38][17][11] + xor_out[39][17][11];
assign sum_out[8][17][11] = xor_out[40][17][11] + xor_out[41][17][11] + xor_out[42][17][11] + xor_out[43][17][11] + xor_out[44][17][11];
assign sum_out[9][17][11] = xor_out[45][17][11] + xor_out[46][17][11] + xor_out[47][17][11] + xor_out[48][17][11] + xor_out[49][17][11];
assign sum_out[10][17][11] = xor_out[50][17][11] + xor_out[51][17][11] + xor_out[52][17][11] + xor_out[53][17][11] + xor_out[54][17][11];
assign sum_out[11][17][11] = xor_out[55][17][11] + xor_out[56][17][11] + xor_out[57][17][11] + xor_out[58][17][11] + xor_out[59][17][11];
assign sum_out[12][17][11] = xor_out[60][17][11] + xor_out[61][17][11] + xor_out[62][17][11] + xor_out[63][17][11] + xor_out[64][17][11];
assign sum_out[13][17][11] = xor_out[65][17][11] + xor_out[66][17][11] + xor_out[67][17][11] + xor_out[68][17][11] + xor_out[69][17][11];
assign sum_out[14][17][11] = xor_out[70][17][11] + xor_out[71][17][11] + xor_out[72][17][11] + xor_out[73][17][11] + xor_out[74][17][11];
assign sum_out[15][17][11] = xor_out[75][17][11] + xor_out[76][17][11] + xor_out[77][17][11] + xor_out[78][17][11] + xor_out[79][17][11];
assign sum_out[16][17][11] = xor_out[80][17][11] + xor_out[81][17][11] + xor_out[82][17][11] + xor_out[83][17][11] + xor_out[84][17][11];
assign sum_out[17][17][11] = xor_out[85][17][11] + xor_out[86][17][11] + xor_out[87][17][11] + xor_out[88][17][11] + xor_out[89][17][11];
assign sum_out[18][17][11] = xor_out[90][17][11] + xor_out[91][17][11] + xor_out[92][17][11] + xor_out[93][17][11] + xor_out[94][17][11];
assign sum_out[19][17][11] = xor_out[95][17][11] + xor_out[96][17][11] + xor_out[97][17][11] + xor_out[98][17][11] + xor_out[99][17][11];

assign sum_out[0][17][12] = xor_out[0][17][12] + xor_out[1][17][12] + xor_out[2][17][12] + xor_out[3][17][12] + xor_out[4][17][12];
assign sum_out[1][17][12] = xor_out[5][17][12] + xor_out[6][17][12] + xor_out[7][17][12] + xor_out[8][17][12] + xor_out[9][17][12];
assign sum_out[2][17][12] = xor_out[10][17][12] + xor_out[11][17][12] + xor_out[12][17][12] + xor_out[13][17][12] + xor_out[14][17][12];
assign sum_out[3][17][12] = xor_out[15][17][12] + xor_out[16][17][12] + xor_out[17][17][12] + xor_out[18][17][12] + xor_out[19][17][12];
assign sum_out[4][17][12] = xor_out[20][17][12] + xor_out[21][17][12] + xor_out[22][17][12] + xor_out[23][17][12] + xor_out[24][17][12];
assign sum_out[5][17][12] = xor_out[25][17][12] + xor_out[26][17][12] + xor_out[27][17][12] + xor_out[28][17][12] + xor_out[29][17][12];
assign sum_out[6][17][12] = xor_out[30][17][12] + xor_out[31][17][12] + xor_out[32][17][12] + xor_out[33][17][12] + xor_out[34][17][12];
assign sum_out[7][17][12] = xor_out[35][17][12] + xor_out[36][17][12] + xor_out[37][17][12] + xor_out[38][17][12] + xor_out[39][17][12];
assign sum_out[8][17][12] = xor_out[40][17][12] + xor_out[41][17][12] + xor_out[42][17][12] + xor_out[43][17][12] + xor_out[44][17][12];
assign sum_out[9][17][12] = xor_out[45][17][12] + xor_out[46][17][12] + xor_out[47][17][12] + xor_out[48][17][12] + xor_out[49][17][12];
assign sum_out[10][17][12] = xor_out[50][17][12] + xor_out[51][17][12] + xor_out[52][17][12] + xor_out[53][17][12] + xor_out[54][17][12];
assign sum_out[11][17][12] = xor_out[55][17][12] + xor_out[56][17][12] + xor_out[57][17][12] + xor_out[58][17][12] + xor_out[59][17][12];
assign sum_out[12][17][12] = xor_out[60][17][12] + xor_out[61][17][12] + xor_out[62][17][12] + xor_out[63][17][12] + xor_out[64][17][12];
assign sum_out[13][17][12] = xor_out[65][17][12] + xor_out[66][17][12] + xor_out[67][17][12] + xor_out[68][17][12] + xor_out[69][17][12];
assign sum_out[14][17][12] = xor_out[70][17][12] + xor_out[71][17][12] + xor_out[72][17][12] + xor_out[73][17][12] + xor_out[74][17][12];
assign sum_out[15][17][12] = xor_out[75][17][12] + xor_out[76][17][12] + xor_out[77][17][12] + xor_out[78][17][12] + xor_out[79][17][12];
assign sum_out[16][17][12] = xor_out[80][17][12] + xor_out[81][17][12] + xor_out[82][17][12] + xor_out[83][17][12] + xor_out[84][17][12];
assign sum_out[17][17][12] = xor_out[85][17][12] + xor_out[86][17][12] + xor_out[87][17][12] + xor_out[88][17][12] + xor_out[89][17][12];
assign sum_out[18][17][12] = xor_out[90][17][12] + xor_out[91][17][12] + xor_out[92][17][12] + xor_out[93][17][12] + xor_out[94][17][12];
assign sum_out[19][17][12] = xor_out[95][17][12] + xor_out[96][17][12] + xor_out[97][17][12] + xor_out[98][17][12] + xor_out[99][17][12];

assign sum_out[0][17][13] = xor_out[0][17][13] + xor_out[1][17][13] + xor_out[2][17][13] + xor_out[3][17][13] + xor_out[4][17][13];
assign sum_out[1][17][13] = xor_out[5][17][13] + xor_out[6][17][13] + xor_out[7][17][13] + xor_out[8][17][13] + xor_out[9][17][13];
assign sum_out[2][17][13] = xor_out[10][17][13] + xor_out[11][17][13] + xor_out[12][17][13] + xor_out[13][17][13] + xor_out[14][17][13];
assign sum_out[3][17][13] = xor_out[15][17][13] + xor_out[16][17][13] + xor_out[17][17][13] + xor_out[18][17][13] + xor_out[19][17][13];
assign sum_out[4][17][13] = xor_out[20][17][13] + xor_out[21][17][13] + xor_out[22][17][13] + xor_out[23][17][13] + xor_out[24][17][13];
assign sum_out[5][17][13] = xor_out[25][17][13] + xor_out[26][17][13] + xor_out[27][17][13] + xor_out[28][17][13] + xor_out[29][17][13];
assign sum_out[6][17][13] = xor_out[30][17][13] + xor_out[31][17][13] + xor_out[32][17][13] + xor_out[33][17][13] + xor_out[34][17][13];
assign sum_out[7][17][13] = xor_out[35][17][13] + xor_out[36][17][13] + xor_out[37][17][13] + xor_out[38][17][13] + xor_out[39][17][13];
assign sum_out[8][17][13] = xor_out[40][17][13] + xor_out[41][17][13] + xor_out[42][17][13] + xor_out[43][17][13] + xor_out[44][17][13];
assign sum_out[9][17][13] = xor_out[45][17][13] + xor_out[46][17][13] + xor_out[47][17][13] + xor_out[48][17][13] + xor_out[49][17][13];
assign sum_out[10][17][13] = xor_out[50][17][13] + xor_out[51][17][13] + xor_out[52][17][13] + xor_out[53][17][13] + xor_out[54][17][13];
assign sum_out[11][17][13] = xor_out[55][17][13] + xor_out[56][17][13] + xor_out[57][17][13] + xor_out[58][17][13] + xor_out[59][17][13];
assign sum_out[12][17][13] = xor_out[60][17][13] + xor_out[61][17][13] + xor_out[62][17][13] + xor_out[63][17][13] + xor_out[64][17][13];
assign sum_out[13][17][13] = xor_out[65][17][13] + xor_out[66][17][13] + xor_out[67][17][13] + xor_out[68][17][13] + xor_out[69][17][13];
assign sum_out[14][17][13] = xor_out[70][17][13] + xor_out[71][17][13] + xor_out[72][17][13] + xor_out[73][17][13] + xor_out[74][17][13];
assign sum_out[15][17][13] = xor_out[75][17][13] + xor_out[76][17][13] + xor_out[77][17][13] + xor_out[78][17][13] + xor_out[79][17][13];
assign sum_out[16][17][13] = xor_out[80][17][13] + xor_out[81][17][13] + xor_out[82][17][13] + xor_out[83][17][13] + xor_out[84][17][13];
assign sum_out[17][17][13] = xor_out[85][17][13] + xor_out[86][17][13] + xor_out[87][17][13] + xor_out[88][17][13] + xor_out[89][17][13];
assign sum_out[18][17][13] = xor_out[90][17][13] + xor_out[91][17][13] + xor_out[92][17][13] + xor_out[93][17][13] + xor_out[94][17][13];
assign sum_out[19][17][13] = xor_out[95][17][13] + xor_out[96][17][13] + xor_out[97][17][13] + xor_out[98][17][13] + xor_out[99][17][13];

assign sum_out[0][17][14] = xor_out[0][17][14] + xor_out[1][17][14] + xor_out[2][17][14] + xor_out[3][17][14] + xor_out[4][17][14];
assign sum_out[1][17][14] = xor_out[5][17][14] + xor_out[6][17][14] + xor_out[7][17][14] + xor_out[8][17][14] + xor_out[9][17][14];
assign sum_out[2][17][14] = xor_out[10][17][14] + xor_out[11][17][14] + xor_out[12][17][14] + xor_out[13][17][14] + xor_out[14][17][14];
assign sum_out[3][17][14] = xor_out[15][17][14] + xor_out[16][17][14] + xor_out[17][17][14] + xor_out[18][17][14] + xor_out[19][17][14];
assign sum_out[4][17][14] = xor_out[20][17][14] + xor_out[21][17][14] + xor_out[22][17][14] + xor_out[23][17][14] + xor_out[24][17][14];
assign sum_out[5][17][14] = xor_out[25][17][14] + xor_out[26][17][14] + xor_out[27][17][14] + xor_out[28][17][14] + xor_out[29][17][14];
assign sum_out[6][17][14] = xor_out[30][17][14] + xor_out[31][17][14] + xor_out[32][17][14] + xor_out[33][17][14] + xor_out[34][17][14];
assign sum_out[7][17][14] = xor_out[35][17][14] + xor_out[36][17][14] + xor_out[37][17][14] + xor_out[38][17][14] + xor_out[39][17][14];
assign sum_out[8][17][14] = xor_out[40][17][14] + xor_out[41][17][14] + xor_out[42][17][14] + xor_out[43][17][14] + xor_out[44][17][14];
assign sum_out[9][17][14] = xor_out[45][17][14] + xor_out[46][17][14] + xor_out[47][17][14] + xor_out[48][17][14] + xor_out[49][17][14];
assign sum_out[10][17][14] = xor_out[50][17][14] + xor_out[51][17][14] + xor_out[52][17][14] + xor_out[53][17][14] + xor_out[54][17][14];
assign sum_out[11][17][14] = xor_out[55][17][14] + xor_out[56][17][14] + xor_out[57][17][14] + xor_out[58][17][14] + xor_out[59][17][14];
assign sum_out[12][17][14] = xor_out[60][17][14] + xor_out[61][17][14] + xor_out[62][17][14] + xor_out[63][17][14] + xor_out[64][17][14];
assign sum_out[13][17][14] = xor_out[65][17][14] + xor_out[66][17][14] + xor_out[67][17][14] + xor_out[68][17][14] + xor_out[69][17][14];
assign sum_out[14][17][14] = xor_out[70][17][14] + xor_out[71][17][14] + xor_out[72][17][14] + xor_out[73][17][14] + xor_out[74][17][14];
assign sum_out[15][17][14] = xor_out[75][17][14] + xor_out[76][17][14] + xor_out[77][17][14] + xor_out[78][17][14] + xor_out[79][17][14];
assign sum_out[16][17][14] = xor_out[80][17][14] + xor_out[81][17][14] + xor_out[82][17][14] + xor_out[83][17][14] + xor_out[84][17][14];
assign sum_out[17][17][14] = xor_out[85][17][14] + xor_out[86][17][14] + xor_out[87][17][14] + xor_out[88][17][14] + xor_out[89][17][14];
assign sum_out[18][17][14] = xor_out[90][17][14] + xor_out[91][17][14] + xor_out[92][17][14] + xor_out[93][17][14] + xor_out[94][17][14];
assign sum_out[19][17][14] = xor_out[95][17][14] + xor_out[96][17][14] + xor_out[97][17][14] + xor_out[98][17][14] + xor_out[99][17][14];

assign sum_out[0][17][15] = xor_out[0][17][15] + xor_out[1][17][15] + xor_out[2][17][15] + xor_out[3][17][15] + xor_out[4][17][15];
assign sum_out[1][17][15] = xor_out[5][17][15] + xor_out[6][17][15] + xor_out[7][17][15] + xor_out[8][17][15] + xor_out[9][17][15];
assign sum_out[2][17][15] = xor_out[10][17][15] + xor_out[11][17][15] + xor_out[12][17][15] + xor_out[13][17][15] + xor_out[14][17][15];
assign sum_out[3][17][15] = xor_out[15][17][15] + xor_out[16][17][15] + xor_out[17][17][15] + xor_out[18][17][15] + xor_out[19][17][15];
assign sum_out[4][17][15] = xor_out[20][17][15] + xor_out[21][17][15] + xor_out[22][17][15] + xor_out[23][17][15] + xor_out[24][17][15];
assign sum_out[5][17][15] = xor_out[25][17][15] + xor_out[26][17][15] + xor_out[27][17][15] + xor_out[28][17][15] + xor_out[29][17][15];
assign sum_out[6][17][15] = xor_out[30][17][15] + xor_out[31][17][15] + xor_out[32][17][15] + xor_out[33][17][15] + xor_out[34][17][15];
assign sum_out[7][17][15] = xor_out[35][17][15] + xor_out[36][17][15] + xor_out[37][17][15] + xor_out[38][17][15] + xor_out[39][17][15];
assign sum_out[8][17][15] = xor_out[40][17][15] + xor_out[41][17][15] + xor_out[42][17][15] + xor_out[43][17][15] + xor_out[44][17][15];
assign sum_out[9][17][15] = xor_out[45][17][15] + xor_out[46][17][15] + xor_out[47][17][15] + xor_out[48][17][15] + xor_out[49][17][15];
assign sum_out[10][17][15] = xor_out[50][17][15] + xor_out[51][17][15] + xor_out[52][17][15] + xor_out[53][17][15] + xor_out[54][17][15];
assign sum_out[11][17][15] = xor_out[55][17][15] + xor_out[56][17][15] + xor_out[57][17][15] + xor_out[58][17][15] + xor_out[59][17][15];
assign sum_out[12][17][15] = xor_out[60][17][15] + xor_out[61][17][15] + xor_out[62][17][15] + xor_out[63][17][15] + xor_out[64][17][15];
assign sum_out[13][17][15] = xor_out[65][17][15] + xor_out[66][17][15] + xor_out[67][17][15] + xor_out[68][17][15] + xor_out[69][17][15];
assign sum_out[14][17][15] = xor_out[70][17][15] + xor_out[71][17][15] + xor_out[72][17][15] + xor_out[73][17][15] + xor_out[74][17][15];
assign sum_out[15][17][15] = xor_out[75][17][15] + xor_out[76][17][15] + xor_out[77][17][15] + xor_out[78][17][15] + xor_out[79][17][15];
assign sum_out[16][17][15] = xor_out[80][17][15] + xor_out[81][17][15] + xor_out[82][17][15] + xor_out[83][17][15] + xor_out[84][17][15];
assign sum_out[17][17][15] = xor_out[85][17][15] + xor_out[86][17][15] + xor_out[87][17][15] + xor_out[88][17][15] + xor_out[89][17][15];
assign sum_out[18][17][15] = xor_out[90][17][15] + xor_out[91][17][15] + xor_out[92][17][15] + xor_out[93][17][15] + xor_out[94][17][15];
assign sum_out[19][17][15] = xor_out[95][17][15] + xor_out[96][17][15] + xor_out[97][17][15] + xor_out[98][17][15] + xor_out[99][17][15];

assign sum_out[0][17][16] = xor_out[0][17][16] + xor_out[1][17][16] + xor_out[2][17][16] + xor_out[3][17][16] + xor_out[4][17][16];
assign sum_out[1][17][16] = xor_out[5][17][16] + xor_out[6][17][16] + xor_out[7][17][16] + xor_out[8][17][16] + xor_out[9][17][16];
assign sum_out[2][17][16] = xor_out[10][17][16] + xor_out[11][17][16] + xor_out[12][17][16] + xor_out[13][17][16] + xor_out[14][17][16];
assign sum_out[3][17][16] = xor_out[15][17][16] + xor_out[16][17][16] + xor_out[17][17][16] + xor_out[18][17][16] + xor_out[19][17][16];
assign sum_out[4][17][16] = xor_out[20][17][16] + xor_out[21][17][16] + xor_out[22][17][16] + xor_out[23][17][16] + xor_out[24][17][16];
assign sum_out[5][17][16] = xor_out[25][17][16] + xor_out[26][17][16] + xor_out[27][17][16] + xor_out[28][17][16] + xor_out[29][17][16];
assign sum_out[6][17][16] = xor_out[30][17][16] + xor_out[31][17][16] + xor_out[32][17][16] + xor_out[33][17][16] + xor_out[34][17][16];
assign sum_out[7][17][16] = xor_out[35][17][16] + xor_out[36][17][16] + xor_out[37][17][16] + xor_out[38][17][16] + xor_out[39][17][16];
assign sum_out[8][17][16] = xor_out[40][17][16] + xor_out[41][17][16] + xor_out[42][17][16] + xor_out[43][17][16] + xor_out[44][17][16];
assign sum_out[9][17][16] = xor_out[45][17][16] + xor_out[46][17][16] + xor_out[47][17][16] + xor_out[48][17][16] + xor_out[49][17][16];
assign sum_out[10][17][16] = xor_out[50][17][16] + xor_out[51][17][16] + xor_out[52][17][16] + xor_out[53][17][16] + xor_out[54][17][16];
assign sum_out[11][17][16] = xor_out[55][17][16] + xor_out[56][17][16] + xor_out[57][17][16] + xor_out[58][17][16] + xor_out[59][17][16];
assign sum_out[12][17][16] = xor_out[60][17][16] + xor_out[61][17][16] + xor_out[62][17][16] + xor_out[63][17][16] + xor_out[64][17][16];
assign sum_out[13][17][16] = xor_out[65][17][16] + xor_out[66][17][16] + xor_out[67][17][16] + xor_out[68][17][16] + xor_out[69][17][16];
assign sum_out[14][17][16] = xor_out[70][17][16] + xor_out[71][17][16] + xor_out[72][17][16] + xor_out[73][17][16] + xor_out[74][17][16];
assign sum_out[15][17][16] = xor_out[75][17][16] + xor_out[76][17][16] + xor_out[77][17][16] + xor_out[78][17][16] + xor_out[79][17][16];
assign sum_out[16][17][16] = xor_out[80][17][16] + xor_out[81][17][16] + xor_out[82][17][16] + xor_out[83][17][16] + xor_out[84][17][16];
assign sum_out[17][17][16] = xor_out[85][17][16] + xor_out[86][17][16] + xor_out[87][17][16] + xor_out[88][17][16] + xor_out[89][17][16];
assign sum_out[18][17][16] = xor_out[90][17][16] + xor_out[91][17][16] + xor_out[92][17][16] + xor_out[93][17][16] + xor_out[94][17][16];
assign sum_out[19][17][16] = xor_out[95][17][16] + xor_out[96][17][16] + xor_out[97][17][16] + xor_out[98][17][16] + xor_out[99][17][16];

assign sum_out[0][17][17] = xor_out[0][17][17] + xor_out[1][17][17] + xor_out[2][17][17] + xor_out[3][17][17] + xor_out[4][17][17];
assign sum_out[1][17][17] = xor_out[5][17][17] + xor_out[6][17][17] + xor_out[7][17][17] + xor_out[8][17][17] + xor_out[9][17][17];
assign sum_out[2][17][17] = xor_out[10][17][17] + xor_out[11][17][17] + xor_out[12][17][17] + xor_out[13][17][17] + xor_out[14][17][17];
assign sum_out[3][17][17] = xor_out[15][17][17] + xor_out[16][17][17] + xor_out[17][17][17] + xor_out[18][17][17] + xor_out[19][17][17];
assign sum_out[4][17][17] = xor_out[20][17][17] + xor_out[21][17][17] + xor_out[22][17][17] + xor_out[23][17][17] + xor_out[24][17][17];
assign sum_out[5][17][17] = xor_out[25][17][17] + xor_out[26][17][17] + xor_out[27][17][17] + xor_out[28][17][17] + xor_out[29][17][17];
assign sum_out[6][17][17] = xor_out[30][17][17] + xor_out[31][17][17] + xor_out[32][17][17] + xor_out[33][17][17] + xor_out[34][17][17];
assign sum_out[7][17][17] = xor_out[35][17][17] + xor_out[36][17][17] + xor_out[37][17][17] + xor_out[38][17][17] + xor_out[39][17][17];
assign sum_out[8][17][17] = xor_out[40][17][17] + xor_out[41][17][17] + xor_out[42][17][17] + xor_out[43][17][17] + xor_out[44][17][17];
assign sum_out[9][17][17] = xor_out[45][17][17] + xor_out[46][17][17] + xor_out[47][17][17] + xor_out[48][17][17] + xor_out[49][17][17];
assign sum_out[10][17][17] = xor_out[50][17][17] + xor_out[51][17][17] + xor_out[52][17][17] + xor_out[53][17][17] + xor_out[54][17][17];
assign sum_out[11][17][17] = xor_out[55][17][17] + xor_out[56][17][17] + xor_out[57][17][17] + xor_out[58][17][17] + xor_out[59][17][17];
assign sum_out[12][17][17] = xor_out[60][17][17] + xor_out[61][17][17] + xor_out[62][17][17] + xor_out[63][17][17] + xor_out[64][17][17];
assign sum_out[13][17][17] = xor_out[65][17][17] + xor_out[66][17][17] + xor_out[67][17][17] + xor_out[68][17][17] + xor_out[69][17][17];
assign sum_out[14][17][17] = xor_out[70][17][17] + xor_out[71][17][17] + xor_out[72][17][17] + xor_out[73][17][17] + xor_out[74][17][17];
assign sum_out[15][17][17] = xor_out[75][17][17] + xor_out[76][17][17] + xor_out[77][17][17] + xor_out[78][17][17] + xor_out[79][17][17];
assign sum_out[16][17][17] = xor_out[80][17][17] + xor_out[81][17][17] + xor_out[82][17][17] + xor_out[83][17][17] + xor_out[84][17][17];
assign sum_out[17][17][17] = xor_out[85][17][17] + xor_out[86][17][17] + xor_out[87][17][17] + xor_out[88][17][17] + xor_out[89][17][17];
assign sum_out[18][17][17] = xor_out[90][17][17] + xor_out[91][17][17] + xor_out[92][17][17] + xor_out[93][17][17] + xor_out[94][17][17];
assign sum_out[19][17][17] = xor_out[95][17][17] + xor_out[96][17][17] + xor_out[97][17][17] + xor_out[98][17][17] + xor_out[99][17][17];

assign sum_out[0][17][18] = xor_out[0][17][18] + xor_out[1][17][18] + xor_out[2][17][18] + xor_out[3][17][18] + xor_out[4][17][18];
assign sum_out[1][17][18] = xor_out[5][17][18] + xor_out[6][17][18] + xor_out[7][17][18] + xor_out[8][17][18] + xor_out[9][17][18];
assign sum_out[2][17][18] = xor_out[10][17][18] + xor_out[11][17][18] + xor_out[12][17][18] + xor_out[13][17][18] + xor_out[14][17][18];
assign sum_out[3][17][18] = xor_out[15][17][18] + xor_out[16][17][18] + xor_out[17][17][18] + xor_out[18][17][18] + xor_out[19][17][18];
assign sum_out[4][17][18] = xor_out[20][17][18] + xor_out[21][17][18] + xor_out[22][17][18] + xor_out[23][17][18] + xor_out[24][17][18];
assign sum_out[5][17][18] = xor_out[25][17][18] + xor_out[26][17][18] + xor_out[27][17][18] + xor_out[28][17][18] + xor_out[29][17][18];
assign sum_out[6][17][18] = xor_out[30][17][18] + xor_out[31][17][18] + xor_out[32][17][18] + xor_out[33][17][18] + xor_out[34][17][18];
assign sum_out[7][17][18] = xor_out[35][17][18] + xor_out[36][17][18] + xor_out[37][17][18] + xor_out[38][17][18] + xor_out[39][17][18];
assign sum_out[8][17][18] = xor_out[40][17][18] + xor_out[41][17][18] + xor_out[42][17][18] + xor_out[43][17][18] + xor_out[44][17][18];
assign sum_out[9][17][18] = xor_out[45][17][18] + xor_out[46][17][18] + xor_out[47][17][18] + xor_out[48][17][18] + xor_out[49][17][18];
assign sum_out[10][17][18] = xor_out[50][17][18] + xor_out[51][17][18] + xor_out[52][17][18] + xor_out[53][17][18] + xor_out[54][17][18];
assign sum_out[11][17][18] = xor_out[55][17][18] + xor_out[56][17][18] + xor_out[57][17][18] + xor_out[58][17][18] + xor_out[59][17][18];
assign sum_out[12][17][18] = xor_out[60][17][18] + xor_out[61][17][18] + xor_out[62][17][18] + xor_out[63][17][18] + xor_out[64][17][18];
assign sum_out[13][17][18] = xor_out[65][17][18] + xor_out[66][17][18] + xor_out[67][17][18] + xor_out[68][17][18] + xor_out[69][17][18];
assign sum_out[14][17][18] = xor_out[70][17][18] + xor_out[71][17][18] + xor_out[72][17][18] + xor_out[73][17][18] + xor_out[74][17][18];
assign sum_out[15][17][18] = xor_out[75][17][18] + xor_out[76][17][18] + xor_out[77][17][18] + xor_out[78][17][18] + xor_out[79][17][18];
assign sum_out[16][17][18] = xor_out[80][17][18] + xor_out[81][17][18] + xor_out[82][17][18] + xor_out[83][17][18] + xor_out[84][17][18];
assign sum_out[17][17][18] = xor_out[85][17][18] + xor_out[86][17][18] + xor_out[87][17][18] + xor_out[88][17][18] + xor_out[89][17][18];
assign sum_out[18][17][18] = xor_out[90][17][18] + xor_out[91][17][18] + xor_out[92][17][18] + xor_out[93][17][18] + xor_out[94][17][18];
assign sum_out[19][17][18] = xor_out[95][17][18] + xor_out[96][17][18] + xor_out[97][17][18] + xor_out[98][17][18] + xor_out[99][17][18];

assign sum_out[0][17][19] = xor_out[0][17][19] + xor_out[1][17][19] + xor_out[2][17][19] + xor_out[3][17][19] + xor_out[4][17][19];
assign sum_out[1][17][19] = xor_out[5][17][19] + xor_out[6][17][19] + xor_out[7][17][19] + xor_out[8][17][19] + xor_out[9][17][19];
assign sum_out[2][17][19] = xor_out[10][17][19] + xor_out[11][17][19] + xor_out[12][17][19] + xor_out[13][17][19] + xor_out[14][17][19];
assign sum_out[3][17][19] = xor_out[15][17][19] + xor_out[16][17][19] + xor_out[17][17][19] + xor_out[18][17][19] + xor_out[19][17][19];
assign sum_out[4][17][19] = xor_out[20][17][19] + xor_out[21][17][19] + xor_out[22][17][19] + xor_out[23][17][19] + xor_out[24][17][19];
assign sum_out[5][17][19] = xor_out[25][17][19] + xor_out[26][17][19] + xor_out[27][17][19] + xor_out[28][17][19] + xor_out[29][17][19];
assign sum_out[6][17][19] = xor_out[30][17][19] + xor_out[31][17][19] + xor_out[32][17][19] + xor_out[33][17][19] + xor_out[34][17][19];
assign sum_out[7][17][19] = xor_out[35][17][19] + xor_out[36][17][19] + xor_out[37][17][19] + xor_out[38][17][19] + xor_out[39][17][19];
assign sum_out[8][17][19] = xor_out[40][17][19] + xor_out[41][17][19] + xor_out[42][17][19] + xor_out[43][17][19] + xor_out[44][17][19];
assign sum_out[9][17][19] = xor_out[45][17][19] + xor_out[46][17][19] + xor_out[47][17][19] + xor_out[48][17][19] + xor_out[49][17][19];
assign sum_out[10][17][19] = xor_out[50][17][19] + xor_out[51][17][19] + xor_out[52][17][19] + xor_out[53][17][19] + xor_out[54][17][19];
assign sum_out[11][17][19] = xor_out[55][17][19] + xor_out[56][17][19] + xor_out[57][17][19] + xor_out[58][17][19] + xor_out[59][17][19];
assign sum_out[12][17][19] = xor_out[60][17][19] + xor_out[61][17][19] + xor_out[62][17][19] + xor_out[63][17][19] + xor_out[64][17][19];
assign sum_out[13][17][19] = xor_out[65][17][19] + xor_out[66][17][19] + xor_out[67][17][19] + xor_out[68][17][19] + xor_out[69][17][19];
assign sum_out[14][17][19] = xor_out[70][17][19] + xor_out[71][17][19] + xor_out[72][17][19] + xor_out[73][17][19] + xor_out[74][17][19];
assign sum_out[15][17][19] = xor_out[75][17][19] + xor_out[76][17][19] + xor_out[77][17][19] + xor_out[78][17][19] + xor_out[79][17][19];
assign sum_out[16][17][19] = xor_out[80][17][19] + xor_out[81][17][19] + xor_out[82][17][19] + xor_out[83][17][19] + xor_out[84][17][19];
assign sum_out[17][17][19] = xor_out[85][17][19] + xor_out[86][17][19] + xor_out[87][17][19] + xor_out[88][17][19] + xor_out[89][17][19];
assign sum_out[18][17][19] = xor_out[90][17][19] + xor_out[91][17][19] + xor_out[92][17][19] + xor_out[93][17][19] + xor_out[94][17][19];
assign sum_out[19][17][19] = xor_out[95][17][19] + xor_out[96][17][19] + xor_out[97][17][19] + xor_out[98][17][19] + xor_out[99][17][19];

assign sum_out[0][17][20] = xor_out[0][17][20] + xor_out[1][17][20] + xor_out[2][17][20] + xor_out[3][17][20] + xor_out[4][17][20];
assign sum_out[1][17][20] = xor_out[5][17][20] + xor_out[6][17][20] + xor_out[7][17][20] + xor_out[8][17][20] + xor_out[9][17][20];
assign sum_out[2][17][20] = xor_out[10][17][20] + xor_out[11][17][20] + xor_out[12][17][20] + xor_out[13][17][20] + xor_out[14][17][20];
assign sum_out[3][17][20] = xor_out[15][17][20] + xor_out[16][17][20] + xor_out[17][17][20] + xor_out[18][17][20] + xor_out[19][17][20];
assign sum_out[4][17][20] = xor_out[20][17][20] + xor_out[21][17][20] + xor_out[22][17][20] + xor_out[23][17][20] + xor_out[24][17][20];
assign sum_out[5][17][20] = xor_out[25][17][20] + xor_out[26][17][20] + xor_out[27][17][20] + xor_out[28][17][20] + xor_out[29][17][20];
assign sum_out[6][17][20] = xor_out[30][17][20] + xor_out[31][17][20] + xor_out[32][17][20] + xor_out[33][17][20] + xor_out[34][17][20];
assign sum_out[7][17][20] = xor_out[35][17][20] + xor_out[36][17][20] + xor_out[37][17][20] + xor_out[38][17][20] + xor_out[39][17][20];
assign sum_out[8][17][20] = xor_out[40][17][20] + xor_out[41][17][20] + xor_out[42][17][20] + xor_out[43][17][20] + xor_out[44][17][20];
assign sum_out[9][17][20] = xor_out[45][17][20] + xor_out[46][17][20] + xor_out[47][17][20] + xor_out[48][17][20] + xor_out[49][17][20];
assign sum_out[10][17][20] = xor_out[50][17][20] + xor_out[51][17][20] + xor_out[52][17][20] + xor_out[53][17][20] + xor_out[54][17][20];
assign sum_out[11][17][20] = xor_out[55][17][20] + xor_out[56][17][20] + xor_out[57][17][20] + xor_out[58][17][20] + xor_out[59][17][20];
assign sum_out[12][17][20] = xor_out[60][17][20] + xor_out[61][17][20] + xor_out[62][17][20] + xor_out[63][17][20] + xor_out[64][17][20];
assign sum_out[13][17][20] = xor_out[65][17][20] + xor_out[66][17][20] + xor_out[67][17][20] + xor_out[68][17][20] + xor_out[69][17][20];
assign sum_out[14][17][20] = xor_out[70][17][20] + xor_out[71][17][20] + xor_out[72][17][20] + xor_out[73][17][20] + xor_out[74][17][20];
assign sum_out[15][17][20] = xor_out[75][17][20] + xor_out[76][17][20] + xor_out[77][17][20] + xor_out[78][17][20] + xor_out[79][17][20];
assign sum_out[16][17][20] = xor_out[80][17][20] + xor_out[81][17][20] + xor_out[82][17][20] + xor_out[83][17][20] + xor_out[84][17][20];
assign sum_out[17][17][20] = xor_out[85][17][20] + xor_out[86][17][20] + xor_out[87][17][20] + xor_out[88][17][20] + xor_out[89][17][20];
assign sum_out[18][17][20] = xor_out[90][17][20] + xor_out[91][17][20] + xor_out[92][17][20] + xor_out[93][17][20] + xor_out[94][17][20];
assign sum_out[19][17][20] = xor_out[95][17][20] + xor_out[96][17][20] + xor_out[97][17][20] + xor_out[98][17][20] + xor_out[99][17][20];

assign sum_out[0][17][21] = xor_out[0][17][21] + xor_out[1][17][21] + xor_out[2][17][21] + xor_out[3][17][21] + xor_out[4][17][21];
assign sum_out[1][17][21] = xor_out[5][17][21] + xor_out[6][17][21] + xor_out[7][17][21] + xor_out[8][17][21] + xor_out[9][17][21];
assign sum_out[2][17][21] = xor_out[10][17][21] + xor_out[11][17][21] + xor_out[12][17][21] + xor_out[13][17][21] + xor_out[14][17][21];
assign sum_out[3][17][21] = xor_out[15][17][21] + xor_out[16][17][21] + xor_out[17][17][21] + xor_out[18][17][21] + xor_out[19][17][21];
assign sum_out[4][17][21] = xor_out[20][17][21] + xor_out[21][17][21] + xor_out[22][17][21] + xor_out[23][17][21] + xor_out[24][17][21];
assign sum_out[5][17][21] = xor_out[25][17][21] + xor_out[26][17][21] + xor_out[27][17][21] + xor_out[28][17][21] + xor_out[29][17][21];
assign sum_out[6][17][21] = xor_out[30][17][21] + xor_out[31][17][21] + xor_out[32][17][21] + xor_out[33][17][21] + xor_out[34][17][21];
assign sum_out[7][17][21] = xor_out[35][17][21] + xor_out[36][17][21] + xor_out[37][17][21] + xor_out[38][17][21] + xor_out[39][17][21];
assign sum_out[8][17][21] = xor_out[40][17][21] + xor_out[41][17][21] + xor_out[42][17][21] + xor_out[43][17][21] + xor_out[44][17][21];
assign sum_out[9][17][21] = xor_out[45][17][21] + xor_out[46][17][21] + xor_out[47][17][21] + xor_out[48][17][21] + xor_out[49][17][21];
assign sum_out[10][17][21] = xor_out[50][17][21] + xor_out[51][17][21] + xor_out[52][17][21] + xor_out[53][17][21] + xor_out[54][17][21];
assign sum_out[11][17][21] = xor_out[55][17][21] + xor_out[56][17][21] + xor_out[57][17][21] + xor_out[58][17][21] + xor_out[59][17][21];
assign sum_out[12][17][21] = xor_out[60][17][21] + xor_out[61][17][21] + xor_out[62][17][21] + xor_out[63][17][21] + xor_out[64][17][21];
assign sum_out[13][17][21] = xor_out[65][17][21] + xor_out[66][17][21] + xor_out[67][17][21] + xor_out[68][17][21] + xor_out[69][17][21];
assign sum_out[14][17][21] = xor_out[70][17][21] + xor_out[71][17][21] + xor_out[72][17][21] + xor_out[73][17][21] + xor_out[74][17][21];
assign sum_out[15][17][21] = xor_out[75][17][21] + xor_out[76][17][21] + xor_out[77][17][21] + xor_out[78][17][21] + xor_out[79][17][21];
assign sum_out[16][17][21] = xor_out[80][17][21] + xor_out[81][17][21] + xor_out[82][17][21] + xor_out[83][17][21] + xor_out[84][17][21];
assign sum_out[17][17][21] = xor_out[85][17][21] + xor_out[86][17][21] + xor_out[87][17][21] + xor_out[88][17][21] + xor_out[89][17][21];
assign sum_out[18][17][21] = xor_out[90][17][21] + xor_out[91][17][21] + xor_out[92][17][21] + xor_out[93][17][21] + xor_out[94][17][21];
assign sum_out[19][17][21] = xor_out[95][17][21] + xor_out[96][17][21] + xor_out[97][17][21] + xor_out[98][17][21] + xor_out[99][17][21];

assign sum_out[0][17][22] = xor_out[0][17][22] + xor_out[1][17][22] + xor_out[2][17][22] + xor_out[3][17][22] + xor_out[4][17][22];
assign sum_out[1][17][22] = xor_out[5][17][22] + xor_out[6][17][22] + xor_out[7][17][22] + xor_out[8][17][22] + xor_out[9][17][22];
assign sum_out[2][17][22] = xor_out[10][17][22] + xor_out[11][17][22] + xor_out[12][17][22] + xor_out[13][17][22] + xor_out[14][17][22];
assign sum_out[3][17][22] = xor_out[15][17][22] + xor_out[16][17][22] + xor_out[17][17][22] + xor_out[18][17][22] + xor_out[19][17][22];
assign sum_out[4][17][22] = xor_out[20][17][22] + xor_out[21][17][22] + xor_out[22][17][22] + xor_out[23][17][22] + xor_out[24][17][22];
assign sum_out[5][17][22] = xor_out[25][17][22] + xor_out[26][17][22] + xor_out[27][17][22] + xor_out[28][17][22] + xor_out[29][17][22];
assign sum_out[6][17][22] = xor_out[30][17][22] + xor_out[31][17][22] + xor_out[32][17][22] + xor_out[33][17][22] + xor_out[34][17][22];
assign sum_out[7][17][22] = xor_out[35][17][22] + xor_out[36][17][22] + xor_out[37][17][22] + xor_out[38][17][22] + xor_out[39][17][22];
assign sum_out[8][17][22] = xor_out[40][17][22] + xor_out[41][17][22] + xor_out[42][17][22] + xor_out[43][17][22] + xor_out[44][17][22];
assign sum_out[9][17][22] = xor_out[45][17][22] + xor_out[46][17][22] + xor_out[47][17][22] + xor_out[48][17][22] + xor_out[49][17][22];
assign sum_out[10][17][22] = xor_out[50][17][22] + xor_out[51][17][22] + xor_out[52][17][22] + xor_out[53][17][22] + xor_out[54][17][22];
assign sum_out[11][17][22] = xor_out[55][17][22] + xor_out[56][17][22] + xor_out[57][17][22] + xor_out[58][17][22] + xor_out[59][17][22];
assign sum_out[12][17][22] = xor_out[60][17][22] + xor_out[61][17][22] + xor_out[62][17][22] + xor_out[63][17][22] + xor_out[64][17][22];
assign sum_out[13][17][22] = xor_out[65][17][22] + xor_out[66][17][22] + xor_out[67][17][22] + xor_out[68][17][22] + xor_out[69][17][22];
assign sum_out[14][17][22] = xor_out[70][17][22] + xor_out[71][17][22] + xor_out[72][17][22] + xor_out[73][17][22] + xor_out[74][17][22];
assign sum_out[15][17][22] = xor_out[75][17][22] + xor_out[76][17][22] + xor_out[77][17][22] + xor_out[78][17][22] + xor_out[79][17][22];
assign sum_out[16][17][22] = xor_out[80][17][22] + xor_out[81][17][22] + xor_out[82][17][22] + xor_out[83][17][22] + xor_out[84][17][22];
assign sum_out[17][17][22] = xor_out[85][17][22] + xor_out[86][17][22] + xor_out[87][17][22] + xor_out[88][17][22] + xor_out[89][17][22];
assign sum_out[18][17][22] = xor_out[90][17][22] + xor_out[91][17][22] + xor_out[92][17][22] + xor_out[93][17][22] + xor_out[94][17][22];
assign sum_out[19][17][22] = xor_out[95][17][22] + xor_out[96][17][22] + xor_out[97][17][22] + xor_out[98][17][22] + xor_out[99][17][22];

assign sum_out[0][17][23] = xor_out[0][17][23] + xor_out[1][17][23] + xor_out[2][17][23] + xor_out[3][17][23] + xor_out[4][17][23];
assign sum_out[1][17][23] = xor_out[5][17][23] + xor_out[6][17][23] + xor_out[7][17][23] + xor_out[8][17][23] + xor_out[9][17][23];
assign sum_out[2][17][23] = xor_out[10][17][23] + xor_out[11][17][23] + xor_out[12][17][23] + xor_out[13][17][23] + xor_out[14][17][23];
assign sum_out[3][17][23] = xor_out[15][17][23] + xor_out[16][17][23] + xor_out[17][17][23] + xor_out[18][17][23] + xor_out[19][17][23];
assign sum_out[4][17][23] = xor_out[20][17][23] + xor_out[21][17][23] + xor_out[22][17][23] + xor_out[23][17][23] + xor_out[24][17][23];
assign sum_out[5][17][23] = xor_out[25][17][23] + xor_out[26][17][23] + xor_out[27][17][23] + xor_out[28][17][23] + xor_out[29][17][23];
assign sum_out[6][17][23] = xor_out[30][17][23] + xor_out[31][17][23] + xor_out[32][17][23] + xor_out[33][17][23] + xor_out[34][17][23];
assign sum_out[7][17][23] = xor_out[35][17][23] + xor_out[36][17][23] + xor_out[37][17][23] + xor_out[38][17][23] + xor_out[39][17][23];
assign sum_out[8][17][23] = xor_out[40][17][23] + xor_out[41][17][23] + xor_out[42][17][23] + xor_out[43][17][23] + xor_out[44][17][23];
assign sum_out[9][17][23] = xor_out[45][17][23] + xor_out[46][17][23] + xor_out[47][17][23] + xor_out[48][17][23] + xor_out[49][17][23];
assign sum_out[10][17][23] = xor_out[50][17][23] + xor_out[51][17][23] + xor_out[52][17][23] + xor_out[53][17][23] + xor_out[54][17][23];
assign sum_out[11][17][23] = xor_out[55][17][23] + xor_out[56][17][23] + xor_out[57][17][23] + xor_out[58][17][23] + xor_out[59][17][23];
assign sum_out[12][17][23] = xor_out[60][17][23] + xor_out[61][17][23] + xor_out[62][17][23] + xor_out[63][17][23] + xor_out[64][17][23];
assign sum_out[13][17][23] = xor_out[65][17][23] + xor_out[66][17][23] + xor_out[67][17][23] + xor_out[68][17][23] + xor_out[69][17][23];
assign sum_out[14][17][23] = xor_out[70][17][23] + xor_out[71][17][23] + xor_out[72][17][23] + xor_out[73][17][23] + xor_out[74][17][23];
assign sum_out[15][17][23] = xor_out[75][17][23] + xor_out[76][17][23] + xor_out[77][17][23] + xor_out[78][17][23] + xor_out[79][17][23];
assign sum_out[16][17][23] = xor_out[80][17][23] + xor_out[81][17][23] + xor_out[82][17][23] + xor_out[83][17][23] + xor_out[84][17][23];
assign sum_out[17][17][23] = xor_out[85][17][23] + xor_out[86][17][23] + xor_out[87][17][23] + xor_out[88][17][23] + xor_out[89][17][23];
assign sum_out[18][17][23] = xor_out[90][17][23] + xor_out[91][17][23] + xor_out[92][17][23] + xor_out[93][17][23] + xor_out[94][17][23];
assign sum_out[19][17][23] = xor_out[95][17][23] + xor_out[96][17][23] + xor_out[97][17][23] + xor_out[98][17][23] + xor_out[99][17][23];

assign sum_out[0][18][0] = xor_out[0][18][0] + xor_out[1][18][0] + xor_out[2][18][0] + xor_out[3][18][0] + xor_out[4][18][0];
assign sum_out[1][18][0] = xor_out[5][18][0] + xor_out[6][18][0] + xor_out[7][18][0] + xor_out[8][18][0] + xor_out[9][18][0];
assign sum_out[2][18][0] = xor_out[10][18][0] + xor_out[11][18][0] + xor_out[12][18][0] + xor_out[13][18][0] + xor_out[14][18][0];
assign sum_out[3][18][0] = xor_out[15][18][0] + xor_out[16][18][0] + xor_out[17][18][0] + xor_out[18][18][0] + xor_out[19][18][0];
assign sum_out[4][18][0] = xor_out[20][18][0] + xor_out[21][18][0] + xor_out[22][18][0] + xor_out[23][18][0] + xor_out[24][18][0];
assign sum_out[5][18][0] = xor_out[25][18][0] + xor_out[26][18][0] + xor_out[27][18][0] + xor_out[28][18][0] + xor_out[29][18][0];
assign sum_out[6][18][0] = xor_out[30][18][0] + xor_out[31][18][0] + xor_out[32][18][0] + xor_out[33][18][0] + xor_out[34][18][0];
assign sum_out[7][18][0] = xor_out[35][18][0] + xor_out[36][18][0] + xor_out[37][18][0] + xor_out[38][18][0] + xor_out[39][18][0];
assign sum_out[8][18][0] = xor_out[40][18][0] + xor_out[41][18][0] + xor_out[42][18][0] + xor_out[43][18][0] + xor_out[44][18][0];
assign sum_out[9][18][0] = xor_out[45][18][0] + xor_out[46][18][0] + xor_out[47][18][0] + xor_out[48][18][0] + xor_out[49][18][0];
assign sum_out[10][18][0] = xor_out[50][18][0] + xor_out[51][18][0] + xor_out[52][18][0] + xor_out[53][18][0] + xor_out[54][18][0];
assign sum_out[11][18][0] = xor_out[55][18][0] + xor_out[56][18][0] + xor_out[57][18][0] + xor_out[58][18][0] + xor_out[59][18][0];
assign sum_out[12][18][0] = xor_out[60][18][0] + xor_out[61][18][0] + xor_out[62][18][0] + xor_out[63][18][0] + xor_out[64][18][0];
assign sum_out[13][18][0] = xor_out[65][18][0] + xor_out[66][18][0] + xor_out[67][18][0] + xor_out[68][18][0] + xor_out[69][18][0];
assign sum_out[14][18][0] = xor_out[70][18][0] + xor_out[71][18][0] + xor_out[72][18][0] + xor_out[73][18][0] + xor_out[74][18][0];
assign sum_out[15][18][0] = xor_out[75][18][0] + xor_out[76][18][0] + xor_out[77][18][0] + xor_out[78][18][0] + xor_out[79][18][0];
assign sum_out[16][18][0] = xor_out[80][18][0] + xor_out[81][18][0] + xor_out[82][18][0] + xor_out[83][18][0] + xor_out[84][18][0];
assign sum_out[17][18][0] = xor_out[85][18][0] + xor_out[86][18][0] + xor_out[87][18][0] + xor_out[88][18][0] + xor_out[89][18][0];
assign sum_out[18][18][0] = xor_out[90][18][0] + xor_out[91][18][0] + xor_out[92][18][0] + xor_out[93][18][0] + xor_out[94][18][0];
assign sum_out[19][18][0] = xor_out[95][18][0] + xor_out[96][18][0] + xor_out[97][18][0] + xor_out[98][18][0] + xor_out[99][18][0];

assign sum_out[0][18][1] = xor_out[0][18][1] + xor_out[1][18][1] + xor_out[2][18][1] + xor_out[3][18][1] + xor_out[4][18][1];
assign sum_out[1][18][1] = xor_out[5][18][1] + xor_out[6][18][1] + xor_out[7][18][1] + xor_out[8][18][1] + xor_out[9][18][1];
assign sum_out[2][18][1] = xor_out[10][18][1] + xor_out[11][18][1] + xor_out[12][18][1] + xor_out[13][18][1] + xor_out[14][18][1];
assign sum_out[3][18][1] = xor_out[15][18][1] + xor_out[16][18][1] + xor_out[17][18][1] + xor_out[18][18][1] + xor_out[19][18][1];
assign sum_out[4][18][1] = xor_out[20][18][1] + xor_out[21][18][1] + xor_out[22][18][1] + xor_out[23][18][1] + xor_out[24][18][1];
assign sum_out[5][18][1] = xor_out[25][18][1] + xor_out[26][18][1] + xor_out[27][18][1] + xor_out[28][18][1] + xor_out[29][18][1];
assign sum_out[6][18][1] = xor_out[30][18][1] + xor_out[31][18][1] + xor_out[32][18][1] + xor_out[33][18][1] + xor_out[34][18][1];
assign sum_out[7][18][1] = xor_out[35][18][1] + xor_out[36][18][1] + xor_out[37][18][1] + xor_out[38][18][1] + xor_out[39][18][1];
assign sum_out[8][18][1] = xor_out[40][18][1] + xor_out[41][18][1] + xor_out[42][18][1] + xor_out[43][18][1] + xor_out[44][18][1];
assign sum_out[9][18][1] = xor_out[45][18][1] + xor_out[46][18][1] + xor_out[47][18][1] + xor_out[48][18][1] + xor_out[49][18][1];
assign sum_out[10][18][1] = xor_out[50][18][1] + xor_out[51][18][1] + xor_out[52][18][1] + xor_out[53][18][1] + xor_out[54][18][1];
assign sum_out[11][18][1] = xor_out[55][18][1] + xor_out[56][18][1] + xor_out[57][18][1] + xor_out[58][18][1] + xor_out[59][18][1];
assign sum_out[12][18][1] = xor_out[60][18][1] + xor_out[61][18][1] + xor_out[62][18][1] + xor_out[63][18][1] + xor_out[64][18][1];
assign sum_out[13][18][1] = xor_out[65][18][1] + xor_out[66][18][1] + xor_out[67][18][1] + xor_out[68][18][1] + xor_out[69][18][1];
assign sum_out[14][18][1] = xor_out[70][18][1] + xor_out[71][18][1] + xor_out[72][18][1] + xor_out[73][18][1] + xor_out[74][18][1];
assign sum_out[15][18][1] = xor_out[75][18][1] + xor_out[76][18][1] + xor_out[77][18][1] + xor_out[78][18][1] + xor_out[79][18][1];
assign sum_out[16][18][1] = xor_out[80][18][1] + xor_out[81][18][1] + xor_out[82][18][1] + xor_out[83][18][1] + xor_out[84][18][1];
assign sum_out[17][18][1] = xor_out[85][18][1] + xor_out[86][18][1] + xor_out[87][18][1] + xor_out[88][18][1] + xor_out[89][18][1];
assign sum_out[18][18][1] = xor_out[90][18][1] + xor_out[91][18][1] + xor_out[92][18][1] + xor_out[93][18][1] + xor_out[94][18][1];
assign sum_out[19][18][1] = xor_out[95][18][1] + xor_out[96][18][1] + xor_out[97][18][1] + xor_out[98][18][1] + xor_out[99][18][1];

assign sum_out[0][18][2] = xor_out[0][18][2] + xor_out[1][18][2] + xor_out[2][18][2] + xor_out[3][18][2] + xor_out[4][18][2];
assign sum_out[1][18][2] = xor_out[5][18][2] + xor_out[6][18][2] + xor_out[7][18][2] + xor_out[8][18][2] + xor_out[9][18][2];
assign sum_out[2][18][2] = xor_out[10][18][2] + xor_out[11][18][2] + xor_out[12][18][2] + xor_out[13][18][2] + xor_out[14][18][2];
assign sum_out[3][18][2] = xor_out[15][18][2] + xor_out[16][18][2] + xor_out[17][18][2] + xor_out[18][18][2] + xor_out[19][18][2];
assign sum_out[4][18][2] = xor_out[20][18][2] + xor_out[21][18][2] + xor_out[22][18][2] + xor_out[23][18][2] + xor_out[24][18][2];
assign sum_out[5][18][2] = xor_out[25][18][2] + xor_out[26][18][2] + xor_out[27][18][2] + xor_out[28][18][2] + xor_out[29][18][2];
assign sum_out[6][18][2] = xor_out[30][18][2] + xor_out[31][18][2] + xor_out[32][18][2] + xor_out[33][18][2] + xor_out[34][18][2];
assign sum_out[7][18][2] = xor_out[35][18][2] + xor_out[36][18][2] + xor_out[37][18][2] + xor_out[38][18][2] + xor_out[39][18][2];
assign sum_out[8][18][2] = xor_out[40][18][2] + xor_out[41][18][2] + xor_out[42][18][2] + xor_out[43][18][2] + xor_out[44][18][2];
assign sum_out[9][18][2] = xor_out[45][18][2] + xor_out[46][18][2] + xor_out[47][18][2] + xor_out[48][18][2] + xor_out[49][18][2];
assign sum_out[10][18][2] = xor_out[50][18][2] + xor_out[51][18][2] + xor_out[52][18][2] + xor_out[53][18][2] + xor_out[54][18][2];
assign sum_out[11][18][2] = xor_out[55][18][2] + xor_out[56][18][2] + xor_out[57][18][2] + xor_out[58][18][2] + xor_out[59][18][2];
assign sum_out[12][18][2] = xor_out[60][18][2] + xor_out[61][18][2] + xor_out[62][18][2] + xor_out[63][18][2] + xor_out[64][18][2];
assign sum_out[13][18][2] = xor_out[65][18][2] + xor_out[66][18][2] + xor_out[67][18][2] + xor_out[68][18][2] + xor_out[69][18][2];
assign sum_out[14][18][2] = xor_out[70][18][2] + xor_out[71][18][2] + xor_out[72][18][2] + xor_out[73][18][2] + xor_out[74][18][2];
assign sum_out[15][18][2] = xor_out[75][18][2] + xor_out[76][18][2] + xor_out[77][18][2] + xor_out[78][18][2] + xor_out[79][18][2];
assign sum_out[16][18][2] = xor_out[80][18][2] + xor_out[81][18][2] + xor_out[82][18][2] + xor_out[83][18][2] + xor_out[84][18][2];
assign sum_out[17][18][2] = xor_out[85][18][2] + xor_out[86][18][2] + xor_out[87][18][2] + xor_out[88][18][2] + xor_out[89][18][2];
assign sum_out[18][18][2] = xor_out[90][18][2] + xor_out[91][18][2] + xor_out[92][18][2] + xor_out[93][18][2] + xor_out[94][18][2];
assign sum_out[19][18][2] = xor_out[95][18][2] + xor_out[96][18][2] + xor_out[97][18][2] + xor_out[98][18][2] + xor_out[99][18][2];

assign sum_out[0][18][3] = xor_out[0][18][3] + xor_out[1][18][3] + xor_out[2][18][3] + xor_out[3][18][3] + xor_out[4][18][3];
assign sum_out[1][18][3] = xor_out[5][18][3] + xor_out[6][18][3] + xor_out[7][18][3] + xor_out[8][18][3] + xor_out[9][18][3];
assign sum_out[2][18][3] = xor_out[10][18][3] + xor_out[11][18][3] + xor_out[12][18][3] + xor_out[13][18][3] + xor_out[14][18][3];
assign sum_out[3][18][3] = xor_out[15][18][3] + xor_out[16][18][3] + xor_out[17][18][3] + xor_out[18][18][3] + xor_out[19][18][3];
assign sum_out[4][18][3] = xor_out[20][18][3] + xor_out[21][18][3] + xor_out[22][18][3] + xor_out[23][18][3] + xor_out[24][18][3];
assign sum_out[5][18][3] = xor_out[25][18][3] + xor_out[26][18][3] + xor_out[27][18][3] + xor_out[28][18][3] + xor_out[29][18][3];
assign sum_out[6][18][3] = xor_out[30][18][3] + xor_out[31][18][3] + xor_out[32][18][3] + xor_out[33][18][3] + xor_out[34][18][3];
assign sum_out[7][18][3] = xor_out[35][18][3] + xor_out[36][18][3] + xor_out[37][18][3] + xor_out[38][18][3] + xor_out[39][18][3];
assign sum_out[8][18][3] = xor_out[40][18][3] + xor_out[41][18][3] + xor_out[42][18][3] + xor_out[43][18][3] + xor_out[44][18][3];
assign sum_out[9][18][3] = xor_out[45][18][3] + xor_out[46][18][3] + xor_out[47][18][3] + xor_out[48][18][3] + xor_out[49][18][3];
assign sum_out[10][18][3] = xor_out[50][18][3] + xor_out[51][18][3] + xor_out[52][18][3] + xor_out[53][18][3] + xor_out[54][18][3];
assign sum_out[11][18][3] = xor_out[55][18][3] + xor_out[56][18][3] + xor_out[57][18][3] + xor_out[58][18][3] + xor_out[59][18][3];
assign sum_out[12][18][3] = xor_out[60][18][3] + xor_out[61][18][3] + xor_out[62][18][3] + xor_out[63][18][3] + xor_out[64][18][3];
assign sum_out[13][18][3] = xor_out[65][18][3] + xor_out[66][18][3] + xor_out[67][18][3] + xor_out[68][18][3] + xor_out[69][18][3];
assign sum_out[14][18][3] = xor_out[70][18][3] + xor_out[71][18][3] + xor_out[72][18][3] + xor_out[73][18][3] + xor_out[74][18][3];
assign sum_out[15][18][3] = xor_out[75][18][3] + xor_out[76][18][3] + xor_out[77][18][3] + xor_out[78][18][3] + xor_out[79][18][3];
assign sum_out[16][18][3] = xor_out[80][18][3] + xor_out[81][18][3] + xor_out[82][18][3] + xor_out[83][18][3] + xor_out[84][18][3];
assign sum_out[17][18][3] = xor_out[85][18][3] + xor_out[86][18][3] + xor_out[87][18][3] + xor_out[88][18][3] + xor_out[89][18][3];
assign sum_out[18][18][3] = xor_out[90][18][3] + xor_out[91][18][3] + xor_out[92][18][3] + xor_out[93][18][3] + xor_out[94][18][3];
assign sum_out[19][18][3] = xor_out[95][18][3] + xor_out[96][18][3] + xor_out[97][18][3] + xor_out[98][18][3] + xor_out[99][18][3];

assign sum_out[0][18][4] = xor_out[0][18][4] + xor_out[1][18][4] + xor_out[2][18][4] + xor_out[3][18][4] + xor_out[4][18][4];
assign sum_out[1][18][4] = xor_out[5][18][4] + xor_out[6][18][4] + xor_out[7][18][4] + xor_out[8][18][4] + xor_out[9][18][4];
assign sum_out[2][18][4] = xor_out[10][18][4] + xor_out[11][18][4] + xor_out[12][18][4] + xor_out[13][18][4] + xor_out[14][18][4];
assign sum_out[3][18][4] = xor_out[15][18][4] + xor_out[16][18][4] + xor_out[17][18][4] + xor_out[18][18][4] + xor_out[19][18][4];
assign sum_out[4][18][4] = xor_out[20][18][4] + xor_out[21][18][4] + xor_out[22][18][4] + xor_out[23][18][4] + xor_out[24][18][4];
assign sum_out[5][18][4] = xor_out[25][18][4] + xor_out[26][18][4] + xor_out[27][18][4] + xor_out[28][18][4] + xor_out[29][18][4];
assign sum_out[6][18][4] = xor_out[30][18][4] + xor_out[31][18][4] + xor_out[32][18][4] + xor_out[33][18][4] + xor_out[34][18][4];
assign sum_out[7][18][4] = xor_out[35][18][4] + xor_out[36][18][4] + xor_out[37][18][4] + xor_out[38][18][4] + xor_out[39][18][4];
assign sum_out[8][18][4] = xor_out[40][18][4] + xor_out[41][18][4] + xor_out[42][18][4] + xor_out[43][18][4] + xor_out[44][18][4];
assign sum_out[9][18][4] = xor_out[45][18][4] + xor_out[46][18][4] + xor_out[47][18][4] + xor_out[48][18][4] + xor_out[49][18][4];
assign sum_out[10][18][4] = xor_out[50][18][4] + xor_out[51][18][4] + xor_out[52][18][4] + xor_out[53][18][4] + xor_out[54][18][4];
assign sum_out[11][18][4] = xor_out[55][18][4] + xor_out[56][18][4] + xor_out[57][18][4] + xor_out[58][18][4] + xor_out[59][18][4];
assign sum_out[12][18][4] = xor_out[60][18][4] + xor_out[61][18][4] + xor_out[62][18][4] + xor_out[63][18][4] + xor_out[64][18][4];
assign sum_out[13][18][4] = xor_out[65][18][4] + xor_out[66][18][4] + xor_out[67][18][4] + xor_out[68][18][4] + xor_out[69][18][4];
assign sum_out[14][18][4] = xor_out[70][18][4] + xor_out[71][18][4] + xor_out[72][18][4] + xor_out[73][18][4] + xor_out[74][18][4];
assign sum_out[15][18][4] = xor_out[75][18][4] + xor_out[76][18][4] + xor_out[77][18][4] + xor_out[78][18][4] + xor_out[79][18][4];
assign sum_out[16][18][4] = xor_out[80][18][4] + xor_out[81][18][4] + xor_out[82][18][4] + xor_out[83][18][4] + xor_out[84][18][4];
assign sum_out[17][18][4] = xor_out[85][18][4] + xor_out[86][18][4] + xor_out[87][18][4] + xor_out[88][18][4] + xor_out[89][18][4];
assign sum_out[18][18][4] = xor_out[90][18][4] + xor_out[91][18][4] + xor_out[92][18][4] + xor_out[93][18][4] + xor_out[94][18][4];
assign sum_out[19][18][4] = xor_out[95][18][4] + xor_out[96][18][4] + xor_out[97][18][4] + xor_out[98][18][4] + xor_out[99][18][4];

assign sum_out[0][18][5] = xor_out[0][18][5] + xor_out[1][18][5] + xor_out[2][18][5] + xor_out[3][18][5] + xor_out[4][18][5];
assign sum_out[1][18][5] = xor_out[5][18][5] + xor_out[6][18][5] + xor_out[7][18][5] + xor_out[8][18][5] + xor_out[9][18][5];
assign sum_out[2][18][5] = xor_out[10][18][5] + xor_out[11][18][5] + xor_out[12][18][5] + xor_out[13][18][5] + xor_out[14][18][5];
assign sum_out[3][18][5] = xor_out[15][18][5] + xor_out[16][18][5] + xor_out[17][18][5] + xor_out[18][18][5] + xor_out[19][18][5];
assign sum_out[4][18][5] = xor_out[20][18][5] + xor_out[21][18][5] + xor_out[22][18][5] + xor_out[23][18][5] + xor_out[24][18][5];
assign sum_out[5][18][5] = xor_out[25][18][5] + xor_out[26][18][5] + xor_out[27][18][5] + xor_out[28][18][5] + xor_out[29][18][5];
assign sum_out[6][18][5] = xor_out[30][18][5] + xor_out[31][18][5] + xor_out[32][18][5] + xor_out[33][18][5] + xor_out[34][18][5];
assign sum_out[7][18][5] = xor_out[35][18][5] + xor_out[36][18][5] + xor_out[37][18][5] + xor_out[38][18][5] + xor_out[39][18][5];
assign sum_out[8][18][5] = xor_out[40][18][5] + xor_out[41][18][5] + xor_out[42][18][5] + xor_out[43][18][5] + xor_out[44][18][5];
assign sum_out[9][18][5] = xor_out[45][18][5] + xor_out[46][18][5] + xor_out[47][18][5] + xor_out[48][18][5] + xor_out[49][18][5];
assign sum_out[10][18][5] = xor_out[50][18][5] + xor_out[51][18][5] + xor_out[52][18][5] + xor_out[53][18][5] + xor_out[54][18][5];
assign sum_out[11][18][5] = xor_out[55][18][5] + xor_out[56][18][5] + xor_out[57][18][5] + xor_out[58][18][5] + xor_out[59][18][5];
assign sum_out[12][18][5] = xor_out[60][18][5] + xor_out[61][18][5] + xor_out[62][18][5] + xor_out[63][18][5] + xor_out[64][18][5];
assign sum_out[13][18][5] = xor_out[65][18][5] + xor_out[66][18][5] + xor_out[67][18][5] + xor_out[68][18][5] + xor_out[69][18][5];
assign sum_out[14][18][5] = xor_out[70][18][5] + xor_out[71][18][5] + xor_out[72][18][5] + xor_out[73][18][5] + xor_out[74][18][5];
assign sum_out[15][18][5] = xor_out[75][18][5] + xor_out[76][18][5] + xor_out[77][18][5] + xor_out[78][18][5] + xor_out[79][18][5];
assign sum_out[16][18][5] = xor_out[80][18][5] + xor_out[81][18][5] + xor_out[82][18][5] + xor_out[83][18][5] + xor_out[84][18][5];
assign sum_out[17][18][5] = xor_out[85][18][5] + xor_out[86][18][5] + xor_out[87][18][5] + xor_out[88][18][5] + xor_out[89][18][5];
assign sum_out[18][18][5] = xor_out[90][18][5] + xor_out[91][18][5] + xor_out[92][18][5] + xor_out[93][18][5] + xor_out[94][18][5];
assign sum_out[19][18][5] = xor_out[95][18][5] + xor_out[96][18][5] + xor_out[97][18][5] + xor_out[98][18][5] + xor_out[99][18][5];

assign sum_out[0][18][6] = xor_out[0][18][6] + xor_out[1][18][6] + xor_out[2][18][6] + xor_out[3][18][6] + xor_out[4][18][6];
assign sum_out[1][18][6] = xor_out[5][18][6] + xor_out[6][18][6] + xor_out[7][18][6] + xor_out[8][18][6] + xor_out[9][18][6];
assign sum_out[2][18][6] = xor_out[10][18][6] + xor_out[11][18][6] + xor_out[12][18][6] + xor_out[13][18][6] + xor_out[14][18][6];
assign sum_out[3][18][6] = xor_out[15][18][6] + xor_out[16][18][6] + xor_out[17][18][6] + xor_out[18][18][6] + xor_out[19][18][6];
assign sum_out[4][18][6] = xor_out[20][18][6] + xor_out[21][18][6] + xor_out[22][18][6] + xor_out[23][18][6] + xor_out[24][18][6];
assign sum_out[5][18][6] = xor_out[25][18][6] + xor_out[26][18][6] + xor_out[27][18][6] + xor_out[28][18][6] + xor_out[29][18][6];
assign sum_out[6][18][6] = xor_out[30][18][6] + xor_out[31][18][6] + xor_out[32][18][6] + xor_out[33][18][6] + xor_out[34][18][6];
assign sum_out[7][18][6] = xor_out[35][18][6] + xor_out[36][18][6] + xor_out[37][18][6] + xor_out[38][18][6] + xor_out[39][18][6];
assign sum_out[8][18][6] = xor_out[40][18][6] + xor_out[41][18][6] + xor_out[42][18][6] + xor_out[43][18][6] + xor_out[44][18][6];
assign sum_out[9][18][6] = xor_out[45][18][6] + xor_out[46][18][6] + xor_out[47][18][6] + xor_out[48][18][6] + xor_out[49][18][6];
assign sum_out[10][18][6] = xor_out[50][18][6] + xor_out[51][18][6] + xor_out[52][18][6] + xor_out[53][18][6] + xor_out[54][18][6];
assign sum_out[11][18][6] = xor_out[55][18][6] + xor_out[56][18][6] + xor_out[57][18][6] + xor_out[58][18][6] + xor_out[59][18][6];
assign sum_out[12][18][6] = xor_out[60][18][6] + xor_out[61][18][6] + xor_out[62][18][6] + xor_out[63][18][6] + xor_out[64][18][6];
assign sum_out[13][18][6] = xor_out[65][18][6] + xor_out[66][18][6] + xor_out[67][18][6] + xor_out[68][18][6] + xor_out[69][18][6];
assign sum_out[14][18][6] = xor_out[70][18][6] + xor_out[71][18][6] + xor_out[72][18][6] + xor_out[73][18][6] + xor_out[74][18][6];
assign sum_out[15][18][6] = xor_out[75][18][6] + xor_out[76][18][6] + xor_out[77][18][6] + xor_out[78][18][6] + xor_out[79][18][6];
assign sum_out[16][18][6] = xor_out[80][18][6] + xor_out[81][18][6] + xor_out[82][18][6] + xor_out[83][18][6] + xor_out[84][18][6];
assign sum_out[17][18][6] = xor_out[85][18][6] + xor_out[86][18][6] + xor_out[87][18][6] + xor_out[88][18][6] + xor_out[89][18][6];
assign sum_out[18][18][6] = xor_out[90][18][6] + xor_out[91][18][6] + xor_out[92][18][6] + xor_out[93][18][6] + xor_out[94][18][6];
assign sum_out[19][18][6] = xor_out[95][18][6] + xor_out[96][18][6] + xor_out[97][18][6] + xor_out[98][18][6] + xor_out[99][18][6];

assign sum_out[0][18][7] = xor_out[0][18][7] + xor_out[1][18][7] + xor_out[2][18][7] + xor_out[3][18][7] + xor_out[4][18][7];
assign sum_out[1][18][7] = xor_out[5][18][7] + xor_out[6][18][7] + xor_out[7][18][7] + xor_out[8][18][7] + xor_out[9][18][7];
assign sum_out[2][18][7] = xor_out[10][18][7] + xor_out[11][18][7] + xor_out[12][18][7] + xor_out[13][18][7] + xor_out[14][18][7];
assign sum_out[3][18][7] = xor_out[15][18][7] + xor_out[16][18][7] + xor_out[17][18][7] + xor_out[18][18][7] + xor_out[19][18][7];
assign sum_out[4][18][7] = xor_out[20][18][7] + xor_out[21][18][7] + xor_out[22][18][7] + xor_out[23][18][7] + xor_out[24][18][7];
assign sum_out[5][18][7] = xor_out[25][18][7] + xor_out[26][18][7] + xor_out[27][18][7] + xor_out[28][18][7] + xor_out[29][18][7];
assign sum_out[6][18][7] = xor_out[30][18][7] + xor_out[31][18][7] + xor_out[32][18][7] + xor_out[33][18][7] + xor_out[34][18][7];
assign sum_out[7][18][7] = xor_out[35][18][7] + xor_out[36][18][7] + xor_out[37][18][7] + xor_out[38][18][7] + xor_out[39][18][7];
assign sum_out[8][18][7] = xor_out[40][18][7] + xor_out[41][18][7] + xor_out[42][18][7] + xor_out[43][18][7] + xor_out[44][18][7];
assign sum_out[9][18][7] = xor_out[45][18][7] + xor_out[46][18][7] + xor_out[47][18][7] + xor_out[48][18][7] + xor_out[49][18][7];
assign sum_out[10][18][7] = xor_out[50][18][7] + xor_out[51][18][7] + xor_out[52][18][7] + xor_out[53][18][7] + xor_out[54][18][7];
assign sum_out[11][18][7] = xor_out[55][18][7] + xor_out[56][18][7] + xor_out[57][18][7] + xor_out[58][18][7] + xor_out[59][18][7];
assign sum_out[12][18][7] = xor_out[60][18][7] + xor_out[61][18][7] + xor_out[62][18][7] + xor_out[63][18][7] + xor_out[64][18][7];
assign sum_out[13][18][7] = xor_out[65][18][7] + xor_out[66][18][7] + xor_out[67][18][7] + xor_out[68][18][7] + xor_out[69][18][7];
assign sum_out[14][18][7] = xor_out[70][18][7] + xor_out[71][18][7] + xor_out[72][18][7] + xor_out[73][18][7] + xor_out[74][18][7];
assign sum_out[15][18][7] = xor_out[75][18][7] + xor_out[76][18][7] + xor_out[77][18][7] + xor_out[78][18][7] + xor_out[79][18][7];
assign sum_out[16][18][7] = xor_out[80][18][7] + xor_out[81][18][7] + xor_out[82][18][7] + xor_out[83][18][7] + xor_out[84][18][7];
assign sum_out[17][18][7] = xor_out[85][18][7] + xor_out[86][18][7] + xor_out[87][18][7] + xor_out[88][18][7] + xor_out[89][18][7];
assign sum_out[18][18][7] = xor_out[90][18][7] + xor_out[91][18][7] + xor_out[92][18][7] + xor_out[93][18][7] + xor_out[94][18][7];
assign sum_out[19][18][7] = xor_out[95][18][7] + xor_out[96][18][7] + xor_out[97][18][7] + xor_out[98][18][7] + xor_out[99][18][7];

assign sum_out[0][18][8] = xor_out[0][18][8] + xor_out[1][18][8] + xor_out[2][18][8] + xor_out[3][18][8] + xor_out[4][18][8];
assign sum_out[1][18][8] = xor_out[5][18][8] + xor_out[6][18][8] + xor_out[7][18][8] + xor_out[8][18][8] + xor_out[9][18][8];
assign sum_out[2][18][8] = xor_out[10][18][8] + xor_out[11][18][8] + xor_out[12][18][8] + xor_out[13][18][8] + xor_out[14][18][8];
assign sum_out[3][18][8] = xor_out[15][18][8] + xor_out[16][18][8] + xor_out[17][18][8] + xor_out[18][18][8] + xor_out[19][18][8];
assign sum_out[4][18][8] = xor_out[20][18][8] + xor_out[21][18][8] + xor_out[22][18][8] + xor_out[23][18][8] + xor_out[24][18][8];
assign sum_out[5][18][8] = xor_out[25][18][8] + xor_out[26][18][8] + xor_out[27][18][8] + xor_out[28][18][8] + xor_out[29][18][8];
assign sum_out[6][18][8] = xor_out[30][18][8] + xor_out[31][18][8] + xor_out[32][18][8] + xor_out[33][18][8] + xor_out[34][18][8];
assign sum_out[7][18][8] = xor_out[35][18][8] + xor_out[36][18][8] + xor_out[37][18][8] + xor_out[38][18][8] + xor_out[39][18][8];
assign sum_out[8][18][8] = xor_out[40][18][8] + xor_out[41][18][8] + xor_out[42][18][8] + xor_out[43][18][8] + xor_out[44][18][8];
assign sum_out[9][18][8] = xor_out[45][18][8] + xor_out[46][18][8] + xor_out[47][18][8] + xor_out[48][18][8] + xor_out[49][18][8];
assign sum_out[10][18][8] = xor_out[50][18][8] + xor_out[51][18][8] + xor_out[52][18][8] + xor_out[53][18][8] + xor_out[54][18][8];
assign sum_out[11][18][8] = xor_out[55][18][8] + xor_out[56][18][8] + xor_out[57][18][8] + xor_out[58][18][8] + xor_out[59][18][8];
assign sum_out[12][18][8] = xor_out[60][18][8] + xor_out[61][18][8] + xor_out[62][18][8] + xor_out[63][18][8] + xor_out[64][18][8];
assign sum_out[13][18][8] = xor_out[65][18][8] + xor_out[66][18][8] + xor_out[67][18][8] + xor_out[68][18][8] + xor_out[69][18][8];
assign sum_out[14][18][8] = xor_out[70][18][8] + xor_out[71][18][8] + xor_out[72][18][8] + xor_out[73][18][8] + xor_out[74][18][8];
assign sum_out[15][18][8] = xor_out[75][18][8] + xor_out[76][18][8] + xor_out[77][18][8] + xor_out[78][18][8] + xor_out[79][18][8];
assign sum_out[16][18][8] = xor_out[80][18][8] + xor_out[81][18][8] + xor_out[82][18][8] + xor_out[83][18][8] + xor_out[84][18][8];
assign sum_out[17][18][8] = xor_out[85][18][8] + xor_out[86][18][8] + xor_out[87][18][8] + xor_out[88][18][8] + xor_out[89][18][8];
assign sum_out[18][18][8] = xor_out[90][18][8] + xor_out[91][18][8] + xor_out[92][18][8] + xor_out[93][18][8] + xor_out[94][18][8];
assign sum_out[19][18][8] = xor_out[95][18][8] + xor_out[96][18][8] + xor_out[97][18][8] + xor_out[98][18][8] + xor_out[99][18][8];

assign sum_out[0][18][9] = xor_out[0][18][9] + xor_out[1][18][9] + xor_out[2][18][9] + xor_out[3][18][9] + xor_out[4][18][9];
assign sum_out[1][18][9] = xor_out[5][18][9] + xor_out[6][18][9] + xor_out[7][18][9] + xor_out[8][18][9] + xor_out[9][18][9];
assign sum_out[2][18][9] = xor_out[10][18][9] + xor_out[11][18][9] + xor_out[12][18][9] + xor_out[13][18][9] + xor_out[14][18][9];
assign sum_out[3][18][9] = xor_out[15][18][9] + xor_out[16][18][9] + xor_out[17][18][9] + xor_out[18][18][9] + xor_out[19][18][9];
assign sum_out[4][18][9] = xor_out[20][18][9] + xor_out[21][18][9] + xor_out[22][18][9] + xor_out[23][18][9] + xor_out[24][18][9];
assign sum_out[5][18][9] = xor_out[25][18][9] + xor_out[26][18][9] + xor_out[27][18][9] + xor_out[28][18][9] + xor_out[29][18][9];
assign sum_out[6][18][9] = xor_out[30][18][9] + xor_out[31][18][9] + xor_out[32][18][9] + xor_out[33][18][9] + xor_out[34][18][9];
assign sum_out[7][18][9] = xor_out[35][18][9] + xor_out[36][18][9] + xor_out[37][18][9] + xor_out[38][18][9] + xor_out[39][18][9];
assign sum_out[8][18][9] = xor_out[40][18][9] + xor_out[41][18][9] + xor_out[42][18][9] + xor_out[43][18][9] + xor_out[44][18][9];
assign sum_out[9][18][9] = xor_out[45][18][9] + xor_out[46][18][9] + xor_out[47][18][9] + xor_out[48][18][9] + xor_out[49][18][9];
assign sum_out[10][18][9] = xor_out[50][18][9] + xor_out[51][18][9] + xor_out[52][18][9] + xor_out[53][18][9] + xor_out[54][18][9];
assign sum_out[11][18][9] = xor_out[55][18][9] + xor_out[56][18][9] + xor_out[57][18][9] + xor_out[58][18][9] + xor_out[59][18][9];
assign sum_out[12][18][9] = xor_out[60][18][9] + xor_out[61][18][9] + xor_out[62][18][9] + xor_out[63][18][9] + xor_out[64][18][9];
assign sum_out[13][18][9] = xor_out[65][18][9] + xor_out[66][18][9] + xor_out[67][18][9] + xor_out[68][18][9] + xor_out[69][18][9];
assign sum_out[14][18][9] = xor_out[70][18][9] + xor_out[71][18][9] + xor_out[72][18][9] + xor_out[73][18][9] + xor_out[74][18][9];
assign sum_out[15][18][9] = xor_out[75][18][9] + xor_out[76][18][9] + xor_out[77][18][9] + xor_out[78][18][9] + xor_out[79][18][9];
assign sum_out[16][18][9] = xor_out[80][18][9] + xor_out[81][18][9] + xor_out[82][18][9] + xor_out[83][18][9] + xor_out[84][18][9];
assign sum_out[17][18][9] = xor_out[85][18][9] + xor_out[86][18][9] + xor_out[87][18][9] + xor_out[88][18][9] + xor_out[89][18][9];
assign sum_out[18][18][9] = xor_out[90][18][9] + xor_out[91][18][9] + xor_out[92][18][9] + xor_out[93][18][9] + xor_out[94][18][9];
assign sum_out[19][18][9] = xor_out[95][18][9] + xor_out[96][18][9] + xor_out[97][18][9] + xor_out[98][18][9] + xor_out[99][18][9];

assign sum_out[0][18][10] = xor_out[0][18][10] + xor_out[1][18][10] + xor_out[2][18][10] + xor_out[3][18][10] + xor_out[4][18][10];
assign sum_out[1][18][10] = xor_out[5][18][10] + xor_out[6][18][10] + xor_out[7][18][10] + xor_out[8][18][10] + xor_out[9][18][10];
assign sum_out[2][18][10] = xor_out[10][18][10] + xor_out[11][18][10] + xor_out[12][18][10] + xor_out[13][18][10] + xor_out[14][18][10];
assign sum_out[3][18][10] = xor_out[15][18][10] + xor_out[16][18][10] + xor_out[17][18][10] + xor_out[18][18][10] + xor_out[19][18][10];
assign sum_out[4][18][10] = xor_out[20][18][10] + xor_out[21][18][10] + xor_out[22][18][10] + xor_out[23][18][10] + xor_out[24][18][10];
assign sum_out[5][18][10] = xor_out[25][18][10] + xor_out[26][18][10] + xor_out[27][18][10] + xor_out[28][18][10] + xor_out[29][18][10];
assign sum_out[6][18][10] = xor_out[30][18][10] + xor_out[31][18][10] + xor_out[32][18][10] + xor_out[33][18][10] + xor_out[34][18][10];
assign sum_out[7][18][10] = xor_out[35][18][10] + xor_out[36][18][10] + xor_out[37][18][10] + xor_out[38][18][10] + xor_out[39][18][10];
assign sum_out[8][18][10] = xor_out[40][18][10] + xor_out[41][18][10] + xor_out[42][18][10] + xor_out[43][18][10] + xor_out[44][18][10];
assign sum_out[9][18][10] = xor_out[45][18][10] + xor_out[46][18][10] + xor_out[47][18][10] + xor_out[48][18][10] + xor_out[49][18][10];
assign sum_out[10][18][10] = xor_out[50][18][10] + xor_out[51][18][10] + xor_out[52][18][10] + xor_out[53][18][10] + xor_out[54][18][10];
assign sum_out[11][18][10] = xor_out[55][18][10] + xor_out[56][18][10] + xor_out[57][18][10] + xor_out[58][18][10] + xor_out[59][18][10];
assign sum_out[12][18][10] = xor_out[60][18][10] + xor_out[61][18][10] + xor_out[62][18][10] + xor_out[63][18][10] + xor_out[64][18][10];
assign sum_out[13][18][10] = xor_out[65][18][10] + xor_out[66][18][10] + xor_out[67][18][10] + xor_out[68][18][10] + xor_out[69][18][10];
assign sum_out[14][18][10] = xor_out[70][18][10] + xor_out[71][18][10] + xor_out[72][18][10] + xor_out[73][18][10] + xor_out[74][18][10];
assign sum_out[15][18][10] = xor_out[75][18][10] + xor_out[76][18][10] + xor_out[77][18][10] + xor_out[78][18][10] + xor_out[79][18][10];
assign sum_out[16][18][10] = xor_out[80][18][10] + xor_out[81][18][10] + xor_out[82][18][10] + xor_out[83][18][10] + xor_out[84][18][10];
assign sum_out[17][18][10] = xor_out[85][18][10] + xor_out[86][18][10] + xor_out[87][18][10] + xor_out[88][18][10] + xor_out[89][18][10];
assign sum_out[18][18][10] = xor_out[90][18][10] + xor_out[91][18][10] + xor_out[92][18][10] + xor_out[93][18][10] + xor_out[94][18][10];
assign sum_out[19][18][10] = xor_out[95][18][10] + xor_out[96][18][10] + xor_out[97][18][10] + xor_out[98][18][10] + xor_out[99][18][10];

assign sum_out[0][18][11] = xor_out[0][18][11] + xor_out[1][18][11] + xor_out[2][18][11] + xor_out[3][18][11] + xor_out[4][18][11];
assign sum_out[1][18][11] = xor_out[5][18][11] + xor_out[6][18][11] + xor_out[7][18][11] + xor_out[8][18][11] + xor_out[9][18][11];
assign sum_out[2][18][11] = xor_out[10][18][11] + xor_out[11][18][11] + xor_out[12][18][11] + xor_out[13][18][11] + xor_out[14][18][11];
assign sum_out[3][18][11] = xor_out[15][18][11] + xor_out[16][18][11] + xor_out[17][18][11] + xor_out[18][18][11] + xor_out[19][18][11];
assign sum_out[4][18][11] = xor_out[20][18][11] + xor_out[21][18][11] + xor_out[22][18][11] + xor_out[23][18][11] + xor_out[24][18][11];
assign sum_out[5][18][11] = xor_out[25][18][11] + xor_out[26][18][11] + xor_out[27][18][11] + xor_out[28][18][11] + xor_out[29][18][11];
assign sum_out[6][18][11] = xor_out[30][18][11] + xor_out[31][18][11] + xor_out[32][18][11] + xor_out[33][18][11] + xor_out[34][18][11];
assign sum_out[7][18][11] = xor_out[35][18][11] + xor_out[36][18][11] + xor_out[37][18][11] + xor_out[38][18][11] + xor_out[39][18][11];
assign sum_out[8][18][11] = xor_out[40][18][11] + xor_out[41][18][11] + xor_out[42][18][11] + xor_out[43][18][11] + xor_out[44][18][11];
assign sum_out[9][18][11] = xor_out[45][18][11] + xor_out[46][18][11] + xor_out[47][18][11] + xor_out[48][18][11] + xor_out[49][18][11];
assign sum_out[10][18][11] = xor_out[50][18][11] + xor_out[51][18][11] + xor_out[52][18][11] + xor_out[53][18][11] + xor_out[54][18][11];
assign sum_out[11][18][11] = xor_out[55][18][11] + xor_out[56][18][11] + xor_out[57][18][11] + xor_out[58][18][11] + xor_out[59][18][11];
assign sum_out[12][18][11] = xor_out[60][18][11] + xor_out[61][18][11] + xor_out[62][18][11] + xor_out[63][18][11] + xor_out[64][18][11];
assign sum_out[13][18][11] = xor_out[65][18][11] + xor_out[66][18][11] + xor_out[67][18][11] + xor_out[68][18][11] + xor_out[69][18][11];
assign sum_out[14][18][11] = xor_out[70][18][11] + xor_out[71][18][11] + xor_out[72][18][11] + xor_out[73][18][11] + xor_out[74][18][11];
assign sum_out[15][18][11] = xor_out[75][18][11] + xor_out[76][18][11] + xor_out[77][18][11] + xor_out[78][18][11] + xor_out[79][18][11];
assign sum_out[16][18][11] = xor_out[80][18][11] + xor_out[81][18][11] + xor_out[82][18][11] + xor_out[83][18][11] + xor_out[84][18][11];
assign sum_out[17][18][11] = xor_out[85][18][11] + xor_out[86][18][11] + xor_out[87][18][11] + xor_out[88][18][11] + xor_out[89][18][11];
assign sum_out[18][18][11] = xor_out[90][18][11] + xor_out[91][18][11] + xor_out[92][18][11] + xor_out[93][18][11] + xor_out[94][18][11];
assign sum_out[19][18][11] = xor_out[95][18][11] + xor_out[96][18][11] + xor_out[97][18][11] + xor_out[98][18][11] + xor_out[99][18][11];

assign sum_out[0][18][12] = xor_out[0][18][12] + xor_out[1][18][12] + xor_out[2][18][12] + xor_out[3][18][12] + xor_out[4][18][12];
assign sum_out[1][18][12] = xor_out[5][18][12] + xor_out[6][18][12] + xor_out[7][18][12] + xor_out[8][18][12] + xor_out[9][18][12];
assign sum_out[2][18][12] = xor_out[10][18][12] + xor_out[11][18][12] + xor_out[12][18][12] + xor_out[13][18][12] + xor_out[14][18][12];
assign sum_out[3][18][12] = xor_out[15][18][12] + xor_out[16][18][12] + xor_out[17][18][12] + xor_out[18][18][12] + xor_out[19][18][12];
assign sum_out[4][18][12] = xor_out[20][18][12] + xor_out[21][18][12] + xor_out[22][18][12] + xor_out[23][18][12] + xor_out[24][18][12];
assign sum_out[5][18][12] = xor_out[25][18][12] + xor_out[26][18][12] + xor_out[27][18][12] + xor_out[28][18][12] + xor_out[29][18][12];
assign sum_out[6][18][12] = xor_out[30][18][12] + xor_out[31][18][12] + xor_out[32][18][12] + xor_out[33][18][12] + xor_out[34][18][12];
assign sum_out[7][18][12] = xor_out[35][18][12] + xor_out[36][18][12] + xor_out[37][18][12] + xor_out[38][18][12] + xor_out[39][18][12];
assign sum_out[8][18][12] = xor_out[40][18][12] + xor_out[41][18][12] + xor_out[42][18][12] + xor_out[43][18][12] + xor_out[44][18][12];
assign sum_out[9][18][12] = xor_out[45][18][12] + xor_out[46][18][12] + xor_out[47][18][12] + xor_out[48][18][12] + xor_out[49][18][12];
assign sum_out[10][18][12] = xor_out[50][18][12] + xor_out[51][18][12] + xor_out[52][18][12] + xor_out[53][18][12] + xor_out[54][18][12];
assign sum_out[11][18][12] = xor_out[55][18][12] + xor_out[56][18][12] + xor_out[57][18][12] + xor_out[58][18][12] + xor_out[59][18][12];
assign sum_out[12][18][12] = xor_out[60][18][12] + xor_out[61][18][12] + xor_out[62][18][12] + xor_out[63][18][12] + xor_out[64][18][12];
assign sum_out[13][18][12] = xor_out[65][18][12] + xor_out[66][18][12] + xor_out[67][18][12] + xor_out[68][18][12] + xor_out[69][18][12];
assign sum_out[14][18][12] = xor_out[70][18][12] + xor_out[71][18][12] + xor_out[72][18][12] + xor_out[73][18][12] + xor_out[74][18][12];
assign sum_out[15][18][12] = xor_out[75][18][12] + xor_out[76][18][12] + xor_out[77][18][12] + xor_out[78][18][12] + xor_out[79][18][12];
assign sum_out[16][18][12] = xor_out[80][18][12] + xor_out[81][18][12] + xor_out[82][18][12] + xor_out[83][18][12] + xor_out[84][18][12];
assign sum_out[17][18][12] = xor_out[85][18][12] + xor_out[86][18][12] + xor_out[87][18][12] + xor_out[88][18][12] + xor_out[89][18][12];
assign sum_out[18][18][12] = xor_out[90][18][12] + xor_out[91][18][12] + xor_out[92][18][12] + xor_out[93][18][12] + xor_out[94][18][12];
assign sum_out[19][18][12] = xor_out[95][18][12] + xor_out[96][18][12] + xor_out[97][18][12] + xor_out[98][18][12] + xor_out[99][18][12];

assign sum_out[0][18][13] = xor_out[0][18][13] + xor_out[1][18][13] + xor_out[2][18][13] + xor_out[3][18][13] + xor_out[4][18][13];
assign sum_out[1][18][13] = xor_out[5][18][13] + xor_out[6][18][13] + xor_out[7][18][13] + xor_out[8][18][13] + xor_out[9][18][13];
assign sum_out[2][18][13] = xor_out[10][18][13] + xor_out[11][18][13] + xor_out[12][18][13] + xor_out[13][18][13] + xor_out[14][18][13];
assign sum_out[3][18][13] = xor_out[15][18][13] + xor_out[16][18][13] + xor_out[17][18][13] + xor_out[18][18][13] + xor_out[19][18][13];
assign sum_out[4][18][13] = xor_out[20][18][13] + xor_out[21][18][13] + xor_out[22][18][13] + xor_out[23][18][13] + xor_out[24][18][13];
assign sum_out[5][18][13] = xor_out[25][18][13] + xor_out[26][18][13] + xor_out[27][18][13] + xor_out[28][18][13] + xor_out[29][18][13];
assign sum_out[6][18][13] = xor_out[30][18][13] + xor_out[31][18][13] + xor_out[32][18][13] + xor_out[33][18][13] + xor_out[34][18][13];
assign sum_out[7][18][13] = xor_out[35][18][13] + xor_out[36][18][13] + xor_out[37][18][13] + xor_out[38][18][13] + xor_out[39][18][13];
assign sum_out[8][18][13] = xor_out[40][18][13] + xor_out[41][18][13] + xor_out[42][18][13] + xor_out[43][18][13] + xor_out[44][18][13];
assign sum_out[9][18][13] = xor_out[45][18][13] + xor_out[46][18][13] + xor_out[47][18][13] + xor_out[48][18][13] + xor_out[49][18][13];
assign sum_out[10][18][13] = xor_out[50][18][13] + xor_out[51][18][13] + xor_out[52][18][13] + xor_out[53][18][13] + xor_out[54][18][13];
assign sum_out[11][18][13] = xor_out[55][18][13] + xor_out[56][18][13] + xor_out[57][18][13] + xor_out[58][18][13] + xor_out[59][18][13];
assign sum_out[12][18][13] = xor_out[60][18][13] + xor_out[61][18][13] + xor_out[62][18][13] + xor_out[63][18][13] + xor_out[64][18][13];
assign sum_out[13][18][13] = xor_out[65][18][13] + xor_out[66][18][13] + xor_out[67][18][13] + xor_out[68][18][13] + xor_out[69][18][13];
assign sum_out[14][18][13] = xor_out[70][18][13] + xor_out[71][18][13] + xor_out[72][18][13] + xor_out[73][18][13] + xor_out[74][18][13];
assign sum_out[15][18][13] = xor_out[75][18][13] + xor_out[76][18][13] + xor_out[77][18][13] + xor_out[78][18][13] + xor_out[79][18][13];
assign sum_out[16][18][13] = xor_out[80][18][13] + xor_out[81][18][13] + xor_out[82][18][13] + xor_out[83][18][13] + xor_out[84][18][13];
assign sum_out[17][18][13] = xor_out[85][18][13] + xor_out[86][18][13] + xor_out[87][18][13] + xor_out[88][18][13] + xor_out[89][18][13];
assign sum_out[18][18][13] = xor_out[90][18][13] + xor_out[91][18][13] + xor_out[92][18][13] + xor_out[93][18][13] + xor_out[94][18][13];
assign sum_out[19][18][13] = xor_out[95][18][13] + xor_out[96][18][13] + xor_out[97][18][13] + xor_out[98][18][13] + xor_out[99][18][13];

assign sum_out[0][18][14] = xor_out[0][18][14] + xor_out[1][18][14] + xor_out[2][18][14] + xor_out[3][18][14] + xor_out[4][18][14];
assign sum_out[1][18][14] = xor_out[5][18][14] + xor_out[6][18][14] + xor_out[7][18][14] + xor_out[8][18][14] + xor_out[9][18][14];
assign sum_out[2][18][14] = xor_out[10][18][14] + xor_out[11][18][14] + xor_out[12][18][14] + xor_out[13][18][14] + xor_out[14][18][14];
assign sum_out[3][18][14] = xor_out[15][18][14] + xor_out[16][18][14] + xor_out[17][18][14] + xor_out[18][18][14] + xor_out[19][18][14];
assign sum_out[4][18][14] = xor_out[20][18][14] + xor_out[21][18][14] + xor_out[22][18][14] + xor_out[23][18][14] + xor_out[24][18][14];
assign sum_out[5][18][14] = xor_out[25][18][14] + xor_out[26][18][14] + xor_out[27][18][14] + xor_out[28][18][14] + xor_out[29][18][14];
assign sum_out[6][18][14] = xor_out[30][18][14] + xor_out[31][18][14] + xor_out[32][18][14] + xor_out[33][18][14] + xor_out[34][18][14];
assign sum_out[7][18][14] = xor_out[35][18][14] + xor_out[36][18][14] + xor_out[37][18][14] + xor_out[38][18][14] + xor_out[39][18][14];
assign sum_out[8][18][14] = xor_out[40][18][14] + xor_out[41][18][14] + xor_out[42][18][14] + xor_out[43][18][14] + xor_out[44][18][14];
assign sum_out[9][18][14] = xor_out[45][18][14] + xor_out[46][18][14] + xor_out[47][18][14] + xor_out[48][18][14] + xor_out[49][18][14];
assign sum_out[10][18][14] = xor_out[50][18][14] + xor_out[51][18][14] + xor_out[52][18][14] + xor_out[53][18][14] + xor_out[54][18][14];
assign sum_out[11][18][14] = xor_out[55][18][14] + xor_out[56][18][14] + xor_out[57][18][14] + xor_out[58][18][14] + xor_out[59][18][14];
assign sum_out[12][18][14] = xor_out[60][18][14] + xor_out[61][18][14] + xor_out[62][18][14] + xor_out[63][18][14] + xor_out[64][18][14];
assign sum_out[13][18][14] = xor_out[65][18][14] + xor_out[66][18][14] + xor_out[67][18][14] + xor_out[68][18][14] + xor_out[69][18][14];
assign sum_out[14][18][14] = xor_out[70][18][14] + xor_out[71][18][14] + xor_out[72][18][14] + xor_out[73][18][14] + xor_out[74][18][14];
assign sum_out[15][18][14] = xor_out[75][18][14] + xor_out[76][18][14] + xor_out[77][18][14] + xor_out[78][18][14] + xor_out[79][18][14];
assign sum_out[16][18][14] = xor_out[80][18][14] + xor_out[81][18][14] + xor_out[82][18][14] + xor_out[83][18][14] + xor_out[84][18][14];
assign sum_out[17][18][14] = xor_out[85][18][14] + xor_out[86][18][14] + xor_out[87][18][14] + xor_out[88][18][14] + xor_out[89][18][14];
assign sum_out[18][18][14] = xor_out[90][18][14] + xor_out[91][18][14] + xor_out[92][18][14] + xor_out[93][18][14] + xor_out[94][18][14];
assign sum_out[19][18][14] = xor_out[95][18][14] + xor_out[96][18][14] + xor_out[97][18][14] + xor_out[98][18][14] + xor_out[99][18][14];

assign sum_out[0][18][15] = xor_out[0][18][15] + xor_out[1][18][15] + xor_out[2][18][15] + xor_out[3][18][15] + xor_out[4][18][15];
assign sum_out[1][18][15] = xor_out[5][18][15] + xor_out[6][18][15] + xor_out[7][18][15] + xor_out[8][18][15] + xor_out[9][18][15];
assign sum_out[2][18][15] = xor_out[10][18][15] + xor_out[11][18][15] + xor_out[12][18][15] + xor_out[13][18][15] + xor_out[14][18][15];
assign sum_out[3][18][15] = xor_out[15][18][15] + xor_out[16][18][15] + xor_out[17][18][15] + xor_out[18][18][15] + xor_out[19][18][15];
assign sum_out[4][18][15] = xor_out[20][18][15] + xor_out[21][18][15] + xor_out[22][18][15] + xor_out[23][18][15] + xor_out[24][18][15];
assign sum_out[5][18][15] = xor_out[25][18][15] + xor_out[26][18][15] + xor_out[27][18][15] + xor_out[28][18][15] + xor_out[29][18][15];
assign sum_out[6][18][15] = xor_out[30][18][15] + xor_out[31][18][15] + xor_out[32][18][15] + xor_out[33][18][15] + xor_out[34][18][15];
assign sum_out[7][18][15] = xor_out[35][18][15] + xor_out[36][18][15] + xor_out[37][18][15] + xor_out[38][18][15] + xor_out[39][18][15];
assign sum_out[8][18][15] = xor_out[40][18][15] + xor_out[41][18][15] + xor_out[42][18][15] + xor_out[43][18][15] + xor_out[44][18][15];
assign sum_out[9][18][15] = xor_out[45][18][15] + xor_out[46][18][15] + xor_out[47][18][15] + xor_out[48][18][15] + xor_out[49][18][15];
assign sum_out[10][18][15] = xor_out[50][18][15] + xor_out[51][18][15] + xor_out[52][18][15] + xor_out[53][18][15] + xor_out[54][18][15];
assign sum_out[11][18][15] = xor_out[55][18][15] + xor_out[56][18][15] + xor_out[57][18][15] + xor_out[58][18][15] + xor_out[59][18][15];
assign sum_out[12][18][15] = xor_out[60][18][15] + xor_out[61][18][15] + xor_out[62][18][15] + xor_out[63][18][15] + xor_out[64][18][15];
assign sum_out[13][18][15] = xor_out[65][18][15] + xor_out[66][18][15] + xor_out[67][18][15] + xor_out[68][18][15] + xor_out[69][18][15];
assign sum_out[14][18][15] = xor_out[70][18][15] + xor_out[71][18][15] + xor_out[72][18][15] + xor_out[73][18][15] + xor_out[74][18][15];
assign sum_out[15][18][15] = xor_out[75][18][15] + xor_out[76][18][15] + xor_out[77][18][15] + xor_out[78][18][15] + xor_out[79][18][15];
assign sum_out[16][18][15] = xor_out[80][18][15] + xor_out[81][18][15] + xor_out[82][18][15] + xor_out[83][18][15] + xor_out[84][18][15];
assign sum_out[17][18][15] = xor_out[85][18][15] + xor_out[86][18][15] + xor_out[87][18][15] + xor_out[88][18][15] + xor_out[89][18][15];
assign sum_out[18][18][15] = xor_out[90][18][15] + xor_out[91][18][15] + xor_out[92][18][15] + xor_out[93][18][15] + xor_out[94][18][15];
assign sum_out[19][18][15] = xor_out[95][18][15] + xor_out[96][18][15] + xor_out[97][18][15] + xor_out[98][18][15] + xor_out[99][18][15];

assign sum_out[0][18][16] = xor_out[0][18][16] + xor_out[1][18][16] + xor_out[2][18][16] + xor_out[3][18][16] + xor_out[4][18][16];
assign sum_out[1][18][16] = xor_out[5][18][16] + xor_out[6][18][16] + xor_out[7][18][16] + xor_out[8][18][16] + xor_out[9][18][16];
assign sum_out[2][18][16] = xor_out[10][18][16] + xor_out[11][18][16] + xor_out[12][18][16] + xor_out[13][18][16] + xor_out[14][18][16];
assign sum_out[3][18][16] = xor_out[15][18][16] + xor_out[16][18][16] + xor_out[17][18][16] + xor_out[18][18][16] + xor_out[19][18][16];
assign sum_out[4][18][16] = xor_out[20][18][16] + xor_out[21][18][16] + xor_out[22][18][16] + xor_out[23][18][16] + xor_out[24][18][16];
assign sum_out[5][18][16] = xor_out[25][18][16] + xor_out[26][18][16] + xor_out[27][18][16] + xor_out[28][18][16] + xor_out[29][18][16];
assign sum_out[6][18][16] = xor_out[30][18][16] + xor_out[31][18][16] + xor_out[32][18][16] + xor_out[33][18][16] + xor_out[34][18][16];
assign sum_out[7][18][16] = xor_out[35][18][16] + xor_out[36][18][16] + xor_out[37][18][16] + xor_out[38][18][16] + xor_out[39][18][16];
assign sum_out[8][18][16] = xor_out[40][18][16] + xor_out[41][18][16] + xor_out[42][18][16] + xor_out[43][18][16] + xor_out[44][18][16];
assign sum_out[9][18][16] = xor_out[45][18][16] + xor_out[46][18][16] + xor_out[47][18][16] + xor_out[48][18][16] + xor_out[49][18][16];
assign sum_out[10][18][16] = xor_out[50][18][16] + xor_out[51][18][16] + xor_out[52][18][16] + xor_out[53][18][16] + xor_out[54][18][16];
assign sum_out[11][18][16] = xor_out[55][18][16] + xor_out[56][18][16] + xor_out[57][18][16] + xor_out[58][18][16] + xor_out[59][18][16];
assign sum_out[12][18][16] = xor_out[60][18][16] + xor_out[61][18][16] + xor_out[62][18][16] + xor_out[63][18][16] + xor_out[64][18][16];
assign sum_out[13][18][16] = xor_out[65][18][16] + xor_out[66][18][16] + xor_out[67][18][16] + xor_out[68][18][16] + xor_out[69][18][16];
assign sum_out[14][18][16] = xor_out[70][18][16] + xor_out[71][18][16] + xor_out[72][18][16] + xor_out[73][18][16] + xor_out[74][18][16];
assign sum_out[15][18][16] = xor_out[75][18][16] + xor_out[76][18][16] + xor_out[77][18][16] + xor_out[78][18][16] + xor_out[79][18][16];
assign sum_out[16][18][16] = xor_out[80][18][16] + xor_out[81][18][16] + xor_out[82][18][16] + xor_out[83][18][16] + xor_out[84][18][16];
assign sum_out[17][18][16] = xor_out[85][18][16] + xor_out[86][18][16] + xor_out[87][18][16] + xor_out[88][18][16] + xor_out[89][18][16];
assign sum_out[18][18][16] = xor_out[90][18][16] + xor_out[91][18][16] + xor_out[92][18][16] + xor_out[93][18][16] + xor_out[94][18][16];
assign sum_out[19][18][16] = xor_out[95][18][16] + xor_out[96][18][16] + xor_out[97][18][16] + xor_out[98][18][16] + xor_out[99][18][16];

assign sum_out[0][18][17] = xor_out[0][18][17] + xor_out[1][18][17] + xor_out[2][18][17] + xor_out[3][18][17] + xor_out[4][18][17];
assign sum_out[1][18][17] = xor_out[5][18][17] + xor_out[6][18][17] + xor_out[7][18][17] + xor_out[8][18][17] + xor_out[9][18][17];
assign sum_out[2][18][17] = xor_out[10][18][17] + xor_out[11][18][17] + xor_out[12][18][17] + xor_out[13][18][17] + xor_out[14][18][17];
assign sum_out[3][18][17] = xor_out[15][18][17] + xor_out[16][18][17] + xor_out[17][18][17] + xor_out[18][18][17] + xor_out[19][18][17];
assign sum_out[4][18][17] = xor_out[20][18][17] + xor_out[21][18][17] + xor_out[22][18][17] + xor_out[23][18][17] + xor_out[24][18][17];
assign sum_out[5][18][17] = xor_out[25][18][17] + xor_out[26][18][17] + xor_out[27][18][17] + xor_out[28][18][17] + xor_out[29][18][17];
assign sum_out[6][18][17] = xor_out[30][18][17] + xor_out[31][18][17] + xor_out[32][18][17] + xor_out[33][18][17] + xor_out[34][18][17];
assign sum_out[7][18][17] = xor_out[35][18][17] + xor_out[36][18][17] + xor_out[37][18][17] + xor_out[38][18][17] + xor_out[39][18][17];
assign sum_out[8][18][17] = xor_out[40][18][17] + xor_out[41][18][17] + xor_out[42][18][17] + xor_out[43][18][17] + xor_out[44][18][17];
assign sum_out[9][18][17] = xor_out[45][18][17] + xor_out[46][18][17] + xor_out[47][18][17] + xor_out[48][18][17] + xor_out[49][18][17];
assign sum_out[10][18][17] = xor_out[50][18][17] + xor_out[51][18][17] + xor_out[52][18][17] + xor_out[53][18][17] + xor_out[54][18][17];
assign sum_out[11][18][17] = xor_out[55][18][17] + xor_out[56][18][17] + xor_out[57][18][17] + xor_out[58][18][17] + xor_out[59][18][17];
assign sum_out[12][18][17] = xor_out[60][18][17] + xor_out[61][18][17] + xor_out[62][18][17] + xor_out[63][18][17] + xor_out[64][18][17];
assign sum_out[13][18][17] = xor_out[65][18][17] + xor_out[66][18][17] + xor_out[67][18][17] + xor_out[68][18][17] + xor_out[69][18][17];
assign sum_out[14][18][17] = xor_out[70][18][17] + xor_out[71][18][17] + xor_out[72][18][17] + xor_out[73][18][17] + xor_out[74][18][17];
assign sum_out[15][18][17] = xor_out[75][18][17] + xor_out[76][18][17] + xor_out[77][18][17] + xor_out[78][18][17] + xor_out[79][18][17];
assign sum_out[16][18][17] = xor_out[80][18][17] + xor_out[81][18][17] + xor_out[82][18][17] + xor_out[83][18][17] + xor_out[84][18][17];
assign sum_out[17][18][17] = xor_out[85][18][17] + xor_out[86][18][17] + xor_out[87][18][17] + xor_out[88][18][17] + xor_out[89][18][17];
assign sum_out[18][18][17] = xor_out[90][18][17] + xor_out[91][18][17] + xor_out[92][18][17] + xor_out[93][18][17] + xor_out[94][18][17];
assign sum_out[19][18][17] = xor_out[95][18][17] + xor_out[96][18][17] + xor_out[97][18][17] + xor_out[98][18][17] + xor_out[99][18][17];

assign sum_out[0][18][18] = xor_out[0][18][18] + xor_out[1][18][18] + xor_out[2][18][18] + xor_out[3][18][18] + xor_out[4][18][18];
assign sum_out[1][18][18] = xor_out[5][18][18] + xor_out[6][18][18] + xor_out[7][18][18] + xor_out[8][18][18] + xor_out[9][18][18];
assign sum_out[2][18][18] = xor_out[10][18][18] + xor_out[11][18][18] + xor_out[12][18][18] + xor_out[13][18][18] + xor_out[14][18][18];
assign sum_out[3][18][18] = xor_out[15][18][18] + xor_out[16][18][18] + xor_out[17][18][18] + xor_out[18][18][18] + xor_out[19][18][18];
assign sum_out[4][18][18] = xor_out[20][18][18] + xor_out[21][18][18] + xor_out[22][18][18] + xor_out[23][18][18] + xor_out[24][18][18];
assign sum_out[5][18][18] = xor_out[25][18][18] + xor_out[26][18][18] + xor_out[27][18][18] + xor_out[28][18][18] + xor_out[29][18][18];
assign sum_out[6][18][18] = xor_out[30][18][18] + xor_out[31][18][18] + xor_out[32][18][18] + xor_out[33][18][18] + xor_out[34][18][18];
assign sum_out[7][18][18] = xor_out[35][18][18] + xor_out[36][18][18] + xor_out[37][18][18] + xor_out[38][18][18] + xor_out[39][18][18];
assign sum_out[8][18][18] = xor_out[40][18][18] + xor_out[41][18][18] + xor_out[42][18][18] + xor_out[43][18][18] + xor_out[44][18][18];
assign sum_out[9][18][18] = xor_out[45][18][18] + xor_out[46][18][18] + xor_out[47][18][18] + xor_out[48][18][18] + xor_out[49][18][18];
assign sum_out[10][18][18] = xor_out[50][18][18] + xor_out[51][18][18] + xor_out[52][18][18] + xor_out[53][18][18] + xor_out[54][18][18];
assign sum_out[11][18][18] = xor_out[55][18][18] + xor_out[56][18][18] + xor_out[57][18][18] + xor_out[58][18][18] + xor_out[59][18][18];
assign sum_out[12][18][18] = xor_out[60][18][18] + xor_out[61][18][18] + xor_out[62][18][18] + xor_out[63][18][18] + xor_out[64][18][18];
assign sum_out[13][18][18] = xor_out[65][18][18] + xor_out[66][18][18] + xor_out[67][18][18] + xor_out[68][18][18] + xor_out[69][18][18];
assign sum_out[14][18][18] = xor_out[70][18][18] + xor_out[71][18][18] + xor_out[72][18][18] + xor_out[73][18][18] + xor_out[74][18][18];
assign sum_out[15][18][18] = xor_out[75][18][18] + xor_out[76][18][18] + xor_out[77][18][18] + xor_out[78][18][18] + xor_out[79][18][18];
assign sum_out[16][18][18] = xor_out[80][18][18] + xor_out[81][18][18] + xor_out[82][18][18] + xor_out[83][18][18] + xor_out[84][18][18];
assign sum_out[17][18][18] = xor_out[85][18][18] + xor_out[86][18][18] + xor_out[87][18][18] + xor_out[88][18][18] + xor_out[89][18][18];
assign sum_out[18][18][18] = xor_out[90][18][18] + xor_out[91][18][18] + xor_out[92][18][18] + xor_out[93][18][18] + xor_out[94][18][18];
assign sum_out[19][18][18] = xor_out[95][18][18] + xor_out[96][18][18] + xor_out[97][18][18] + xor_out[98][18][18] + xor_out[99][18][18];

assign sum_out[0][18][19] = xor_out[0][18][19] + xor_out[1][18][19] + xor_out[2][18][19] + xor_out[3][18][19] + xor_out[4][18][19];
assign sum_out[1][18][19] = xor_out[5][18][19] + xor_out[6][18][19] + xor_out[7][18][19] + xor_out[8][18][19] + xor_out[9][18][19];
assign sum_out[2][18][19] = xor_out[10][18][19] + xor_out[11][18][19] + xor_out[12][18][19] + xor_out[13][18][19] + xor_out[14][18][19];
assign sum_out[3][18][19] = xor_out[15][18][19] + xor_out[16][18][19] + xor_out[17][18][19] + xor_out[18][18][19] + xor_out[19][18][19];
assign sum_out[4][18][19] = xor_out[20][18][19] + xor_out[21][18][19] + xor_out[22][18][19] + xor_out[23][18][19] + xor_out[24][18][19];
assign sum_out[5][18][19] = xor_out[25][18][19] + xor_out[26][18][19] + xor_out[27][18][19] + xor_out[28][18][19] + xor_out[29][18][19];
assign sum_out[6][18][19] = xor_out[30][18][19] + xor_out[31][18][19] + xor_out[32][18][19] + xor_out[33][18][19] + xor_out[34][18][19];
assign sum_out[7][18][19] = xor_out[35][18][19] + xor_out[36][18][19] + xor_out[37][18][19] + xor_out[38][18][19] + xor_out[39][18][19];
assign sum_out[8][18][19] = xor_out[40][18][19] + xor_out[41][18][19] + xor_out[42][18][19] + xor_out[43][18][19] + xor_out[44][18][19];
assign sum_out[9][18][19] = xor_out[45][18][19] + xor_out[46][18][19] + xor_out[47][18][19] + xor_out[48][18][19] + xor_out[49][18][19];
assign sum_out[10][18][19] = xor_out[50][18][19] + xor_out[51][18][19] + xor_out[52][18][19] + xor_out[53][18][19] + xor_out[54][18][19];
assign sum_out[11][18][19] = xor_out[55][18][19] + xor_out[56][18][19] + xor_out[57][18][19] + xor_out[58][18][19] + xor_out[59][18][19];
assign sum_out[12][18][19] = xor_out[60][18][19] + xor_out[61][18][19] + xor_out[62][18][19] + xor_out[63][18][19] + xor_out[64][18][19];
assign sum_out[13][18][19] = xor_out[65][18][19] + xor_out[66][18][19] + xor_out[67][18][19] + xor_out[68][18][19] + xor_out[69][18][19];
assign sum_out[14][18][19] = xor_out[70][18][19] + xor_out[71][18][19] + xor_out[72][18][19] + xor_out[73][18][19] + xor_out[74][18][19];
assign sum_out[15][18][19] = xor_out[75][18][19] + xor_out[76][18][19] + xor_out[77][18][19] + xor_out[78][18][19] + xor_out[79][18][19];
assign sum_out[16][18][19] = xor_out[80][18][19] + xor_out[81][18][19] + xor_out[82][18][19] + xor_out[83][18][19] + xor_out[84][18][19];
assign sum_out[17][18][19] = xor_out[85][18][19] + xor_out[86][18][19] + xor_out[87][18][19] + xor_out[88][18][19] + xor_out[89][18][19];
assign sum_out[18][18][19] = xor_out[90][18][19] + xor_out[91][18][19] + xor_out[92][18][19] + xor_out[93][18][19] + xor_out[94][18][19];
assign sum_out[19][18][19] = xor_out[95][18][19] + xor_out[96][18][19] + xor_out[97][18][19] + xor_out[98][18][19] + xor_out[99][18][19];

assign sum_out[0][18][20] = xor_out[0][18][20] + xor_out[1][18][20] + xor_out[2][18][20] + xor_out[3][18][20] + xor_out[4][18][20];
assign sum_out[1][18][20] = xor_out[5][18][20] + xor_out[6][18][20] + xor_out[7][18][20] + xor_out[8][18][20] + xor_out[9][18][20];
assign sum_out[2][18][20] = xor_out[10][18][20] + xor_out[11][18][20] + xor_out[12][18][20] + xor_out[13][18][20] + xor_out[14][18][20];
assign sum_out[3][18][20] = xor_out[15][18][20] + xor_out[16][18][20] + xor_out[17][18][20] + xor_out[18][18][20] + xor_out[19][18][20];
assign sum_out[4][18][20] = xor_out[20][18][20] + xor_out[21][18][20] + xor_out[22][18][20] + xor_out[23][18][20] + xor_out[24][18][20];
assign sum_out[5][18][20] = xor_out[25][18][20] + xor_out[26][18][20] + xor_out[27][18][20] + xor_out[28][18][20] + xor_out[29][18][20];
assign sum_out[6][18][20] = xor_out[30][18][20] + xor_out[31][18][20] + xor_out[32][18][20] + xor_out[33][18][20] + xor_out[34][18][20];
assign sum_out[7][18][20] = xor_out[35][18][20] + xor_out[36][18][20] + xor_out[37][18][20] + xor_out[38][18][20] + xor_out[39][18][20];
assign sum_out[8][18][20] = xor_out[40][18][20] + xor_out[41][18][20] + xor_out[42][18][20] + xor_out[43][18][20] + xor_out[44][18][20];
assign sum_out[9][18][20] = xor_out[45][18][20] + xor_out[46][18][20] + xor_out[47][18][20] + xor_out[48][18][20] + xor_out[49][18][20];
assign sum_out[10][18][20] = xor_out[50][18][20] + xor_out[51][18][20] + xor_out[52][18][20] + xor_out[53][18][20] + xor_out[54][18][20];
assign sum_out[11][18][20] = xor_out[55][18][20] + xor_out[56][18][20] + xor_out[57][18][20] + xor_out[58][18][20] + xor_out[59][18][20];
assign sum_out[12][18][20] = xor_out[60][18][20] + xor_out[61][18][20] + xor_out[62][18][20] + xor_out[63][18][20] + xor_out[64][18][20];
assign sum_out[13][18][20] = xor_out[65][18][20] + xor_out[66][18][20] + xor_out[67][18][20] + xor_out[68][18][20] + xor_out[69][18][20];
assign sum_out[14][18][20] = xor_out[70][18][20] + xor_out[71][18][20] + xor_out[72][18][20] + xor_out[73][18][20] + xor_out[74][18][20];
assign sum_out[15][18][20] = xor_out[75][18][20] + xor_out[76][18][20] + xor_out[77][18][20] + xor_out[78][18][20] + xor_out[79][18][20];
assign sum_out[16][18][20] = xor_out[80][18][20] + xor_out[81][18][20] + xor_out[82][18][20] + xor_out[83][18][20] + xor_out[84][18][20];
assign sum_out[17][18][20] = xor_out[85][18][20] + xor_out[86][18][20] + xor_out[87][18][20] + xor_out[88][18][20] + xor_out[89][18][20];
assign sum_out[18][18][20] = xor_out[90][18][20] + xor_out[91][18][20] + xor_out[92][18][20] + xor_out[93][18][20] + xor_out[94][18][20];
assign sum_out[19][18][20] = xor_out[95][18][20] + xor_out[96][18][20] + xor_out[97][18][20] + xor_out[98][18][20] + xor_out[99][18][20];

assign sum_out[0][18][21] = xor_out[0][18][21] + xor_out[1][18][21] + xor_out[2][18][21] + xor_out[3][18][21] + xor_out[4][18][21];
assign sum_out[1][18][21] = xor_out[5][18][21] + xor_out[6][18][21] + xor_out[7][18][21] + xor_out[8][18][21] + xor_out[9][18][21];
assign sum_out[2][18][21] = xor_out[10][18][21] + xor_out[11][18][21] + xor_out[12][18][21] + xor_out[13][18][21] + xor_out[14][18][21];
assign sum_out[3][18][21] = xor_out[15][18][21] + xor_out[16][18][21] + xor_out[17][18][21] + xor_out[18][18][21] + xor_out[19][18][21];
assign sum_out[4][18][21] = xor_out[20][18][21] + xor_out[21][18][21] + xor_out[22][18][21] + xor_out[23][18][21] + xor_out[24][18][21];
assign sum_out[5][18][21] = xor_out[25][18][21] + xor_out[26][18][21] + xor_out[27][18][21] + xor_out[28][18][21] + xor_out[29][18][21];
assign sum_out[6][18][21] = xor_out[30][18][21] + xor_out[31][18][21] + xor_out[32][18][21] + xor_out[33][18][21] + xor_out[34][18][21];
assign sum_out[7][18][21] = xor_out[35][18][21] + xor_out[36][18][21] + xor_out[37][18][21] + xor_out[38][18][21] + xor_out[39][18][21];
assign sum_out[8][18][21] = xor_out[40][18][21] + xor_out[41][18][21] + xor_out[42][18][21] + xor_out[43][18][21] + xor_out[44][18][21];
assign sum_out[9][18][21] = xor_out[45][18][21] + xor_out[46][18][21] + xor_out[47][18][21] + xor_out[48][18][21] + xor_out[49][18][21];
assign sum_out[10][18][21] = xor_out[50][18][21] + xor_out[51][18][21] + xor_out[52][18][21] + xor_out[53][18][21] + xor_out[54][18][21];
assign sum_out[11][18][21] = xor_out[55][18][21] + xor_out[56][18][21] + xor_out[57][18][21] + xor_out[58][18][21] + xor_out[59][18][21];
assign sum_out[12][18][21] = xor_out[60][18][21] + xor_out[61][18][21] + xor_out[62][18][21] + xor_out[63][18][21] + xor_out[64][18][21];
assign sum_out[13][18][21] = xor_out[65][18][21] + xor_out[66][18][21] + xor_out[67][18][21] + xor_out[68][18][21] + xor_out[69][18][21];
assign sum_out[14][18][21] = xor_out[70][18][21] + xor_out[71][18][21] + xor_out[72][18][21] + xor_out[73][18][21] + xor_out[74][18][21];
assign sum_out[15][18][21] = xor_out[75][18][21] + xor_out[76][18][21] + xor_out[77][18][21] + xor_out[78][18][21] + xor_out[79][18][21];
assign sum_out[16][18][21] = xor_out[80][18][21] + xor_out[81][18][21] + xor_out[82][18][21] + xor_out[83][18][21] + xor_out[84][18][21];
assign sum_out[17][18][21] = xor_out[85][18][21] + xor_out[86][18][21] + xor_out[87][18][21] + xor_out[88][18][21] + xor_out[89][18][21];
assign sum_out[18][18][21] = xor_out[90][18][21] + xor_out[91][18][21] + xor_out[92][18][21] + xor_out[93][18][21] + xor_out[94][18][21];
assign sum_out[19][18][21] = xor_out[95][18][21] + xor_out[96][18][21] + xor_out[97][18][21] + xor_out[98][18][21] + xor_out[99][18][21];

assign sum_out[0][18][22] = xor_out[0][18][22] + xor_out[1][18][22] + xor_out[2][18][22] + xor_out[3][18][22] + xor_out[4][18][22];
assign sum_out[1][18][22] = xor_out[5][18][22] + xor_out[6][18][22] + xor_out[7][18][22] + xor_out[8][18][22] + xor_out[9][18][22];
assign sum_out[2][18][22] = xor_out[10][18][22] + xor_out[11][18][22] + xor_out[12][18][22] + xor_out[13][18][22] + xor_out[14][18][22];
assign sum_out[3][18][22] = xor_out[15][18][22] + xor_out[16][18][22] + xor_out[17][18][22] + xor_out[18][18][22] + xor_out[19][18][22];
assign sum_out[4][18][22] = xor_out[20][18][22] + xor_out[21][18][22] + xor_out[22][18][22] + xor_out[23][18][22] + xor_out[24][18][22];
assign sum_out[5][18][22] = xor_out[25][18][22] + xor_out[26][18][22] + xor_out[27][18][22] + xor_out[28][18][22] + xor_out[29][18][22];
assign sum_out[6][18][22] = xor_out[30][18][22] + xor_out[31][18][22] + xor_out[32][18][22] + xor_out[33][18][22] + xor_out[34][18][22];
assign sum_out[7][18][22] = xor_out[35][18][22] + xor_out[36][18][22] + xor_out[37][18][22] + xor_out[38][18][22] + xor_out[39][18][22];
assign sum_out[8][18][22] = xor_out[40][18][22] + xor_out[41][18][22] + xor_out[42][18][22] + xor_out[43][18][22] + xor_out[44][18][22];
assign sum_out[9][18][22] = xor_out[45][18][22] + xor_out[46][18][22] + xor_out[47][18][22] + xor_out[48][18][22] + xor_out[49][18][22];
assign sum_out[10][18][22] = xor_out[50][18][22] + xor_out[51][18][22] + xor_out[52][18][22] + xor_out[53][18][22] + xor_out[54][18][22];
assign sum_out[11][18][22] = xor_out[55][18][22] + xor_out[56][18][22] + xor_out[57][18][22] + xor_out[58][18][22] + xor_out[59][18][22];
assign sum_out[12][18][22] = xor_out[60][18][22] + xor_out[61][18][22] + xor_out[62][18][22] + xor_out[63][18][22] + xor_out[64][18][22];
assign sum_out[13][18][22] = xor_out[65][18][22] + xor_out[66][18][22] + xor_out[67][18][22] + xor_out[68][18][22] + xor_out[69][18][22];
assign sum_out[14][18][22] = xor_out[70][18][22] + xor_out[71][18][22] + xor_out[72][18][22] + xor_out[73][18][22] + xor_out[74][18][22];
assign sum_out[15][18][22] = xor_out[75][18][22] + xor_out[76][18][22] + xor_out[77][18][22] + xor_out[78][18][22] + xor_out[79][18][22];
assign sum_out[16][18][22] = xor_out[80][18][22] + xor_out[81][18][22] + xor_out[82][18][22] + xor_out[83][18][22] + xor_out[84][18][22];
assign sum_out[17][18][22] = xor_out[85][18][22] + xor_out[86][18][22] + xor_out[87][18][22] + xor_out[88][18][22] + xor_out[89][18][22];
assign sum_out[18][18][22] = xor_out[90][18][22] + xor_out[91][18][22] + xor_out[92][18][22] + xor_out[93][18][22] + xor_out[94][18][22];
assign sum_out[19][18][22] = xor_out[95][18][22] + xor_out[96][18][22] + xor_out[97][18][22] + xor_out[98][18][22] + xor_out[99][18][22];

assign sum_out[0][18][23] = xor_out[0][18][23] + xor_out[1][18][23] + xor_out[2][18][23] + xor_out[3][18][23] + xor_out[4][18][23];
assign sum_out[1][18][23] = xor_out[5][18][23] + xor_out[6][18][23] + xor_out[7][18][23] + xor_out[8][18][23] + xor_out[9][18][23];
assign sum_out[2][18][23] = xor_out[10][18][23] + xor_out[11][18][23] + xor_out[12][18][23] + xor_out[13][18][23] + xor_out[14][18][23];
assign sum_out[3][18][23] = xor_out[15][18][23] + xor_out[16][18][23] + xor_out[17][18][23] + xor_out[18][18][23] + xor_out[19][18][23];
assign sum_out[4][18][23] = xor_out[20][18][23] + xor_out[21][18][23] + xor_out[22][18][23] + xor_out[23][18][23] + xor_out[24][18][23];
assign sum_out[5][18][23] = xor_out[25][18][23] + xor_out[26][18][23] + xor_out[27][18][23] + xor_out[28][18][23] + xor_out[29][18][23];
assign sum_out[6][18][23] = xor_out[30][18][23] + xor_out[31][18][23] + xor_out[32][18][23] + xor_out[33][18][23] + xor_out[34][18][23];
assign sum_out[7][18][23] = xor_out[35][18][23] + xor_out[36][18][23] + xor_out[37][18][23] + xor_out[38][18][23] + xor_out[39][18][23];
assign sum_out[8][18][23] = xor_out[40][18][23] + xor_out[41][18][23] + xor_out[42][18][23] + xor_out[43][18][23] + xor_out[44][18][23];
assign sum_out[9][18][23] = xor_out[45][18][23] + xor_out[46][18][23] + xor_out[47][18][23] + xor_out[48][18][23] + xor_out[49][18][23];
assign sum_out[10][18][23] = xor_out[50][18][23] + xor_out[51][18][23] + xor_out[52][18][23] + xor_out[53][18][23] + xor_out[54][18][23];
assign sum_out[11][18][23] = xor_out[55][18][23] + xor_out[56][18][23] + xor_out[57][18][23] + xor_out[58][18][23] + xor_out[59][18][23];
assign sum_out[12][18][23] = xor_out[60][18][23] + xor_out[61][18][23] + xor_out[62][18][23] + xor_out[63][18][23] + xor_out[64][18][23];
assign sum_out[13][18][23] = xor_out[65][18][23] + xor_out[66][18][23] + xor_out[67][18][23] + xor_out[68][18][23] + xor_out[69][18][23];
assign sum_out[14][18][23] = xor_out[70][18][23] + xor_out[71][18][23] + xor_out[72][18][23] + xor_out[73][18][23] + xor_out[74][18][23];
assign sum_out[15][18][23] = xor_out[75][18][23] + xor_out[76][18][23] + xor_out[77][18][23] + xor_out[78][18][23] + xor_out[79][18][23];
assign sum_out[16][18][23] = xor_out[80][18][23] + xor_out[81][18][23] + xor_out[82][18][23] + xor_out[83][18][23] + xor_out[84][18][23];
assign sum_out[17][18][23] = xor_out[85][18][23] + xor_out[86][18][23] + xor_out[87][18][23] + xor_out[88][18][23] + xor_out[89][18][23];
assign sum_out[18][18][23] = xor_out[90][18][23] + xor_out[91][18][23] + xor_out[92][18][23] + xor_out[93][18][23] + xor_out[94][18][23];
assign sum_out[19][18][23] = xor_out[95][18][23] + xor_out[96][18][23] + xor_out[97][18][23] + xor_out[98][18][23] + xor_out[99][18][23];

assign sum_out[0][19][0] = xor_out[0][19][0] + xor_out[1][19][0] + xor_out[2][19][0] + xor_out[3][19][0] + xor_out[4][19][0];
assign sum_out[1][19][0] = xor_out[5][19][0] + xor_out[6][19][0] + xor_out[7][19][0] + xor_out[8][19][0] + xor_out[9][19][0];
assign sum_out[2][19][0] = xor_out[10][19][0] + xor_out[11][19][0] + xor_out[12][19][0] + xor_out[13][19][0] + xor_out[14][19][0];
assign sum_out[3][19][0] = xor_out[15][19][0] + xor_out[16][19][0] + xor_out[17][19][0] + xor_out[18][19][0] + xor_out[19][19][0];
assign sum_out[4][19][0] = xor_out[20][19][0] + xor_out[21][19][0] + xor_out[22][19][0] + xor_out[23][19][0] + xor_out[24][19][0];
assign sum_out[5][19][0] = xor_out[25][19][0] + xor_out[26][19][0] + xor_out[27][19][0] + xor_out[28][19][0] + xor_out[29][19][0];
assign sum_out[6][19][0] = xor_out[30][19][0] + xor_out[31][19][0] + xor_out[32][19][0] + xor_out[33][19][0] + xor_out[34][19][0];
assign sum_out[7][19][0] = xor_out[35][19][0] + xor_out[36][19][0] + xor_out[37][19][0] + xor_out[38][19][0] + xor_out[39][19][0];
assign sum_out[8][19][0] = xor_out[40][19][0] + xor_out[41][19][0] + xor_out[42][19][0] + xor_out[43][19][0] + xor_out[44][19][0];
assign sum_out[9][19][0] = xor_out[45][19][0] + xor_out[46][19][0] + xor_out[47][19][0] + xor_out[48][19][0] + xor_out[49][19][0];
assign sum_out[10][19][0] = xor_out[50][19][0] + xor_out[51][19][0] + xor_out[52][19][0] + xor_out[53][19][0] + xor_out[54][19][0];
assign sum_out[11][19][0] = xor_out[55][19][0] + xor_out[56][19][0] + xor_out[57][19][0] + xor_out[58][19][0] + xor_out[59][19][0];
assign sum_out[12][19][0] = xor_out[60][19][0] + xor_out[61][19][0] + xor_out[62][19][0] + xor_out[63][19][0] + xor_out[64][19][0];
assign sum_out[13][19][0] = xor_out[65][19][0] + xor_out[66][19][0] + xor_out[67][19][0] + xor_out[68][19][0] + xor_out[69][19][0];
assign sum_out[14][19][0] = xor_out[70][19][0] + xor_out[71][19][0] + xor_out[72][19][0] + xor_out[73][19][0] + xor_out[74][19][0];
assign sum_out[15][19][0] = xor_out[75][19][0] + xor_out[76][19][0] + xor_out[77][19][0] + xor_out[78][19][0] + xor_out[79][19][0];
assign sum_out[16][19][0] = xor_out[80][19][0] + xor_out[81][19][0] + xor_out[82][19][0] + xor_out[83][19][0] + xor_out[84][19][0];
assign sum_out[17][19][0] = xor_out[85][19][0] + xor_out[86][19][0] + xor_out[87][19][0] + xor_out[88][19][0] + xor_out[89][19][0];
assign sum_out[18][19][0] = xor_out[90][19][0] + xor_out[91][19][0] + xor_out[92][19][0] + xor_out[93][19][0] + xor_out[94][19][0];
assign sum_out[19][19][0] = xor_out[95][19][0] + xor_out[96][19][0] + xor_out[97][19][0] + xor_out[98][19][0] + xor_out[99][19][0];

assign sum_out[0][19][1] = xor_out[0][19][1] + xor_out[1][19][1] + xor_out[2][19][1] + xor_out[3][19][1] + xor_out[4][19][1];
assign sum_out[1][19][1] = xor_out[5][19][1] + xor_out[6][19][1] + xor_out[7][19][1] + xor_out[8][19][1] + xor_out[9][19][1];
assign sum_out[2][19][1] = xor_out[10][19][1] + xor_out[11][19][1] + xor_out[12][19][1] + xor_out[13][19][1] + xor_out[14][19][1];
assign sum_out[3][19][1] = xor_out[15][19][1] + xor_out[16][19][1] + xor_out[17][19][1] + xor_out[18][19][1] + xor_out[19][19][1];
assign sum_out[4][19][1] = xor_out[20][19][1] + xor_out[21][19][1] + xor_out[22][19][1] + xor_out[23][19][1] + xor_out[24][19][1];
assign sum_out[5][19][1] = xor_out[25][19][1] + xor_out[26][19][1] + xor_out[27][19][1] + xor_out[28][19][1] + xor_out[29][19][1];
assign sum_out[6][19][1] = xor_out[30][19][1] + xor_out[31][19][1] + xor_out[32][19][1] + xor_out[33][19][1] + xor_out[34][19][1];
assign sum_out[7][19][1] = xor_out[35][19][1] + xor_out[36][19][1] + xor_out[37][19][1] + xor_out[38][19][1] + xor_out[39][19][1];
assign sum_out[8][19][1] = xor_out[40][19][1] + xor_out[41][19][1] + xor_out[42][19][1] + xor_out[43][19][1] + xor_out[44][19][1];
assign sum_out[9][19][1] = xor_out[45][19][1] + xor_out[46][19][1] + xor_out[47][19][1] + xor_out[48][19][1] + xor_out[49][19][1];
assign sum_out[10][19][1] = xor_out[50][19][1] + xor_out[51][19][1] + xor_out[52][19][1] + xor_out[53][19][1] + xor_out[54][19][1];
assign sum_out[11][19][1] = xor_out[55][19][1] + xor_out[56][19][1] + xor_out[57][19][1] + xor_out[58][19][1] + xor_out[59][19][1];
assign sum_out[12][19][1] = xor_out[60][19][1] + xor_out[61][19][1] + xor_out[62][19][1] + xor_out[63][19][1] + xor_out[64][19][1];
assign sum_out[13][19][1] = xor_out[65][19][1] + xor_out[66][19][1] + xor_out[67][19][1] + xor_out[68][19][1] + xor_out[69][19][1];
assign sum_out[14][19][1] = xor_out[70][19][1] + xor_out[71][19][1] + xor_out[72][19][1] + xor_out[73][19][1] + xor_out[74][19][1];
assign sum_out[15][19][1] = xor_out[75][19][1] + xor_out[76][19][1] + xor_out[77][19][1] + xor_out[78][19][1] + xor_out[79][19][1];
assign sum_out[16][19][1] = xor_out[80][19][1] + xor_out[81][19][1] + xor_out[82][19][1] + xor_out[83][19][1] + xor_out[84][19][1];
assign sum_out[17][19][1] = xor_out[85][19][1] + xor_out[86][19][1] + xor_out[87][19][1] + xor_out[88][19][1] + xor_out[89][19][1];
assign sum_out[18][19][1] = xor_out[90][19][1] + xor_out[91][19][1] + xor_out[92][19][1] + xor_out[93][19][1] + xor_out[94][19][1];
assign sum_out[19][19][1] = xor_out[95][19][1] + xor_out[96][19][1] + xor_out[97][19][1] + xor_out[98][19][1] + xor_out[99][19][1];

assign sum_out[0][19][2] = xor_out[0][19][2] + xor_out[1][19][2] + xor_out[2][19][2] + xor_out[3][19][2] + xor_out[4][19][2];
assign sum_out[1][19][2] = xor_out[5][19][2] + xor_out[6][19][2] + xor_out[7][19][2] + xor_out[8][19][2] + xor_out[9][19][2];
assign sum_out[2][19][2] = xor_out[10][19][2] + xor_out[11][19][2] + xor_out[12][19][2] + xor_out[13][19][2] + xor_out[14][19][2];
assign sum_out[3][19][2] = xor_out[15][19][2] + xor_out[16][19][2] + xor_out[17][19][2] + xor_out[18][19][2] + xor_out[19][19][2];
assign sum_out[4][19][2] = xor_out[20][19][2] + xor_out[21][19][2] + xor_out[22][19][2] + xor_out[23][19][2] + xor_out[24][19][2];
assign sum_out[5][19][2] = xor_out[25][19][2] + xor_out[26][19][2] + xor_out[27][19][2] + xor_out[28][19][2] + xor_out[29][19][2];
assign sum_out[6][19][2] = xor_out[30][19][2] + xor_out[31][19][2] + xor_out[32][19][2] + xor_out[33][19][2] + xor_out[34][19][2];
assign sum_out[7][19][2] = xor_out[35][19][2] + xor_out[36][19][2] + xor_out[37][19][2] + xor_out[38][19][2] + xor_out[39][19][2];
assign sum_out[8][19][2] = xor_out[40][19][2] + xor_out[41][19][2] + xor_out[42][19][2] + xor_out[43][19][2] + xor_out[44][19][2];
assign sum_out[9][19][2] = xor_out[45][19][2] + xor_out[46][19][2] + xor_out[47][19][2] + xor_out[48][19][2] + xor_out[49][19][2];
assign sum_out[10][19][2] = xor_out[50][19][2] + xor_out[51][19][2] + xor_out[52][19][2] + xor_out[53][19][2] + xor_out[54][19][2];
assign sum_out[11][19][2] = xor_out[55][19][2] + xor_out[56][19][2] + xor_out[57][19][2] + xor_out[58][19][2] + xor_out[59][19][2];
assign sum_out[12][19][2] = xor_out[60][19][2] + xor_out[61][19][2] + xor_out[62][19][2] + xor_out[63][19][2] + xor_out[64][19][2];
assign sum_out[13][19][2] = xor_out[65][19][2] + xor_out[66][19][2] + xor_out[67][19][2] + xor_out[68][19][2] + xor_out[69][19][2];
assign sum_out[14][19][2] = xor_out[70][19][2] + xor_out[71][19][2] + xor_out[72][19][2] + xor_out[73][19][2] + xor_out[74][19][2];
assign sum_out[15][19][2] = xor_out[75][19][2] + xor_out[76][19][2] + xor_out[77][19][2] + xor_out[78][19][2] + xor_out[79][19][2];
assign sum_out[16][19][2] = xor_out[80][19][2] + xor_out[81][19][2] + xor_out[82][19][2] + xor_out[83][19][2] + xor_out[84][19][2];
assign sum_out[17][19][2] = xor_out[85][19][2] + xor_out[86][19][2] + xor_out[87][19][2] + xor_out[88][19][2] + xor_out[89][19][2];
assign sum_out[18][19][2] = xor_out[90][19][2] + xor_out[91][19][2] + xor_out[92][19][2] + xor_out[93][19][2] + xor_out[94][19][2];
assign sum_out[19][19][2] = xor_out[95][19][2] + xor_out[96][19][2] + xor_out[97][19][2] + xor_out[98][19][2] + xor_out[99][19][2];

assign sum_out[0][19][3] = xor_out[0][19][3] + xor_out[1][19][3] + xor_out[2][19][3] + xor_out[3][19][3] + xor_out[4][19][3];
assign sum_out[1][19][3] = xor_out[5][19][3] + xor_out[6][19][3] + xor_out[7][19][3] + xor_out[8][19][3] + xor_out[9][19][3];
assign sum_out[2][19][3] = xor_out[10][19][3] + xor_out[11][19][3] + xor_out[12][19][3] + xor_out[13][19][3] + xor_out[14][19][3];
assign sum_out[3][19][3] = xor_out[15][19][3] + xor_out[16][19][3] + xor_out[17][19][3] + xor_out[18][19][3] + xor_out[19][19][3];
assign sum_out[4][19][3] = xor_out[20][19][3] + xor_out[21][19][3] + xor_out[22][19][3] + xor_out[23][19][3] + xor_out[24][19][3];
assign sum_out[5][19][3] = xor_out[25][19][3] + xor_out[26][19][3] + xor_out[27][19][3] + xor_out[28][19][3] + xor_out[29][19][3];
assign sum_out[6][19][3] = xor_out[30][19][3] + xor_out[31][19][3] + xor_out[32][19][3] + xor_out[33][19][3] + xor_out[34][19][3];
assign sum_out[7][19][3] = xor_out[35][19][3] + xor_out[36][19][3] + xor_out[37][19][3] + xor_out[38][19][3] + xor_out[39][19][3];
assign sum_out[8][19][3] = xor_out[40][19][3] + xor_out[41][19][3] + xor_out[42][19][3] + xor_out[43][19][3] + xor_out[44][19][3];
assign sum_out[9][19][3] = xor_out[45][19][3] + xor_out[46][19][3] + xor_out[47][19][3] + xor_out[48][19][3] + xor_out[49][19][3];
assign sum_out[10][19][3] = xor_out[50][19][3] + xor_out[51][19][3] + xor_out[52][19][3] + xor_out[53][19][3] + xor_out[54][19][3];
assign sum_out[11][19][3] = xor_out[55][19][3] + xor_out[56][19][3] + xor_out[57][19][3] + xor_out[58][19][3] + xor_out[59][19][3];
assign sum_out[12][19][3] = xor_out[60][19][3] + xor_out[61][19][3] + xor_out[62][19][3] + xor_out[63][19][3] + xor_out[64][19][3];
assign sum_out[13][19][3] = xor_out[65][19][3] + xor_out[66][19][3] + xor_out[67][19][3] + xor_out[68][19][3] + xor_out[69][19][3];
assign sum_out[14][19][3] = xor_out[70][19][3] + xor_out[71][19][3] + xor_out[72][19][3] + xor_out[73][19][3] + xor_out[74][19][3];
assign sum_out[15][19][3] = xor_out[75][19][3] + xor_out[76][19][3] + xor_out[77][19][3] + xor_out[78][19][3] + xor_out[79][19][3];
assign sum_out[16][19][3] = xor_out[80][19][3] + xor_out[81][19][3] + xor_out[82][19][3] + xor_out[83][19][3] + xor_out[84][19][3];
assign sum_out[17][19][3] = xor_out[85][19][3] + xor_out[86][19][3] + xor_out[87][19][3] + xor_out[88][19][3] + xor_out[89][19][3];
assign sum_out[18][19][3] = xor_out[90][19][3] + xor_out[91][19][3] + xor_out[92][19][3] + xor_out[93][19][3] + xor_out[94][19][3];
assign sum_out[19][19][3] = xor_out[95][19][3] + xor_out[96][19][3] + xor_out[97][19][3] + xor_out[98][19][3] + xor_out[99][19][3];

assign sum_out[0][19][4] = xor_out[0][19][4] + xor_out[1][19][4] + xor_out[2][19][4] + xor_out[3][19][4] + xor_out[4][19][4];
assign sum_out[1][19][4] = xor_out[5][19][4] + xor_out[6][19][4] + xor_out[7][19][4] + xor_out[8][19][4] + xor_out[9][19][4];
assign sum_out[2][19][4] = xor_out[10][19][4] + xor_out[11][19][4] + xor_out[12][19][4] + xor_out[13][19][4] + xor_out[14][19][4];
assign sum_out[3][19][4] = xor_out[15][19][4] + xor_out[16][19][4] + xor_out[17][19][4] + xor_out[18][19][4] + xor_out[19][19][4];
assign sum_out[4][19][4] = xor_out[20][19][4] + xor_out[21][19][4] + xor_out[22][19][4] + xor_out[23][19][4] + xor_out[24][19][4];
assign sum_out[5][19][4] = xor_out[25][19][4] + xor_out[26][19][4] + xor_out[27][19][4] + xor_out[28][19][4] + xor_out[29][19][4];
assign sum_out[6][19][4] = xor_out[30][19][4] + xor_out[31][19][4] + xor_out[32][19][4] + xor_out[33][19][4] + xor_out[34][19][4];
assign sum_out[7][19][4] = xor_out[35][19][4] + xor_out[36][19][4] + xor_out[37][19][4] + xor_out[38][19][4] + xor_out[39][19][4];
assign sum_out[8][19][4] = xor_out[40][19][4] + xor_out[41][19][4] + xor_out[42][19][4] + xor_out[43][19][4] + xor_out[44][19][4];
assign sum_out[9][19][4] = xor_out[45][19][4] + xor_out[46][19][4] + xor_out[47][19][4] + xor_out[48][19][4] + xor_out[49][19][4];
assign sum_out[10][19][4] = xor_out[50][19][4] + xor_out[51][19][4] + xor_out[52][19][4] + xor_out[53][19][4] + xor_out[54][19][4];
assign sum_out[11][19][4] = xor_out[55][19][4] + xor_out[56][19][4] + xor_out[57][19][4] + xor_out[58][19][4] + xor_out[59][19][4];
assign sum_out[12][19][4] = xor_out[60][19][4] + xor_out[61][19][4] + xor_out[62][19][4] + xor_out[63][19][4] + xor_out[64][19][4];
assign sum_out[13][19][4] = xor_out[65][19][4] + xor_out[66][19][4] + xor_out[67][19][4] + xor_out[68][19][4] + xor_out[69][19][4];
assign sum_out[14][19][4] = xor_out[70][19][4] + xor_out[71][19][4] + xor_out[72][19][4] + xor_out[73][19][4] + xor_out[74][19][4];
assign sum_out[15][19][4] = xor_out[75][19][4] + xor_out[76][19][4] + xor_out[77][19][4] + xor_out[78][19][4] + xor_out[79][19][4];
assign sum_out[16][19][4] = xor_out[80][19][4] + xor_out[81][19][4] + xor_out[82][19][4] + xor_out[83][19][4] + xor_out[84][19][4];
assign sum_out[17][19][4] = xor_out[85][19][4] + xor_out[86][19][4] + xor_out[87][19][4] + xor_out[88][19][4] + xor_out[89][19][4];
assign sum_out[18][19][4] = xor_out[90][19][4] + xor_out[91][19][4] + xor_out[92][19][4] + xor_out[93][19][4] + xor_out[94][19][4];
assign sum_out[19][19][4] = xor_out[95][19][4] + xor_out[96][19][4] + xor_out[97][19][4] + xor_out[98][19][4] + xor_out[99][19][4];

assign sum_out[0][19][5] = xor_out[0][19][5] + xor_out[1][19][5] + xor_out[2][19][5] + xor_out[3][19][5] + xor_out[4][19][5];
assign sum_out[1][19][5] = xor_out[5][19][5] + xor_out[6][19][5] + xor_out[7][19][5] + xor_out[8][19][5] + xor_out[9][19][5];
assign sum_out[2][19][5] = xor_out[10][19][5] + xor_out[11][19][5] + xor_out[12][19][5] + xor_out[13][19][5] + xor_out[14][19][5];
assign sum_out[3][19][5] = xor_out[15][19][5] + xor_out[16][19][5] + xor_out[17][19][5] + xor_out[18][19][5] + xor_out[19][19][5];
assign sum_out[4][19][5] = xor_out[20][19][5] + xor_out[21][19][5] + xor_out[22][19][5] + xor_out[23][19][5] + xor_out[24][19][5];
assign sum_out[5][19][5] = xor_out[25][19][5] + xor_out[26][19][5] + xor_out[27][19][5] + xor_out[28][19][5] + xor_out[29][19][5];
assign sum_out[6][19][5] = xor_out[30][19][5] + xor_out[31][19][5] + xor_out[32][19][5] + xor_out[33][19][5] + xor_out[34][19][5];
assign sum_out[7][19][5] = xor_out[35][19][5] + xor_out[36][19][5] + xor_out[37][19][5] + xor_out[38][19][5] + xor_out[39][19][5];
assign sum_out[8][19][5] = xor_out[40][19][5] + xor_out[41][19][5] + xor_out[42][19][5] + xor_out[43][19][5] + xor_out[44][19][5];
assign sum_out[9][19][5] = xor_out[45][19][5] + xor_out[46][19][5] + xor_out[47][19][5] + xor_out[48][19][5] + xor_out[49][19][5];
assign sum_out[10][19][5] = xor_out[50][19][5] + xor_out[51][19][5] + xor_out[52][19][5] + xor_out[53][19][5] + xor_out[54][19][5];
assign sum_out[11][19][5] = xor_out[55][19][5] + xor_out[56][19][5] + xor_out[57][19][5] + xor_out[58][19][5] + xor_out[59][19][5];
assign sum_out[12][19][5] = xor_out[60][19][5] + xor_out[61][19][5] + xor_out[62][19][5] + xor_out[63][19][5] + xor_out[64][19][5];
assign sum_out[13][19][5] = xor_out[65][19][5] + xor_out[66][19][5] + xor_out[67][19][5] + xor_out[68][19][5] + xor_out[69][19][5];
assign sum_out[14][19][5] = xor_out[70][19][5] + xor_out[71][19][5] + xor_out[72][19][5] + xor_out[73][19][5] + xor_out[74][19][5];
assign sum_out[15][19][5] = xor_out[75][19][5] + xor_out[76][19][5] + xor_out[77][19][5] + xor_out[78][19][5] + xor_out[79][19][5];
assign sum_out[16][19][5] = xor_out[80][19][5] + xor_out[81][19][5] + xor_out[82][19][5] + xor_out[83][19][5] + xor_out[84][19][5];
assign sum_out[17][19][5] = xor_out[85][19][5] + xor_out[86][19][5] + xor_out[87][19][5] + xor_out[88][19][5] + xor_out[89][19][5];
assign sum_out[18][19][5] = xor_out[90][19][5] + xor_out[91][19][5] + xor_out[92][19][5] + xor_out[93][19][5] + xor_out[94][19][5];
assign sum_out[19][19][5] = xor_out[95][19][5] + xor_out[96][19][5] + xor_out[97][19][5] + xor_out[98][19][5] + xor_out[99][19][5];

assign sum_out[0][19][6] = xor_out[0][19][6] + xor_out[1][19][6] + xor_out[2][19][6] + xor_out[3][19][6] + xor_out[4][19][6];
assign sum_out[1][19][6] = xor_out[5][19][6] + xor_out[6][19][6] + xor_out[7][19][6] + xor_out[8][19][6] + xor_out[9][19][6];
assign sum_out[2][19][6] = xor_out[10][19][6] + xor_out[11][19][6] + xor_out[12][19][6] + xor_out[13][19][6] + xor_out[14][19][6];
assign sum_out[3][19][6] = xor_out[15][19][6] + xor_out[16][19][6] + xor_out[17][19][6] + xor_out[18][19][6] + xor_out[19][19][6];
assign sum_out[4][19][6] = xor_out[20][19][6] + xor_out[21][19][6] + xor_out[22][19][6] + xor_out[23][19][6] + xor_out[24][19][6];
assign sum_out[5][19][6] = xor_out[25][19][6] + xor_out[26][19][6] + xor_out[27][19][6] + xor_out[28][19][6] + xor_out[29][19][6];
assign sum_out[6][19][6] = xor_out[30][19][6] + xor_out[31][19][6] + xor_out[32][19][6] + xor_out[33][19][6] + xor_out[34][19][6];
assign sum_out[7][19][6] = xor_out[35][19][6] + xor_out[36][19][6] + xor_out[37][19][6] + xor_out[38][19][6] + xor_out[39][19][6];
assign sum_out[8][19][6] = xor_out[40][19][6] + xor_out[41][19][6] + xor_out[42][19][6] + xor_out[43][19][6] + xor_out[44][19][6];
assign sum_out[9][19][6] = xor_out[45][19][6] + xor_out[46][19][6] + xor_out[47][19][6] + xor_out[48][19][6] + xor_out[49][19][6];
assign sum_out[10][19][6] = xor_out[50][19][6] + xor_out[51][19][6] + xor_out[52][19][6] + xor_out[53][19][6] + xor_out[54][19][6];
assign sum_out[11][19][6] = xor_out[55][19][6] + xor_out[56][19][6] + xor_out[57][19][6] + xor_out[58][19][6] + xor_out[59][19][6];
assign sum_out[12][19][6] = xor_out[60][19][6] + xor_out[61][19][6] + xor_out[62][19][6] + xor_out[63][19][6] + xor_out[64][19][6];
assign sum_out[13][19][6] = xor_out[65][19][6] + xor_out[66][19][6] + xor_out[67][19][6] + xor_out[68][19][6] + xor_out[69][19][6];
assign sum_out[14][19][6] = xor_out[70][19][6] + xor_out[71][19][6] + xor_out[72][19][6] + xor_out[73][19][6] + xor_out[74][19][6];
assign sum_out[15][19][6] = xor_out[75][19][6] + xor_out[76][19][6] + xor_out[77][19][6] + xor_out[78][19][6] + xor_out[79][19][6];
assign sum_out[16][19][6] = xor_out[80][19][6] + xor_out[81][19][6] + xor_out[82][19][6] + xor_out[83][19][6] + xor_out[84][19][6];
assign sum_out[17][19][6] = xor_out[85][19][6] + xor_out[86][19][6] + xor_out[87][19][6] + xor_out[88][19][6] + xor_out[89][19][6];
assign sum_out[18][19][6] = xor_out[90][19][6] + xor_out[91][19][6] + xor_out[92][19][6] + xor_out[93][19][6] + xor_out[94][19][6];
assign sum_out[19][19][6] = xor_out[95][19][6] + xor_out[96][19][6] + xor_out[97][19][6] + xor_out[98][19][6] + xor_out[99][19][6];

assign sum_out[0][19][7] = xor_out[0][19][7] + xor_out[1][19][7] + xor_out[2][19][7] + xor_out[3][19][7] + xor_out[4][19][7];
assign sum_out[1][19][7] = xor_out[5][19][7] + xor_out[6][19][7] + xor_out[7][19][7] + xor_out[8][19][7] + xor_out[9][19][7];
assign sum_out[2][19][7] = xor_out[10][19][7] + xor_out[11][19][7] + xor_out[12][19][7] + xor_out[13][19][7] + xor_out[14][19][7];
assign sum_out[3][19][7] = xor_out[15][19][7] + xor_out[16][19][7] + xor_out[17][19][7] + xor_out[18][19][7] + xor_out[19][19][7];
assign sum_out[4][19][7] = xor_out[20][19][7] + xor_out[21][19][7] + xor_out[22][19][7] + xor_out[23][19][7] + xor_out[24][19][7];
assign sum_out[5][19][7] = xor_out[25][19][7] + xor_out[26][19][7] + xor_out[27][19][7] + xor_out[28][19][7] + xor_out[29][19][7];
assign sum_out[6][19][7] = xor_out[30][19][7] + xor_out[31][19][7] + xor_out[32][19][7] + xor_out[33][19][7] + xor_out[34][19][7];
assign sum_out[7][19][7] = xor_out[35][19][7] + xor_out[36][19][7] + xor_out[37][19][7] + xor_out[38][19][7] + xor_out[39][19][7];
assign sum_out[8][19][7] = xor_out[40][19][7] + xor_out[41][19][7] + xor_out[42][19][7] + xor_out[43][19][7] + xor_out[44][19][7];
assign sum_out[9][19][7] = xor_out[45][19][7] + xor_out[46][19][7] + xor_out[47][19][7] + xor_out[48][19][7] + xor_out[49][19][7];
assign sum_out[10][19][7] = xor_out[50][19][7] + xor_out[51][19][7] + xor_out[52][19][7] + xor_out[53][19][7] + xor_out[54][19][7];
assign sum_out[11][19][7] = xor_out[55][19][7] + xor_out[56][19][7] + xor_out[57][19][7] + xor_out[58][19][7] + xor_out[59][19][7];
assign sum_out[12][19][7] = xor_out[60][19][7] + xor_out[61][19][7] + xor_out[62][19][7] + xor_out[63][19][7] + xor_out[64][19][7];
assign sum_out[13][19][7] = xor_out[65][19][7] + xor_out[66][19][7] + xor_out[67][19][7] + xor_out[68][19][7] + xor_out[69][19][7];
assign sum_out[14][19][7] = xor_out[70][19][7] + xor_out[71][19][7] + xor_out[72][19][7] + xor_out[73][19][7] + xor_out[74][19][7];
assign sum_out[15][19][7] = xor_out[75][19][7] + xor_out[76][19][7] + xor_out[77][19][7] + xor_out[78][19][7] + xor_out[79][19][7];
assign sum_out[16][19][7] = xor_out[80][19][7] + xor_out[81][19][7] + xor_out[82][19][7] + xor_out[83][19][7] + xor_out[84][19][7];
assign sum_out[17][19][7] = xor_out[85][19][7] + xor_out[86][19][7] + xor_out[87][19][7] + xor_out[88][19][7] + xor_out[89][19][7];
assign sum_out[18][19][7] = xor_out[90][19][7] + xor_out[91][19][7] + xor_out[92][19][7] + xor_out[93][19][7] + xor_out[94][19][7];
assign sum_out[19][19][7] = xor_out[95][19][7] + xor_out[96][19][7] + xor_out[97][19][7] + xor_out[98][19][7] + xor_out[99][19][7];

assign sum_out[0][19][8] = xor_out[0][19][8] + xor_out[1][19][8] + xor_out[2][19][8] + xor_out[3][19][8] + xor_out[4][19][8];
assign sum_out[1][19][8] = xor_out[5][19][8] + xor_out[6][19][8] + xor_out[7][19][8] + xor_out[8][19][8] + xor_out[9][19][8];
assign sum_out[2][19][8] = xor_out[10][19][8] + xor_out[11][19][8] + xor_out[12][19][8] + xor_out[13][19][8] + xor_out[14][19][8];
assign sum_out[3][19][8] = xor_out[15][19][8] + xor_out[16][19][8] + xor_out[17][19][8] + xor_out[18][19][8] + xor_out[19][19][8];
assign sum_out[4][19][8] = xor_out[20][19][8] + xor_out[21][19][8] + xor_out[22][19][8] + xor_out[23][19][8] + xor_out[24][19][8];
assign sum_out[5][19][8] = xor_out[25][19][8] + xor_out[26][19][8] + xor_out[27][19][8] + xor_out[28][19][8] + xor_out[29][19][8];
assign sum_out[6][19][8] = xor_out[30][19][8] + xor_out[31][19][8] + xor_out[32][19][8] + xor_out[33][19][8] + xor_out[34][19][8];
assign sum_out[7][19][8] = xor_out[35][19][8] + xor_out[36][19][8] + xor_out[37][19][8] + xor_out[38][19][8] + xor_out[39][19][8];
assign sum_out[8][19][8] = xor_out[40][19][8] + xor_out[41][19][8] + xor_out[42][19][8] + xor_out[43][19][8] + xor_out[44][19][8];
assign sum_out[9][19][8] = xor_out[45][19][8] + xor_out[46][19][8] + xor_out[47][19][8] + xor_out[48][19][8] + xor_out[49][19][8];
assign sum_out[10][19][8] = xor_out[50][19][8] + xor_out[51][19][8] + xor_out[52][19][8] + xor_out[53][19][8] + xor_out[54][19][8];
assign sum_out[11][19][8] = xor_out[55][19][8] + xor_out[56][19][8] + xor_out[57][19][8] + xor_out[58][19][8] + xor_out[59][19][8];
assign sum_out[12][19][8] = xor_out[60][19][8] + xor_out[61][19][8] + xor_out[62][19][8] + xor_out[63][19][8] + xor_out[64][19][8];
assign sum_out[13][19][8] = xor_out[65][19][8] + xor_out[66][19][8] + xor_out[67][19][8] + xor_out[68][19][8] + xor_out[69][19][8];
assign sum_out[14][19][8] = xor_out[70][19][8] + xor_out[71][19][8] + xor_out[72][19][8] + xor_out[73][19][8] + xor_out[74][19][8];
assign sum_out[15][19][8] = xor_out[75][19][8] + xor_out[76][19][8] + xor_out[77][19][8] + xor_out[78][19][8] + xor_out[79][19][8];
assign sum_out[16][19][8] = xor_out[80][19][8] + xor_out[81][19][8] + xor_out[82][19][8] + xor_out[83][19][8] + xor_out[84][19][8];
assign sum_out[17][19][8] = xor_out[85][19][8] + xor_out[86][19][8] + xor_out[87][19][8] + xor_out[88][19][8] + xor_out[89][19][8];
assign sum_out[18][19][8] = xor_out[90][19][8] + xor_out[91][19][8] + xor_out[92][19][8] + xor_out[93][19][8] + xor_out[94][19][8];
assign sum_out[19][19][8] = xor_out[95][19][8] + xor_out[96][19][8] + xor_out[97][19][8] + xor_out[98][19][8] + xor_out[99][19][8];

assign sum_out[0][19][9] = xor_out[0][19][9] + xor_out[1][19][9] + xor_out[2][19][9] + xor_out[3][19][9] + xor_out[4][19][9];
assign sum_out[1][19][9] = xor_out[5][19][9] + xor_out[6][19][9] + xor_out[7][19][9] + xor_out[8][19][9] + xor_out[9][19][9];
assign sum_out[2][19][9] = xor_out[10][19][9] + xor_out[11][19][9] + xor_out[12][19][9] + xor_out[13][19][9] + xor_out[14][19][9];
assign sum_out[3][19][9] = xor_out[15][19][9] + xor_out[16][19][9] + xor_out[17][19][9] + xor_out[18][19][9] + xor_out[19][19][9];
assign sum_out[4][19][9] = xor_out[20][19][9] + xor_out[21][19][9] + xor_out[22][19][9] + xor_out[23][19][9] + xor_out[24][19][9];
assign sum_out[5][19][9] = xor_out[25][19][9] + xor_out[26][19][9] + xor_out[27][19][9] + xor_out[28][19][9] + xor_out[29][19][9];
assign sum_out[6][19][9] = xor_out[30][19][9] + xor_out[31][19][9] + xor_out[32][19][9] + xor_out[33][19][9] + xor_out[34][19][9];
assign sum_out[7][19][9] = xor_out[35][19][9] + xor_out[36][19][9] + xor_out[37][19][9] + xor_out[38][19][9] + xor_out[39][19][9];
assign sum_out[8][19][9] = xor_out[40][19][9] + xor_out[41][19][9] + xor_out[42][19][9] + xor_out[43][19][9] + xor_out[44][19][9];
assign sum_out[9][19][9] = xor_out[45][19][9] + xor_out[46][19][9] + xor_out[47][19][9] + xor_out[48][19][9] + xor_out[49][19][9];
assign sum_out[10][19][9] = xor_out[50][19][9] + xor_out[51][19][9] + xor_out[52][19][9] + xor_out[53][19][9] + xor_out[54][19][9];
assign sum_out[11][19][9] = xor_out[55][19][9] + xor_out[56][19][9] + xor_out[57][19][9] + xor_out[58][19][9] + xor_out[59][19][9];
assign sum_out[12][19][9] = xor_out[60][19][9] + xor_out[61][19][9] + xor_out[62][19][9] + xor_out[63][19][9] + xor_out[64][19][9];
assign sum_out[13][19][9] = xor_out[65][19][9] + xor_out[66][19][9] + xor_out[67][19][9] + xor_out[68][19][9] + xor_out[69][19][9];
assign sum_out[14][19][9] = xor_out[70][19][9] + xor_out[71][19][9] + xor_out[72][19][9] + xor_out[73][19][9] + xor_out[74][19][9];
assign sum_out[15][19][9] = xor_out[75][19][9] + xor_out[76][19][9] + xor_out[77][19][9] + xor_out[78][19][9] + xor_out[79][19][9];
assign sum_out[16][19][9] = xor_out[80][19][9] + xor_out[81][19][9] + xor_out[82][19][9] + xor_out[83][19][9] + xor_out[84][19][9];
assign sum_out[17][19][9] = xor_out[85][19][9] + xor_out[86][19][9] + xor_out[87][19][9] + xor_out[88][19][9] + xor_out[89][19][9];
assign sum_out[18][19][9] = xor_out[90][19][9] + xor_out[91][19][9] + xor_out[92][19][9] + xor_out[93][19][9] + xor_out[94][19][9];
assign sum_out[19][19][9] = xor_out[95][19][9] + xor_out[96][19][9] + xor_out[97][19][9] + xor_out[98][19][9] + xor_out[99][19][9];

assign sum_out[0][19][10] = xor_out[0][19][10] + xor_out[1][19][10] + xor_out[2][19][10] + xor_out[3][19][10] + xor_out[4][19][10];
assign sum_out[1][19][10] = xor_out[5][19][10] + xor_out[6][19][10] + xor_out[7][19][10] + xor_out[8][19][10] + xor_out[9][19][10];
assign sum_out[2][19][10] = xor_out[10][19][10] + xor_out[11][19][10] + xor_out[12][19][10] + xor_out[13][19][10] + xor_out[14][19][10];
assign sum_out[3][19][10] = xor_out[15][19][10] + xor_out[16][19][10] + xor_out[17][19][10] + xor_out[18][19][10] + xor_out[19][19][10];
assign sum_out[4][19][10] = xor_out[20][19][10] + xor_out[21][19][10] + xor_out[22][19][10] + xor_out[23][19][10] + xor_out[24][19][10];
assign sum_out[5][19][10] = xor_out[25][19][10] + xor_out[26][19][10] + xor_out[27][19][10] + xor_out[28][19][10] + xor_out[29][19][10];
assign sum_out[6][19][10] = xor_out[30][19][10] + xor_out[31][19][10] + xor_out[32][19][10] + xor_out[33][19][10] + xor_out[34][19][10];
assign sum_out[7][19][10] = xor_out[35][19][10] + xor_out[36][19][10] + xor_out[37][19][10] + xor_out[38][19][10] + xor_out[39][19][10];
assign sum_out[8][19][10] = xor_out[40][19][10] + xor_out[41][19][10] + xor_out[42][19][10] + xor_out[43][19][10] + xor_out[44][19][10];
assign sum_out[9][19][10] = xor_out[45][19][10] + xor_out[46][19][10] + xor_out[47][19][10] + xor_out[48][19][10] + xor_out[49][19][10];
assign sum_out[10][19][10] = xor_out[50][19][10] + xor_out[51][19][10] + xor_out[52][19][10] + xor_out[53][19][10] + xor_out[54][19][10];
assign sum_out[11][19][10] = xor_out[55][19][10] + xor_out[56][19][10] + xor_out[57][19][10] + xor_out[58][19][10] + xor_out[59][19][10];
assign sum_out[12][19][10] = xor_out[60][19][10] + xor_out[61][19][10] + xor_out[62][19][10] + xor_out[63][19][10] + xor_out[64][19][10];
assign sum_out[13][19][10] = xor_out[65][19][10] + xor_out[66][19][10] + xor_out[67][19][10] + xor_out[68][19][10] + xor_out[69][19][10];
assign sum_out[14][19][10] = xor_out[70][19][10] + xor_out[71][19][10] + xor_out[72][19][10] + xor_out[73][19][10] + xor_out[74][19][10];
assign sum_out[15][19][10] = xor_out[75][19][10] + xor_out[76][19][10] + xor_out[77][19][10] + xor_out[78][19][10] + xor_out[79][19][10];
assign sum_out[16][19][10] = xor_out[80][19][10] + xor_out[81][19][10] + xor_out[82][19][10] + xor_out[83][19][10] + xor_out[84][19][10];
assign sum_out[17][19][10] = xor_out[85][19][10] + xor_out[86][19][10] + xor_out[87][19][10] + xor_out[88][19][10] + xor_out[89][19][10];
assign sum_out[18][19][10] = xor_out[90][19][10] + xor_out[91][19][10] + xor_out[92][19][10] + xor_out[93][19][10] + xor_out[94][19][10];
assign sum_out[19][19][10] = xor_out[95][19][10] + xor_out[96][19][10] + xor_out[97][19][10] + xor_out[98][19][10] + xor_out[99][19][10];

assign sum_out[0][19][11] = xor_out[0][19][11] + xor_out[1][19][11] + xor_out[2][19][11] + xor_out[3][19][11] + xor_out[4][19][11];
assign sum_out[1][19][11] = xor_out[5][19][11] + xor_out[6][19][11] + xor_out[7][19][11] + xor_out[8][19][11] + xor_out[9][19][11];
assign sum_out[2][19][11] = xor_out[10][19][11] + xor_out[11][19][11] + xor_out[12][19][11] + xor_out[13][19][11] + xor_out[14][19][11];
assign sum_out[3][19][11] = xor_out[15][19][11] + xor_out[16][19][11] + xor_out[17][19][11] + xor_out[18][19][11] + xor_out[19][19][11];
assign sum_out[4][19][11] = xor_out[20][19][11] + xor_out[21][19][11] + xor_out[22][19][11] + xor_out[23][19][11] + xor_out[24][19][11];
assign sum_out[5][19][11] = xor_out[25][19][11] + xor_out[26][19][11] + xor_out[27][19][11] + xor_out[28][19][11] + xor_out[29][19][11];
assign sum_out[6][19][11] = xor_out[30][19][11] + xor_out[31][19][11] + xor_out[32][19][11] + xor_out[33][19][11] + xor_out[34][19][11];
assign sum_out[7][19][11] = xor_out[35][19][11] + xor_out[36][19][11] + xor_out[37][19][11] + xor_out[38][19][11] + xor_out[39][19][11];
assign sum_out[8][19][11] = xor_out[40][19][11] + xor_out[41][19][11] + xor_out[42][19][11] + xor_out[43][19][11] + xor_out[44][19][11];
assign sum_out[9][19][11] = xor_out[45][19][11] + xor_out[46][19][11] + xor_out[47][19][11] + xor_out[48][19][11] + xor_out[49][19][11];
assign sum_out[10][19][11] = xor_out[50][19][11] + xor_out[51][19][11] + xor_out[52][19][11] + xor_out[53][19][11] + xor_out[54][19][11];
assign sum_out[11][19][11] = xor_out[55][19][11] + xor_out[56][19][11] + xor_out[57][19][11] + xor_out[58][19][11] + xor_out[59][19][11];
assign sum_out[12][19][11] = xor_out[60][19][11] + xor_out[61][19][11] + xor_out[62][19][11] + xor_out[63][19][11] + xor_out[64][19][11];
assign sum_out[13][19][11] = xor_out[65][19][11] + xor_out[66][19][11] + xor_out[67][19][11] + xor_out[68][19][11] + xor_out[69][19][11];
assign sum_out[14][19][11] = xor_out[70][19][11] + xor_out[71][19][11] + xor_out[72][19][11] + xor_out[73][19][11] + xor_out[74][19][11];
assign sum_out[15][19][11] = xor_out[75][19][11] + xor_out[76][19][11] + xor_out[77][19][11] + xor_out[78][19][11] + xor_out[79][19][11];
assign sum_out[16][19][11] = xor_out[80][19][11] + xor_out[81][19][11] + xor_out[82][19][11] + xor_out[83][19][11] + xor_out[84][19][11];
assign sum_out[17][19][11] = xor_out[85][19][11] + xor_out[86][19][11] + xor_out[87][19][11] + xor_out[88][19][11] + xor_out[89][19][11];
assign sum_out[18][19][11] = xor_out[90][19][11] + xor_out[91][19][11] + xor_out[92][19][11] + xor_out[93][19][11] + xor_out[94][19][11];
assign sum_out[19][19][11] = xor_out[95][19][11] + xor_out[96][19][11] + xor_out[97][19][11] + xor_out[98][19][11] + xor_out[99][19][11];

assign sum_out[0][19][12] = xor_out[0][19][12] + xor_out[1][19][12] + xor_out[2][19][12] + xor_out[3][19][12] + xor_out[4][19][12];
assign sum_out[1][19][12] = xor_out[5][19][12] + xor_out[6][19][12] + xor_out[7][19][12] + xor_out[8][19][12] + xor_out[9][19][12];
assign sum_out[2][19][12] = xor_out[10][19][12] + xor_out[11][19][12] + xor_out[12][19][12] + xor_out[13][19][12] + xor_out[14][19][12];
assign sum_out[3][19][12] = xor_out[15][19][12] + xor_out[16][19][12] + xor_out[17][19][12] + xor_out[18][19][12] + xor_out[19][19][12];
assign sum_out[4][19][12] = xor_out[20][19][12] + xor_out[21][19][12] + xor_out[22][19][12] + xor_out[23][19][12] + xor_out[24][19][12];
assign sum_out[5][19][12] = xor_out[25][19][12] + xor_out[26][19][12] + xor_out[27][19][12] + xor_out[28][19][12] + xor_out[29][19][12];
assign sum_out[6][19][12] = xor_out[30][19][12] + xor_out[31][19][12] + xor_out[32][19][12] + xor_out[33][19][12] + xor_out[34][19][12];
assign sum_out[7][19][12] = xor_out[35][19][12] + xor_out[36][19][12] + xor_out[37][19][12] + xor_out[38][19][12] + xor_out[39][19][12];
assign sum_out[8][19][12] = xor_out[40][19][12] + xor_out[41][19][12] + xor_out[42][19][12] + xor_out[43][19][12] + xor_out[44][19][12];
assign sum_out[9][19][12] = xor_out[45][19][12] + xor_out[46][19][12] + xor_out[47][19][12] + xor_out[48][19][12] + xor_out[49][19][12];
assign sum_out[10][19][12] = xor_out[50][19][12] + xor_out[51][19][12] + xor_out[52][19][12] + xor_out[53][19][12] + xor_out[54][19][12];
assign sum_out[11][19][12] = xor_out[55][19][12] + xor_out[56][19][12] + xor_out[57][19][12] + xor_out[58][19][12] + xor_out[59][19][12];
assign sum_out[12][19][12] = xor_out[60][19][12] + xor_out[61][19][12] + xor_out[62][19][12] + xor_out[63][19][12] + xor_out[64][19][12];
assign sum_out[13][19][12] = xor_out[65][19][12] + xor_out[66][19][12] + xor_out[67][19][12] + xor_out[68][19][12] + xor_out[69][19][12];
assign sum_out[14][19][12] = xor_out[70][19][12] + xor_out[71][19][12] + xor_out[72][19][12] + xor_out[73][19][12] + xor_out[74][19][12];
assign sum_out[15][19][12] = xor_out[75][19][12] + xor_out[76][19][12] + xor_out[77][19][12] + xor_out[78][19][12] + xor_out[79][19][12];
assign sum_out[16][19][12] = xor_out[80][19][12] + xor_out[81][19][12] + xor_out[82][19][12] + xor_out[83][19][12] + xor_out[84][19][12];
assign sum_out[17][19][12] = xor_out[85][19][12] + xor_out[86][19][12] + xor_out[87][19][12] + xor_out[88][19][12] + xor_out[89][19][12];
assign sum_out[18][19][12] = xor_out[90][19][12] + xor_out[91][19][12] + xor_out[92][19][12] + xor_out[93][19][12] + xor_out[94][19][12];
assign sum_out[19][19][12] = xor_out[95][19][12] + xor_out[96][19][12] + xor_out[97][19][12] + xor_out[98][19][12] + xor_out[99][19][12];

assign sum_out[0][19][13] = xor_out[0][19][13] + xor_out[1][19][13] + xor_out[2][19][13] + xor_out[3][19][13] + xor_out[4][19][13];
assign sum_out[1][19][13] = xor_out[5][19][13] + xor_out[6][19][13] + xor_out[7][19][13] + xor_out[8][19][13] + xor_out[9][19][13];
assign sum_out[2][19][13] = xor_out[10][19][13] + xor_out[11][19][13] + xor_out[12][19][13] + xor_out[13][19][13] + xor_out[14][19][13];
assign sum_out[3][19][13] = xor_out[15][19][13] + xor_out[16][19][13] + xor_out[17][19][13] + xor_out[18][19][13] + xor_out[19][19][13];
assign sum_out[4][19][13] = xor_out[20][19][13] + xor_out[21][19][13] + xor_out[22][19][13] + xor_out[23][19][13] + xor_out[24][19][13];
assign sum_out[5][19][13] = xor_out[25][19][13] + xor_out[26][19][13] + xor_out[27][19][13] + xor_out[28][19][13] + xor_out[29][19][13];
assign sum_out[6][19][13] = xor_out[30][19][13] + xor_out[31][19][13] + xor_out[32][19][13] + xor_out[33][19][13] + xor_out[34][19][13];
assign sum_out[7][19][13] = xor_out[35][19][13] + xor_out[36][19][13] + xor_out[37][19][13] + xor_out[38][19][13] + xor_out[39][19][13];
assign sum_out[8][19][13] = xor_out[40][19][13] + xor_out[41][19][13] + xor_out[42][19][13] + xor_out[43][19][13] + xor_out[44][19][13];
assign sum_out[9][19][13] = xor_out[45][19][13] + xor_out[46][19][13] + xor_out[47][19][13] + xor_out[48][19][13] + xor_out[49][19][13];
assign sum_out[10][19][13] = xor_out[50][19][13] + xor_out[51][19][13] + xor_out[52][19][13] + xor_out[53][19][13] + xor_out[54][19][13];
assign sum_out[11][19][13] = xor_out[55][19][13] + xor_out[56][19][13] + xor_out[57][19][13] + xor_out[58][19][13] + xor_out[59][19][13];
assign sum_out[12][19][13] = xor_out[60][19][13] + xor_out[61][19][13] + xor_out[62][19][13] + xor_out[63][19][13] + xor_out[64][19][13];
assign sum_out[13][19][13] = xor_out[65][19][13] + xor_out[66][19][13] + xor_out[67][19][13] + xor_out[68][19][13] + xor_out[69][19][13];
assign sum_out[14][19][13] = xor_out[70][19][13] + xor_out[71][19][13] + xor_out[72][19][13] + xor_out[73][19][13] + xor_out[74][19][13];
assign sum_out[15][19][13] = xor_out[75][19][13] + xor_out[76][19][13] + xor_out[77][19][13] + xor_out[78][19][13] + xor_out[79][19][13];
assign sum_out[16][19][13] = xor_out[80][19][13] + xor_out[81][19][13] + xor_out[82][19][13] + xor_out[83][19][13] + xor_out[84][19][13];
assign sum_out[17][19][13] = xor_out[85][19][13] + xor_out[86][19][13] + xor_out[87][19][13] + xor_out[88][19][13] + xor_out[89][19][13];
assign sum_out[18][19][13] = xor_out[90][19][13] + xor_out[91][19][13] + xor_out[92][19][13] + xor_out[93][19][13] + xor_out[94][19][13];
assign sum_out[19][19][13] = xor_out[95][19][13] + xor_out[96][19][13] + xor_out[97][19][13] + xor_out[98][19][13] + xor_out[99][19][13];

assign sum_out[0][19][14] = xor_out[0][19][14] + xor_out[1][19][14] + xor_out[2][19][14] + xor_out[3][19][14] + xor_out[4][19][14];
assign sum_out[1][19][14] = xor_out[5][19][14] + xor_out[6][19][14] + xor_out[7][19][14] + xor_out[8][19][14] + xor_out[9][19][14];
assign sum_out[2][19][14] = xor_out[10][19][14] + xor_out[11][19][14] + xor_out[12][19][14] + xor_out[13][19][14] + xor_out[14][19][14];
assign sum_out[3][19][14] = xor_out[15][19][14] + xor_out[16][19][14] + xor_out[17][19][14] + xor_out[18][19][14] + xor_out[19][19][14];
assign sum_out[4][19][14] = xor_out[20][19][14] + xor_out[21][19][14] + xor_out[22][19][14] + xor_out[23][19][14] + xor_out[24][19][14];
assign sum_out[5][19][14] = xor_out[25][19][14] + xor_out[26][19][14] + xor_out[27][19][14] + xor_out[28][19][14] + xor_out[29][19][14];
assign sum_out[6][19][14] = xor_out[30][19][14] + xor_out[31][19][14] + xor_out[32][19][14] + xor_out[33][19][14] + xor_out[34][19][14];
assign sum_out[7][19][14] = xor_out[35][19][14] + xor_out[36][19][14] + xor_out[37][19][14] + xor_out[38][19][14] + xor_out[39][19][14];
assign sum_out[8][19][14] = xor_out[40][19][14] + xor_out[41][19][14] + xor_out[42][19][14] + xor_out[43][19][14] + xor_out[44][19][14];
assign sum_out[9][19][14] = xor_out[45][19][14] + xor_out[46][19][14] + xor_out[47][19][14] + xor_out[48][19][14] + xor_out[49][19][14];
assign sum_out[10][19][14] = xor_out[50][19][14] + xor_out[51][19][14] + xor_out[52][19][14] + xor_out[53][19][14] + xor_out[54][19][14];
assign sum_out[11][19][14] = xor_out[55][19][14] + xor_out[56][19][14] + xor_out[57][19][14] + xor_out[58][19][14] + xor_out[59][19][14];
assign sum_out[12][19][14] = xor_out[60][19][14] + xor_out[61][19][14] + xor_out[62][19][14] + xor_out[63][19][14] + xor_out[64][19][14];
assign sum_out[13][19][14] = xor_out[65][19][14] + xor_out[66][19][14] + xor_out[67][19][14] + xor_out[68][19][14] + xor_out[69][19][14];
assign sum_out[14][19][14] = xor_out[70][19][14] + xor_out[71][19][14] + xor_out[72][19][14] + xor_out[73][19][14] + xor_out[74][19][14];
assign sum_out[15][19][14] = xor_out[75][19][14] + xor_out[76][19][14] + xor_out[77][19][14] + xor_out[78][19][14] + xor_out[79][19][14];
assign sum_out[16][19][14] = xor_out[80][19][14] + xor_out[81][19][14] + xor_out[82][19][14] + xor_out[83][19][14] + xor_out[84][19][14];
assign sum_out[17][19][14] = xor_out[85][19][14] + xor_out[86][19][14] + xor_out[87][19][14] + xor_out[88][19][14] + xor_out[89][19][14];
assign sum_out[18][19][14] = xor_out[90][19][14] + xor_out[91][19][14] + xor_out[92][19][14] + xor_out[93][19][14] + xor_out[94][19][14];
assign sum_out[19][19][14] = xor_out[95][19][14] + xor_out[96][19][14] + xor_out[97][19][14] + xor_out[98][19][14] + xor_out[99][19][14];

assign sum_out[0][19][15] = xor_out[0][19][15] + xor_out[1][19][15] + xor_out[2][19][15] + xor_out[3][19][15] + xor_out[4][19][15];
assign sum_out[1][19][15] = xor_out[5][19][15] + xor_out[6][19][15] + xor_out[7][19][15] + xor_out[8][19][15] + xor_out[9][19][15];
assign sum_out[2][19][15] = xor_out[10][19][15] + xor_out[11][19][15] + xor_out[12][19][15] + xor_out[13][19][15] + xor_out[14][19][15];
assign sum_out[3][19][15] = xor_out[15][19][15] + xor_out[16][19][15] + xor_out[17][19][15] + xor_out[18][19][15] + xor_out[19][19][15];
assign sum_out[4][19][15] = xor_out[20][19][15] + xor_out[21][19][15] + xor_out[22][19][15] + xor_out[23][19][15] + xor_out[24][19][15];
assign sum_out[5][19][15] = xor_out[25][19][15] + xor_out[26][19][15] + xor_out[27][19][15] + xor_out[28][19][15] + xor_out[29][19][15];
assign sum_out[6][19][15] = xor_out[30][19][15] + xor_out[31][19][15] + xor_out[32][19][15] + xor_out[33][19][15] + xor_out[34][19][15];
assign sum_out[7][19][15] = xor_out[35][19][15] + xor_out[36][19][15] + xor_out[37][19][15] + xor_out[38][19][15] + xor_out[39][19][15];
assign sum_out[8][19][15] = xor_out[40][19][15] + xor_out[41][19][15] + xor_out[42][19][15] + xor_out[43][19][15] + xor_out[44][19][15];
assign sum_out[9][19][15] = xor_out[45][19][15] + xor_out[46][19][15] + xor_out[47][19][15] + xor_out[48][19][15] + xor_out[49][19][15];
assign sum_out[10][19][15] = xor_out[50][19][15] + xor_out[51][19][15] + xor_out[52][19][15] + xor_out[53][19][15] + xor_out[54][19][15];
assign sum_out[11][19][15] = xor_out[55][19][15] + xor_out[56][19][15] + xor_out[57][19][15] + xor_out[58][19][15] + xor_out[59][19][15];
assign sum_out[12][19][15] = xor_out[60][19][15] + xor_out[61][19][15] + xor_out[62][19][15] + xor_out[63][19][15] + xor_out[64][19][15];
assign sum_out[13][19][15] = xor_out[65][19][15] + xor_out[66][19][15] + xor_out[67][19][15] + xor_out[68][19][15] + xor_out[69][19][15];
assign sum_out[14][19][15] = xor_out[70][19][15] + xor_out[71][19][15] + xor_out[72][19][15] + xor_out[73][19][15] + xor_out[74][19][15];
assign sum_out[15][19][15] = xor_out[75][19][15] + xor_out[76][19][15] + xor_out[77][19][15] + xor_out[78][19][15] + xor_out[79][19][15];
assign sum_out[16][19][15] = xor_out[80][19][15] + xor_out[81][19][15] + xor_out[82][19][15] + xor_out[83][19][15] + xor_out[84][19][15];
assign sum_out[17][19][15] = xor_out[85][19][15] + xor_out[86][19][15] + xor_out[87][19][15] + xor_out[88][19][15] + xor_out[89][19][15];
assign sum_out[18][19][15] = xor_out[90][19][15] + xor_out[91][19][15] + xor_out[92][19][15] + xor_out[93][19][15] + xor_out[94][19][15];
assign sum_out[19][19][15] = xor_out[95][19][15] + xor_out[96][19][15] + xor_out[97][19][15] + xor_out[98][19][15] + xor_out[99][19][15];

assign sum_out[0][19][16] = xor_out[0][19][16] + xor_out[1][19][16] + xor_out[2][19][16] + xor_out[3][19][16] + xor_out[4][19][16];
assign sum_out[1][19][16] = xor_out[5][19][16] + xor_out[6][19][16] + xor_out[7][19][16] + xor_out[8][19][16] + xor_out[9][19][16];
assign sum_out[2][19][16] = xor_out[10][19][16] + xor_out[11][19][16] + xor_out[12][19][16] + xor_out[13][19][16] + xor_out[14][19][16];
assign sum_out[3][19][16] = xor_out[15][19][16] + xor_out[16][19][16] + xor_out[17][19][16] + xor_out[18][19][16] + xor_out[19][19][16];
assign sum_out[4][19][16] = xor_out[20][19][16] + xor_out[21][19][16] + xor_out[22][19][16] + xor_out[23][19][16] + xor_out[24][19][16];
assign sum_out[5][19][16] = xor_out[25][19][16] + xor_out[26][19][16] + xor_out[27][19][16] + xor_out[28][19][16] + xor_out[29][19][16];
assign sum_out[6][19][16] = xor_out[30][19][16] + xor_out[31][19][16] + xor_out[32][19][16] + xor_out[33][19][16] + xor_out[34][19][16];
assign sum_out[7][19][16] = xor_out[35][19][16] + xor_out[36][19][16] + xor_out[37][19][16] + xor_out[38][19][16] + xor_out[39][19][16];
assign sum_out[8][19][16] = xor_out[40][19][16] + xor_out[41][19][16] + xor_out[42][19][16] + xor_out[43][19][16] + xor_out[44][19][16];
assign sum_out[9][19][16] = xor_out[45][19][16] + xor_out[46][19][16] + xor_out[47][19][16] + xor_out[48][19][16] + xor_out[49][19][16];
assign sum_out[10][19][16] = xor_out[50][19][16] + xor_out[51][19][16] + xor_out[52][19][16] + xor_out[53][19][16] + xor_out[54][19][16];
assign sum_out[11][19][16] = xor_out[55][19][16] + xor_out[56][19][16] + xor_out[57][19][16] + xor_out[58][19][16] + xor_out[59][19][16];
assign sum_out[12][19][16] = xor_out[60][19][16] + xor_out[61][19][16] + xor_out[62][19][16] + xor_out[63][19][16] + xor_out[64][19][16];
assign sum_out[13][19][16] = xor_out[65][19][16] + xor_out[66][19][16] + xor_out[67][19][16] + xor_out[68][19][16] + xor_out[69][19][16];
assign sum_out[14][19][16] = xor_out[70][19][16] + xor_out[71][19][16] + xor_out[72][19][16] + xor_out[73][19][16] + xor_out[74][19][16];
assign sum_out[15][19][16] = xor_out[75][19][16] + xor_out[76][19][16] + xor_out[77][19][16] + xor_out[78][19][16] + xor_out[79][19][16];
assign sum_out[16][19][16] = xor_out[80][19][16] + xor_out[81][19][16] + xor_out[82][19][16] + xor_out[83][19][16] + xor_out[84][19][16];
assign sum_out[17][19][16] = xor_out[85][19][16] + xor_out[86][19][16] + xor_out[87][19][16] + xor_out[88][19][16] + xor_out[89][19][16];
assign sum_out[18][19][16] = xor_out[90][19][16] + xor_out[91][19][16] + xor_out[92][19][16] + xor_out[93][19][16] + xor_out[94][19][16];
assign sum_out[19][19][16] = xor_out[95][19][16] + xor_out[96][19][16] + xor_out[97][19][16] + xor_out[98][19][16] + xor_out[99][19][16];

assign sum_out[0][19][17] = xor_out[0][19][17] + xor_out[1][19][17] + xor_out[2][19][17] + xor_out[3][19][17] + xor_out[4][19][17];
assign sum_out[1][19][17] = xor_out[5][19][17] + xor_out[6][19][17] + xor_out[7][19][17] + xor_out[8][19][17] + xor_out[9][19][17];
assign sum_out[2][19][17] = xor_out[10][19][17] + xor_out[11][19][17] + xor_out[12][19][17] + xor_out[13][19][17] + xor_out[14][19][17];
assign sum_out[3][19][17] = xor_out[15][19][17] + xor_out[16][19][17] + xor_out[17][19][17] + xor_out[18][19][17] + xor_out[19][19][17];
assign sum_out[4][19][17] = xor_out[20][19][17] + xor_out[21][19][17] + xor_out[22][19][17] + xor_out[23][19][17] + xor_out[24][19][17];
assign sum_out[5][19][17] = xor_out[25][19][17] + xor_out[26][19][17] + xor_out[27][19][17] + xor_out[28][19][17] + xor_out[29][19][17];
assign sum_out[6][19][17] = xor_out[30][19][17] + xor_out[31][19][17] + xor_out[32][19][17] + xor_out[33][19][17] + xor_out[34][19][17];
assign sum_out[7][19][17] = xor_out[35][19][17] + xor_out[36][19][17] + xor_out[37][19][17] + xor_out[38][19][17] + xor_out[39][19][17];
assign sum_out[8][19][17] = xor_out[40][19][17] + xor_out[41][19][17] + xor_out[42][19][17] + xor_out[43][19][17] + xor_out[44][19][17];
assign sum_out[9][19][17] = xor_out[45][19][17] + xor_out[46][19][17] + xor_out[47][19][17] + xor_out[48][19][17] + xor_out[49][19][17];
assign sum_out[10][19][17] = xor_out[50][19][17] + xor_out[51][19][17] + xor_out[52][19][17] + xor_out[53][19][17] + xor_out[54][19][17];
assign sum_out[11][19][17] = xor_out[55][19][17] + xor_out[56][19][17] + xor_out[57][19][17] + xor_out[58][19][17] + xor_out[59][19][17];
assign sum_out[12][19][17] = xor_out[60][19][17] + xor_out[61][19][17] + xor_out[62][19][17] + xor_out[63][19][17] + xor_out[64][19][17];
assign sum_out[13][19][17] = xor_out[65][19][17] + xor_out[66][19][17] + xor_out[67][19][17] + xor_out[68][19][17] + xor_out[69][19][17];
assign sum_out[14][19][17] = xor_out[70][19][17] + xor_out[71][19][17] + xor_out[72][19][17] + xor_out[73][19][17] + xor_out[74][19][17];
assign sum_out[15][19][17] = xor_out[75][19][17] + xor_out[76][19][17] + xor_out[77][19][17] + xor_out[78][19][17] + xor_out[79][19][17];
assign sum_out[16][19][17] = xor_out[80][19][17] + xor_out[81][19][17] + xor_out[82][19][17] + xor_out[83][19][17] + xor_out[84][19][17];
assign sum_out[17][19][17] = xor_out[85][19][17] + xor_out[86][19][17] + xor_out[87][19][17] + xor_out[88][19][17] + xor_out[89][19][17];
assign sum_out[18][19][17] = xor_out[90][19][17] + xor_out[91][19][17] + xor_out[92][19][17] + xor_out[93][19][17] + xor_out[94][19][17];
assign sum_out[19][19][17] = xor_out[95][19][17] + xor_out[96][19][17] + xor_out[97][19][17] + xor_out[98][19][17] + xor_out[99][19][17];

assign sum_out[0][19][18] = xor_out[0][19][18] + xor_out[1][19][18] + xor_out[2][19][18] + xor_out[3][19][18] + xor_out[4][19][18];
assign sum_out[1][19][18] = xor_out[5][19][18] + xor_out[6][19][18] + xor_out[7][19][18] + xor_out[8][19][18] + xor_out[9][19][18];
assign sum_out[2][19][18] = xor_out[10][19][18] + xor_out[11][19][18] + xor_out[12][19][18] + xor_out[13][19][18] + xor_out[14][19][18];
assign sum_out[3][19][18] = xor_out[15][19][18] + xor_out[16][19][18] + xor_out[17][19][18] + xor_out[18][19][18] + xor_out[19][19][18];
assign sum_out[4][19][18] = xor_out[20][19][18] + xor_out[21][19][18] + xor_out[22][19][18] + xor_out[23][19][18] + xor_out[24][19][18];
assign sum_out[5][19][18] = xor_out[25][19][18] + xor_out[26][19][18] + xor_out[27][19][18] + xor_out[28][19][18] + xor_out[29][19][18];
assign sum_out[6][19][18] = xor_out[30][19][18] + xor_out[31][19][18] + xor_out[32][19][18] + xor_out[33][19][18] + xor_out[34][19][18];
assign sum_out[7][19][18] = xor_out[35][19][18] + xor_out[36][19][18] + xor_out[37][19][18] + xor_out[38][19][18] + xor_out[39][19][18];
assign sum_out[8][19][18] = xor_out[40][19][18] + xor_out[41][19][18] + xor_out[42][19][18] + xor_out[43][19][18] + xor_out[44][19][18];
assign sum_out[9][19][18] = xor_out[45][19][18] + xor_out[46][19][18] + xor_out[47][19][18] + xor_out[48][19][18] + xor_out[49][19][18];
assign sum_out[10][19][18] = xor_out[50][19][18] + xor_out[51][19][18] + xor_out[52][19][18] + xor_out[53][19][18] + xor_out[54][19][18];
assign sum_out[11][19][18] = xor_out[55][19][18] + xor_out[56][19][18] + xor_out[57][19][18] + xor_out[58][19][18] + xor_out[59][19][18];
assign sum_out[12][19][18] = xor_out[60][19][18] + xor_out[61][19][18] + xor_out[62][19][18] + xor_out[63][19][18] + xor_out[64][19][18];
assign sum_out[13][19][18] = xor_out[65][19][18] + xor_out[66][19][18] + xor_out[67][19][18] + xor_out[68][19][18] + xor_out[69][19][18];
assign sum_out[14][19][18] = xor_out[70][19][18] + xor_out[71][19][18] + xor_out[72][19][18] + xor_out[73][19][18] + xor_out[74][19][18];
assign sum_out[15][19][18] = xor_out[75][19][18] + xor_out[76][19][18] + xor_out[77][19][18] + xor_out[78][19][18] + xor_out[79][19][18];
assign sum_out[16][19][18] = xor_out[80][19][18] + xor_out[81][19][18] + xor_out[82][19][18] + xor_out[83][19][18] + xor_out[84][19][18];
assign sum_out[17][19][18] = xor_out[85][19][18] + xor_out[86][19][18] + xor_out[87][19][18] + xor_out[88][19][18] + xor_out[89][19][18];
assign sum_out[18][19][18] = xor_out[90][19][18] + xor_out[91][19][18] + xor_out[92][19][18] + xor_out[93][19][18] + xor_out[94][19][18];
assign sum_out[19][19][18] = xor_out[95][19][18] + xor_out[96][19][18] + xor_out[97][19][18] + xor_out[98][19][18] + xor_out[99][19][18];

assign sum_out[0][19][19] = xor_out[0][19][19] + xor_out[1][19][19] + xor_out[2][19][19] + xor_out[3][19][19] + xor_out[4][19][19];
assign sum_out[1][19][19] = xor_out[5][19][19] + xor_out[6][19][19] + xor_out[7][19][19] + xor_out[8][19][19] + xor_out[9][19][19];
assign sum_out[2][19][19] = xor_out[10][19][19] + xor_out[11][19][19] + xor_out[12][19][19] + xor_out[13][19][19] + xor_out[14][19][19];
assign sum_out[3][19][19] = xor_out[15][19][19] + xor_out[16][19][19] + xor_out[17][19][19] + xor_out[18][19][19] + xor_out[19][19][19];
assign sum_out[4][19][19] = xor_out[20][19][19] + xor_out[21][19][19] + xor_out[22][19][19] + xor_out[23][19][19] + xor_out[24][19][19];
assign sum_out[5][19][19] = xor_out[25][19][19] + xor_out[26][19][19] + xor_out[27][19][19] + xor_out[28][19][19] + xor_out[29][19][19];
assign sum_out[6][19][19] = xor_out[30][19][19] + xor_out[31][19][19] + xor_out[32][19][19] + xor_out[33][19][19] + xor_out[34][19][19];
assign sum_out[7][19][19] = xor_out[35][19][19] + xor_out[36][19][19] + xor_out[37][19][19] + xor_out[38][19][19] + xor_out[39][19][19];
assign sum_out[8][19][19] = xor_out[40][19][19] + xor_out[41][19][19] + xor_out[42][19][19] + xor_out[43][19][19] + xor_out[44][19][19];
assign sum_out[9][19][19] = xor_out[45][19][19] + xor_out[46][19][19] + xor_out[47][19][19] + xor_out[48][19][19] + xor_out[49][19][19];
assign sum_out[10][19][19] = xor_out[50][19][19] + xor_out[51][19][19] + xor_out[52][19][19] + xor_out[53][19][19] + xor_out[54][19][19];
assign sum_out[11][19][19] = xor_out[55][19][19] + xor_out[56][19][19] + xor_out[57][19][19] + xor_out[58][19][19] + xor_out[59][19][19];
assign sum_out[12][19][19] = xor_out[60][19][19] + xor_out[61][19][19] + xor_out[62][19][19] + xor_out[63][19][19] + xor_out[64][19][19];
assign sum_out[13][19][19] = xor_out[65][19][19] + xor_out[66][19][19] + xor_out[67][19][19] + xor_out[68][19][19] + xor_out[69][19][19];
assign sum_out[14][19][19] = xor_out[70][19][19] + xor_out[71][19][19] + xor_out[72][19][19] + xor_out[73][19][19] + xor_out[74][19][19];
assign sum_out[15][19][19] = xor_out[75][19][19] + xor_out[76][19][19] + xor_out[77][19][19] + xor_out[78][19][19] + xor_out[79][19][19];
assign sum_out[16][19][19] = xor_out[80][19][19] + xor_out[81][19][19] + xor_out[82][19][19] + xor_out[83][19][19] + xor_out[84][19][19];
assign sum_out[17][19][19] = xor_out[85][19][19] + xor_out[86][19][19] + xor_out[87][19][19] + xor_out[88][19][19] + xor_out[89][19][19];
assign sum_out[18][19][19] = xor_out[90][19][19] + xor_out[91][19][19] + xor_out[92][19][19] + xor_out[93][19][19] + xor_out[94][19][19];
assign sum_out[19][19][19] = xor_out[95][19][19] + xor_out[96][19][19] + xor_out[97][19][19] + xor_out[98][19][19] + xor_out[99][19][19];

assign sum_out[0][19][20] = xor_out[0][19][20] + xor_out[1][19][20] + xor_out[2][19][20] + xor_out[3][19][20] + xor_out[4][19][20];
assign sum_out[1][19][20] = xor_out[5][19][20] + xor_out[6][19][20] + xor_out[7][19][20] + xor_out[8][19][20] + xor_out[9][19][20];
assign sum_out[2][19][20] = xor_out[10][19][20] + xor_out[11][19][20] + xor_out[12][19][20] + xor_out[13][19][20] + xor_out[14][19][20];
assign sum_out[3][19][20] = xor_out[15][19][20] + xor_out[16][19][20] + xor_out[17][19][20] + xor_out[18][19][20] + xor_out[19][19][20];
assign sum_out[4][19][20] = xor_out[20][19][20] + xor_out[21][19][20] + xor_out[22][19][20] + xor_out[23][19][20] + xor_out[24][19][20];
assign sum_out[5][19][20] = xor_out[25][19][20] + xor_out[26][19][20] + xor_out[27][19][20] + xor_out[28][19][20] + xor_out[29][19][20];
assign sum_out[6][19][20] = xor_out[30][19][20] + xor_out[31][19][20] + xor_out[32][19][20] + xor_out[33][19][20] + xor_out[34][19][20];
assign sum_out[7][19][20] = xor_out[35][19][20] + xor_out[36][19][20] + xor_out[37][19][20] + xor_out[38][19][20] + xor_out[39][19][20];
assign sum_out[8][19][20] = xor_out[40][19][20] + xor_out[41][19][20] + xor_out[42][19][20] + xor_out[43][19][20] + xor_out[44][19][20];
assign sum_out[9][19][20] = xor_out[45][19][20] + xor_out[46][19][20] + xor_out[47][19][20] + xor_out[48][19][20] + xor_out[49][19][20];
assign sum_out[10][19][20] = xor_out[50][19][20] + xor_out[51][19][20] + xor_out[52][19][20] + xor_out[53][19][20] + xor_out[54][19][20];
assign sum_out[11][19][20] = xor_out[55][19][20] + xor_out[56][19][20] + xor_out[57][19][20] + xor_out[58][19][20] + xor_out[59][19][20];
assign sum_out[12][19][20] = xor_out[60][19][20] + xor_out[61][19][20] + xor_out[62][19][20] + xor_out[63][19][20] + xor_out[64][19][20];
assign sum_out[13][19][20] = xor_out[65][19][20] + xor_out[66][19][20] + xor_out[67][19][20] + xor_out[68][19][20] + xor_out[69][19][20];
assign sum_out[14][19][20] = xor_out[70][19][20] + xor_out[71][19][20] + xor_out[72][19][20] + xor_out[73][19][20] + xor_out[74][19][20];
assign sum_out[15][19][20] = xor_out[75][19][20] + xor_out[76][19][20] + xor_out[77][19][20] + xor_out[78][19][20] + xor_out[79][19][20];
assign sum_out[16][19][20] = xor_out[80][19][20] + xor_out[81][19][20] + xor_out[82][19][20] + xor_out[83][19][20] + xor_out[84][19][20];
assign sum_out[17][19][20] = xor_out[85][19][20] + xor_out[86][19][20] + xor_out[87][19][20] + xor_out[88][19][20] + xor_out[89][19][20];
assign sum_out[18][19][20] = xor_out[90][19][20] + xor_out[91][19][20] + xor_out[92][19][20] + xor_out[93][19][20] + xor_out[94][19][20];
assign sum_out[19][19][20] = xor_out[95][19][20] + xor_out[96][19][20] + xor_out[97][19][20] + xor_out[98][19][20] + xor_out[99][19][20];

assign sum_out[0][19][21] = xor_out[0][19][21] + xor_out[1][19][21] + xor_out[2][19][21] + xor_out[3][19][21] + xor_out[4][19][21];
assign sum_out[1][19][21] = xor_out[5][19][21] + xor_out[6][19][21] + xor_out[7][19][21] + xor_out[8][19][21] + xor_out[9][19][21];
assign sum_out[2][19][21] = xor_out[10][19][21] + xor_out[11][19][21] + xor_out[12][19][21] + xor_out[13][19][21] + xor_out[14][19][21];
assign sum_out[3][19][21] = xor_out[15][19][21] + xor_out[16][19][21] + xor_out[17][19][21] + xor_out[18][19][21] + xor_out[19][19][21];
assign sum_out[4][19][21] = xor_out[20][19][21] + xor_out[21][19][21] + xor_out[22][19][21] + xor_out[23][19][21] + xor_out[24][19][21];
assign sum_out[5][19][21] = xor_out[25][19][21] + xor_out[26][19][21] + xor_out[27][19][21] + xor_out[28][19][21] + xor_out[29][19][21];
assign sum_out[6][19][21] = xor_out[30][19][21] + xor_out[31][19][21] + xor_out[32][19][21] + xor_out[33][19][21] + xor_out[34][19][21];
assign sum_out[7][19][21] = xor_out[35][19][21] + xor_out[36][19][21] + xor_out[37][19][21] + xor_out[38][19][21] + xor_out[39][19][21];
assign sum_out[8][19][21] = xor_out[40][19][21] + xor_out[41][19][21] + xor_out[42][19][21] + xor_out[43][19][21] + xor_out[44][19][21];
assign sum_out[9][19][21] = xor_out[45][19][21] + xor_out[46][19][21] + xor_out[47][19][21] + xor_out[48][19][21] + xor_out[49][19][21];
assign sum_out[10][19][21] = xor_out[50][19][21] + xor_out[51][19][21] + xor_out[52][19][21] + xor_out[53][19][21] + xor_out[54][19][21];
assign sum_out[11][19][21] = xor_out[55][19][21] + xor_out[56][19][21] + xor_out[57][19][21] + xor_out[58][19][21] + xor_out[59][19][21];
assign sum_out[12][19][21] = xor_out[60][19][21] + xor_out[61][19][21] + xor_out[62][19][21] + xor_out[63][19][21] + xor_out[64][19][21];
assign sum_out[13][19][21] = xor_out[65][19][21] + xor_out[66][19][21] + xor_out[67][19][21] + xor_out[68][19][21] + xor_out[69][19][21];
assign sum_out[14][19][21] = xor_out[70][19][21] + xor_out[71][19][21] + xor_out[72][19][21] + xor_out[73][19][21] + xor_out[74][19][21];
assign sum_out[15][19][21] = xor_out[75][19][21] + xor_out[76][19][21] + xor_out[77][19][21] + xor_out[78][19][21] + xor_out[79][19][21];
assign sum_out[16][19][21] = xor_out[80][19][21] + xor_out[81][19][21] + xor_out[82][19][21] + xor_out[83][19][21] + xor_out[84][19][21];
assign sum_out[17][19][21] = xor_out[85][19][21] + xor_out[86][19][21] + xor_out[87][19][21] + xor_out[88][19][21] + xor_out[89][19][21];
assign sum_out[18][19][21] = xor_out[90][19][21] + xor_out[91][19][21] + xor_out[92][19][21] + xor_out[93][19][21] + xor_out[94][19][21];
assign sum_out[19][19][21] = xor_out[95][19][21] + xor_out[96][19][21] + xor_out[97][19][21] + xor_out[98][19][21] + xor_out[99][19][21];

assign sum_out[0][19][22] = xor_out[0][19][22] + xor_out[1][19][22] + xor_out[2][19][22] + xor_out[3][19][22] + xor_out[4][19][22];
assign sum_out[1][19][22] = xor_out[5][19][22] + xor_out[6][19][22] + xor_out[7][19][22] + xor_out[8][19][22] + xor_out[9][19][22];
assign sum_out[2][19][22] = xor_out[10][19][22] + xor_out[11][19][22] + xor_out[12][19][22] + xor_out[13][19][22] + xor_out[14][19][22];
assign sum_out[3][19][22] = xor_out[15][19][22] + xor_out[16][19][22] + xor_out[17][19][22] + xor_out[18][19][22] + xor_out[19][19][22];
assign sum_out[4][19][22] = xor_out[20][19][22] + xor_out[21][19][22] + xor_out[22][19][22] + xor_out[23][19][22] + xor_out[24][19][22];
assign sum_out[5][19][22] = xor_out[25][19][22] + xor_out[26][19][22] + xor_out[27][19][22] + xor_out[28][19][22] + xor_out[29][19][22];
assign sum_out[6][19][22] = xor_out[30][19][22] + xor_out[31][19][22] + xor_out[32][19][22] + xor_out[33][19][22] + xor_out[34][19][22];
assign sum_out[7][19][22] = xor_out[35][19][22] + xor_out[36][19][22] + xor_out[37][19][22] + xor_out[38][19][22] + xor_out[39][19][22];
assign sum_out[8][19][22] = xor_out[40][19][22] + xor_out[41][19][22] + xor_out[42][19][22] + xor_out[43][19][22] + xor_out[44][19][22];
assign sum_out[9][19][22] = xor_out[45][19][22] + xor_out[46][19][22] + xor_out[47][19][22] + xor_out[48][19][22] + xor_out[49][19][22];
assign sum_out[10][19][22] = xor_out[50][19][22] + xor_out[51][19][22] + xor_out[52][19][22] + xor_out[53][19][22] + xor_out[54][19][22];
assign sum_out[11][19][22] = xor_out[55][19][22] + xor_out[56][19][22] + xor_out[57][19][22] + xor_out[58][19][22] + xor_out[59][19][22];
assign sum_out[12][19][22] = xor_out[60][19][22] + xor_out[61][19][22] + xor_out[62][19][22] + xor_out[63][19][22] + xor_out[64][19][22];
assign sum_out[13][19][22] = xor_out[65][19][22] + xor_out[66][19][22] + xor_out[67][19][22] + xor_out[68][19][22] + xor_out[69][19][22];
assign sum_out[14][19][22] = xor_out[70][19][22] + xor_out[71][19][22] + xor_out[72][19][22] + xor_out[73][19][22] + xor_out[74][19][22];
assign sum_out[15][19][22] = xor_out[75][19][22] + xor_out[76][19][22] + xor_out[77][19][22] + xor_out[78][19][22] + xor_out[79][19][22];
assign sum_out[16][19][22] = xor_out[80][19][22] + xor_out[81][19][22] + xor_out[82][19][22] + xor_out[83][19][22] + xor_out[84][19][22];
assign sum_out[17][19][22] = xor_out[85][19][22] + xor_out[86][19][22] + xor_out[87][19][22] + xor_out[88][19][22] + xor_out[89][19][22];
assign sum_out[18][19][22] = xor_out[90][19][22] + xor_out[91][19][22] + xor_out[92][19][22] + xor_out[93][19][22] + xor_out[94][19][22];
assign sum_out[19][19][22] = xor_out[95][19][22] + xor_out[96][19][22] + xor_out[97][19][22] + xor_out[98][19][22] + xor_out[99][19][22];

assign sum_out[0][19][23] = xor_out[0][19][23] + xor_out[1][19][23] + xor_out[2][19][23] + xor_out[3][19][23] + xor_out[4][19][23];
assign sum_out[1][19][23] = xor_out[5][19][23] + xor_out[6][19][23] + xor_out[7][19][23] + xor_out[8][19][23] + xor_out[9][19][23];
assign sum_out[2][19][23] = xor_out[10][19][23] + xor_out[11][19][23] + xor_out[12][19][23] + xor_out[13][19][23] + xor_out[14][19][23];
assign sum_out[3][19][23] = xor_out[15][19][23] + xor_out[16][19][23] + xor_out[17][19][23] + xor_out[18][19][23] + xor_out[19][19][23];
assign sum_out[4][19][23] = xor_out[20][19][23] + xor_out[21][19][23] + xor_out[22][19][23] + xor_out[23][19][23] + xor_out[24][19][23];
assign sum_out[5][19][23] = xor_out[25][19][23] + xor_out[26][19][23] + xor_out[27][19][23] + xor_out[28][19][23] + xor_out[29][19][23];
assign sum_out[6][19][23] = xor_out[30][19][23] + xor_out[31][19][23] + xor_out[32][19][23] + xor_out[33][19][23] + xor_out[34][19][23];
assign sum_out[7][19][23] = xor_out[35][19][23] + xor_out[36][19][23] + xor_out[37][19][23] + xor_out[38][19][23] + xor_out[39][19][23];
assign sum_out[8][19][23] = xor_out[40][19][23] + xor_out[41][19][23] + xor_out[42][19][23] + xor_out[43][19][23] + xor_out[44][19][23];
assign sum_out[9][19][23] = xor_out[45][19][23] + xor_out[46][19][23] + xor_out[47][19][23] + xor_out[48][19][23] + xor_out[49][19][23];
assign sum_out[10][19][23] = xor_out[50][19][23] + xor_out[51][19][23] + xor_out[52][19][23] + xor_out[53][19][23] + xor_out[54][19][23];
assign sum_out[11][19][23] = xor_out[55][19][23] + xor_out[56][19][23] + xor_out[57][19][23] + xor_out[58][19][23] + xor_out[59][19][23];
assign sum_out[12][19][23] = xor_out[60][19][23] + xor_out[61][19][23] + xor_out[62][19][23] + xor_out[63][19][23] + xor_out[64][19][23];
assign sum_out[13][19][23] = xor_out[65][19][23] + xor_out[66][19][23] + xor_out[67][19][23] + xor_out[68][19][23] + xor_out[69][19][23];
assign sum_out[14][19][23] = xor_out[70][19][23] + xor_out[71][19][23] + xor_out[72][19][23] + xor_out[73][19][23] + xor_out[74][19][23];
assign sum_out[15][19][23] = xor_out[75][19][23] + xor_out[76][19][23] + xor_out[77][19][23] + xor_out[78][19][23] + xor_out[79][19][23];
assign sum_out[16][19][23] = xor_out[80][19][23] + xor_out[81][19][23] + xor_out[82][19][23] + xor_out[83][19][23] + xor_out[84][19][23];
assign sum_out[17][19][23] = xor_out[85][19][23] + xor_out[86][19][23] + xor_out[87][19][23] + xor_out[88][19][23] + xor_out[89][19][23];
assign sum_out[18][19][23] = xor_out[90][19][23] + xor_out[91][19][23] + xor_out[92][19][23] + xor_out[93][19][23] + xor_out[94][19][23];
assign sum_out[19][19][23] = xor_out[95][19][23] + xor_out[96][19][23] + xor_out[97][19][23] + xor_out[98][19][23] + xor_out[99][19][23];

assign sum_out[0][20][0] = xor_out[0][20][0] + xor_out[1][20][0] + xor_out[2][20][0] + xor_out[3][20][0] + xor_out[4][20][0];
assign sum_out[1][20][0] = xor_out[5][20][0] + xor_out[6][20][0] + xor_out[7][20][0] + xor_out[8][20][0] + xor_out[9][20][0];
assign sum_out[2][20][0] = xor_out[10][20][0] + xor_out[11][20][0] + xor_out[12][20][0] + xor_out[13][20][0] + xor_out[14][20][0];
assign sum_out[3][20][0] = xor_out[15][20][0] + xor_out[16][20][0] + xor_out[17][20][0] + xor_out[18][20][0] + xor_out[19][20][0];
assign sum_out[4][20][0] = xor_out[20][20][0] + xor_out[21][20][0] + xor_out[22][20][0] + xor_out[23][20][0] + xor_out[24][20][0];
assign sum_out[5][20][0] = xor_out[25][20][0] + xor_out[26][20][0] + xor_out[27][20][0] + xor_out[28][20][0] + xor_out[29][20][0];
assign sum_out[6][20][0] = xor_out[30][20][0] + xor_out[31][20][0] + xor_out[32][20][0] + xor_out[33][20][0] + xor_out[34][20][0];
assign sum_out[7][20][0] = xor_out[35][20][0] + xor_out[36][20][0] + xor_out[37][20][0] + xor_out[38][20][0] + xor_out[39][20][0];
assign sum_out[8][20][0] = xor_out[40][20][0] + xor_out[41][20][0] + xor_out[42][20][0] + xor_out[43][20][0] + xor_out[44][20][0];
assign sum_out[9][20][0] = xor_out[45][20][0] + xor_out[46][20][0] + xor_out[47][20][0] + xor_out[48][20][0] + xor_out[49][20][0];
assign sum_out[10][20][0] = xor_out[50][20][0] + xor_out[51][20][0] + xor_out[52][20][0] + xor_out[53][20][0] + xor_out[54][20][0];
assign sum_out[11][20][0] = xor_out[55][20][0] + xor_out[56][20][0] + xor_out[57][20][0] + xor_out[58][20][0] + xor_out[59][20][0];
assign sum_out[12][20][0] = xor_out[60][20][0] + xor_out[61][20][0] + xor_out[62][20][0] + xor_out[63][20][0] + xor_out[64][20][0];
assign sum_out[13][20][0] = xor_out[65][20][0] + xor_out[66][20][0] + xor_out[67][20][0] + xor_out[68][20][0] + xor_out[69][20][0];
assign sum_out[14][20][0] = xor_out[70][20][0] + xor_out[71][20][0] + xor_out[72][20][0] + xor_out[73][20][0] + xor_out[74][20][0];
assign sum_out[15][20][0] = xor_out[75][20][0] + xor_out[76][20][0] + xor_out[77][20][0] + xor_out[78][20][0] + xor_out[79][20][0];
assign sum_out[16][20][0] = xor_out[80][20][0] + xor_out[81][20][0] + xor_out[82][20][0] + xor_out[83][20][0] + xor_out[84][20][0];
assign sum_out[17][20][0] = xor_out[85][20][0] + xor_out[86][20][0] + xor_out[87][20][0] + xor_out[88][20][0] + xor_out[89][20][0];
assign sum_out[18][20][0] = xor_out[90][20][0] + xor_out[91][20][0] + xor_out[92][20][0] + xor_out[93][20][0] + xor_out[94][20][0];
assign sum_out[19][20][0] = xor_out[95][20][0] + xor_out[96][20][0] + xor_out[97][20][0] + xor_out[98][20][0] + xor_out[99][20][0];

assign sum_out[0][20][1] = xor_out[0][20][1] + xor_out[1][20][1] + xor_out[2][20][1] + xor_out[3][20][1] + xor_out[4][20][1];
assign sum_out[1][20][1] = xor_out[5][20][1] + xor_out[6][20][1] + xor_out[7][20][1] + xor_out[8][20][1] + xor_out[9][20][1];
assign sum_out[2][20][1] = xor_out[10][20][1] + xor_out[11][20][1] + xor_out[12][20][1] + xor_out[13][20][1] + xor_out[14][20][1];
assign sum_out[3][20][1] = xor_out[15][20][1] + xor_out[16][20][1] + xor_out[17][20][1] + xor_out[18][20][1] + xor_out[19][20][1];
assign sum_out[4][20][1] = xor_out[20][20][1] + xor_out[21][20][1] + xor_out[22][20][1] + xor_out[23][20][1] + xor_out[24][20][1];
assign sum_out[5][20][1] = xor_out[25][20][1] + xor_out[26][20][1] + xor_out[27][20][1] + xor_out[28][20][1] + xor_out[29][20][1];
assign sum_out[6][20][1] = xor_out[30][20][1] + xor_out[31][20][1] + xor_out[32][20][1] + xor_out[33][20][1] + xor_out[34][20][1];
assign sum_out[7][20][1] = xor_out[35][20][1] + xor_out[36][20][1] + xor_out[37][20][1] + xor_out[38][20][1] + xor_out[39][20][1];
assign sum_out[8][20][1] = xor_out[40][20][1] + xor_out[41][20][1] + xor_out[42][20][1] + xor_out[43][20][1] + xor_out[44][20][1];
assign sum_out[9][20][1] = xor_out[45][20][1] + xor_out[46][20][1] + xor_out[47][20][1] + xor_out[48][20][1] + xor_out[49][20][1];
assign sum_out[10][20][1] = xor_out[50][20][1] + xor_out[51][20][1] + xor_out[52][20][1] + xor_out[53][20][1] + xor_out[54][20][1];
assign sum_out[11][20][1] = xor_out[55][20][1] + xor_out[56][20][1] + xor_out[57][20][1] + xor_out[58][20][1] + xor_out[59][20][1];
assign sum_out[12][20][1] = xor_out[60][20][1] + xor_out[61][20][1] + xor_out[62][20][1] + xor_out[63][20][1] + xor_out[64][20][1];
assign sum_out[13][20][1] = xor_out[65][20][1] + xor_out[66][20][1] + xor_out[67][20][1] + xor_out[68][20][1] + xor_out[69][20][1];
assign sum_out[14][20][1] = xor_out[70][20][1] + xor_out[71][20][1] + xor_out[72][20][1] + xor_out[73][20][1] + xor_out[74][20][1];
assign sum_out[15][20][1] = xor_out[75][20][1] + xor_out[76][20][1] + xor_out[77][20][1] + xor_out[78][20][1] + xor_out[79][20][1];
assign sum_out[16][20][1] = xor_out[80][20][1] + xor_out[81][20][1] + xor_out[82][20][1] + xor_out[83][20][1] + xor_out[84][20][1];
assign sum_out[17][20][1] = xor_out[85][20][1] + xor_out[86][20][1] + xor_out[87][20][1] + xor_out[88][20][1] + xor_out[89][20][1];
assign sum_out[18][20][1] = xor_out[90][20][1] + xor_out[91][20][1] + xor_out[92][20][1] + xor_out[93][20][1] + xor_out[94][20][1];
assign sum_out[19][20][1] = xor_out[95][20][1] + xor_out[96][20][1] + xor_out[97][20][1] + xor_out[98][20][1] + xor_out[99][20][1];

assign sum_out[0][20][2] = xor_out[0][20][2] + xor_out[1][20][2] + xor_out[2][20][2] + xor_out[3][20][2] + xor_out[4][20][2];
assign sum_out[1][20][2] = xor_out[5][20][2] + xor_out[6][20][2] + xor_out[7][20][2] + xor_out[8][20][2] + xor_out[9][20][2];
assign sum_out[2][20][2] = xor_out[10][20][2] + xor_out[11][20][2] + xor_out[12][20][2] + xor_out[13][20][2] + xor_out[14][20][2];
assign sum_out[3][20][2] = xor_out[15][20][2] + xor_out[16][20][2] + xor_out[17][20][2] + xor_out[18][20][2] + xor_out[19][20][2];
assign sum_out[4][20][2] = xor_out[20][20][2] + xor_out[21][20][2] + xor_out[22][20][2] + xor_out[23][20][2] + xor_out[24][20][2];
assign sum_out[5][20][2] = xor_out[25][20][2] + xor_out[26][20][2] + xor_out[27][20][2] + xor_out[28][20][2] + xor_out[29][20][2];
assign sum_out[6][20][2] = xor_out[30][20][2] + xor_out[31][20][2] + xor_out[32][20][2] + xor_out[33][20][2] + xor_out[34][20][2];
assign sum_out[7][20][2] = xor_out[35][20][2] + xor_out[36][20][2] + xor_out[37][20][2] + xor_out[38][20][2] + xor_out[39][20][2];
assign sum_out[8][20][2] = xor_out[40][20][2] + xor_out[41][20][2] + xor_out[42][20][2] + xor_out[43][20][2] + xor_out[44][20][2];
assign sum_out[9][20][2] = xor_out[45][20][2] + xor_out[46][20][2] + xor_out[47][20][2] + xor_out[48][20][2] + xor_out[49][20][2];
assign sum_out[10][20][2] = xor_out[50][20][2] + xor_out[51][20][2] + xor_out[52][20][2] + xor_out[53][20][2] + xor_out[54][20][2];
assign sum_out[11][20][2] = xor_out[55][20][2] + xor_out[56][20][2] + xor_out[57][20][2] + xor_out[58][20][2] + xor_out[59][20][2];
assign sum_out[12][20][2] = xor_out[60][20][2] + xor_out[61][20][2] + xor_out[62][20][2] + xor_out[63][20][2] + xor_out[64][20][2];
assign sum_out[13][20][2] = xor_out[65][20][2] + xor_out[66][20][2] + xor_out[67][20][2] + xor_out[68][20][2] + xor_out[69][20][2];
assign sum_out[14][20][2] = xor_out[70][20][2] + xor_out[71][20][2] + xor_out[72][20][2] + xor_out[73][20][2] + xor_out[74][20][2];
assign sum_out[15][20][2] = xor_out[75][20][2] + xor_out[76][20][2] + xor_out[77][20][2] + xor_out[78][20][2] + xor_out[79][20][2];
assign sum_out[16][20][2] = xor_out[80][20][2] + xor_out[81][20][2] + xor_out[82][20][2] + xor_out[83][20][2] + xor_out[84][20][2];
assign sum_out[17][20][2] = xor_out[85][20][2] + xor_out[86][20][2] + xor_out[87][20][2] + xor_out[88][20][2] + xor_out[89][20][2];
assign sum_out[18][20][2] = xor_out[90][20][2] + xor_out[91][20][2] + xor_out[92][20][2] + xor_out[93][20][2] + xor_out[94][20][2];
assign sum_out[19][20][2] = xor_out[95][20][2] + xor_out[96][20][2] + xor_out[97][20][2] + xor_out[98][20][2] + xor_out[99][20][2];

assign sum_out[0][20][3] = xor_out[0][20][3] + xor_out[1][20][3] + xor_out[2][20][3] + xor_out[3][20][3] + xor_out[4][20][3];
assign sum_out[1][20][3] = xor_out[5][20][3] + xor_out[6][20][3] + xor_out[7][20][3] + xor_out[8][20][3] + xor_out[9][20][3];
assign sum_out[2][20][3] = xor_out[10][20][3] + xor_out[11][20][3] + xor_out[12][20][3] + xor_out[13][20][3] + xor_out[14][20][3];
assign sum_out[3][20][3] = xor_out[15][20][3] + xor_out[16][20][3] + xor_out[17][20][3] + xor_out[18][20][3] + xor_out[19][20][3];
assign sum_out[4][20][3] = xor_out[20][20][3] + xor_out[21][20][3] + xor_out[22][20][3] + xor_out[23][20][3] + xor_out[24][20][3];
assign sum_out[5][20][3] = xor_out[25][20][3] + xor_out[26][20][3] + xor_out[27][20][3] + xor_out[28][20][3] + xor_out[29][20][3];
assign sum_out[6][20][3] = xor_out[30][20][3] + xor_out[31][20][3] + xor_out[32][20][3] + xor_out[33][20][3] + xor_out[34][20][3];
assign sum_out[7][20][3] = xor_out[35][20][3] + xor_out[36][20][3] + xor_out[37][20][3] + xor_out[38][20][3] + xor_out[39][20][3];
assign sum_out[8][20][3] = xor_out[40][20][3] + xor_out[41][20][3] + xor_out[42][20][3] + xor_out[43][20][3] + xor_out[44][20][3];
assign sum_out[9][20][3] = xor_out[45][20][3] + xor_out[46][20][3] + xor_out[47][20][3] + xor_out[48][20][3] + xor_out[49][20][3];
assign sum_out[10][20][3] = xor_out[50][20][3] + xor_out[51][20][3] + xor_out[52][20][3] + xor_out[53][20][3] + xor_out[54][20][3];
assign sum_out[11][20][3] = xor_out[55][20][3] + xor_out[56][20][3] + xor_out[57][20][3] + xor_out[58][20][3] + xor_out[59][20][3];
assign sum_out[12][20][3] = xor_out[60][20][3] + xor_out[61][20][3] + xor_out[62][20][3] + xor_out[63][20][3] + xor_out[64][20][3];
assign sum_out[13][20][3] = xor_out[65][20][3] + xor_out[66][20][3] + xor_out[67][20][3] + xor_out[68][20][3] + xor_out[69][20][3];
assign sum_out[14][20][3] = xor_out[70][20][3] + xor_out[71][20][3] + xor_out[72][20][3] + xor_out[73][20][3] + xor_out[74][20][3];
assign sum_out[15][20][3] = xor_out[75][20][3] + xor_out[76][20][3] + xor_out[77][20][3] + xor_out[78][20][3] + xor_out[79][20][3];
assign sum_out[16][20][3] = xor_out[80][20][3] + xor_out[81][20][3] + xor_out[82][20][3] + xor_out[83][20][3] + xor_out[84][20][3];
assign sum_out[17][20][3] = xor_out[85][20][3] + xor_out[86][20][3] + xor_out[87][20][3] + xor_out[88][20][3] + xor_out[89][20][3];
assign sum_out[18][20][3] = xor_out[90][20][3] + xor_out[91][20][3] + xor_out[92][20][3] + xor_out[93][20][3] + xor_out[94][20][3];
assign sum_out[19][20][3] = xor_out[95][20][3] + xor_out[96][20][3] + xor_out[97][20][3] + xor_out[98][20][3] + xor_out[99][20][3];

assign sum_out[0][20][4] = xor_out[0][20][4] + xor_out[1][20][4] + xor_out[2][20][4] + xor_out[3][20][4] + xor_out[4][20][4];
assign sum_out[1][20][4] = xor_out[5][20][4] + xor_out[6][20][4] + xor_out[7][20][4] + xor_out[8][20][4] + xor_out[9][20][4];
assign sum_out[2][20][4] = xor_out[10][20][4] + xor_out[11][20][4] + xor_out[12][20][4] + xor_out[13][20][4] + xor_out[14][20][4];
assign sum_out[3][20][4] = xor_out[15][20][4] + xor_out[16][20][4] + xor_out[17][20][4] + xor_out[18][20][4] + xor_out[19][20][4];
assign sum_out[4][20][4] = xor_out[20][20][4] + xor_out[21][20][4] + xor_out[22][20][4] + xor_out[23][20][4] + xor_out[24][20][4];
assign sum_out[5][20][4] = xor_out[25][20][4] + xor_out[26][20][4] + xor_out[27][20][4] + xor_out[28][20][4] + xor_out[29][20][4];
assign sum_out[6][20][4] = xor_out[30][20][4] + xor_out[31][20][4] + xor_out[32][20][4] + xor_out[33][20][4] + xor_out[34][20][4];
assign sum_out[7][20][4] = xor_out[35][20][4] + xor_out[36][20][4] + xor_out[37][20][4] + xor_out[38][20][4] + xor_out[39][20][4];
assign sum_out[8][20][4] = xor_out[40][20][4] + xor_out[41][20][4] + xor_out[42][20][4] + xor_out[43][20][4] + xor_out[44][20][4];
assign sum_out[9][20][4] = xor_out[45][20][4] + xor_out[46][20][4] + xor_out[47][20][4] + xor_out[48][20][4] + xor_out[49][20][4];
assign sum_out[10][20][4] = xor_out[50][20][4] + xor_out[51][20][4] + xor_out[52][20][4] + xor_out[53][20][4] + xor_out[54][20][4];
assign sum_out[11][20][4] = xor_out[55][20][4] + xor_out[56][20][4] + xor_out[57][20][4] + xor_out[58][20][4] + xor_out[59][20][4];
assign sum_out[12][20][4] = xor_out[60][20][4] + xor_out[61][20][4] + xor_out[62][20][4] + xor_out[63][20][4] + xor_out[64][20][4];
assign sum_out[13][20][4] = xor_out[65][20][4] + xor_out[66][20][4] + xor_out[67][20][4] + xor_out[68][20][4] + xor_out[69][20][4];
assign sum_out[14][20][4] = xor_out[70][20][4] + xor_out[71][20][4] + xor_out[72][20][4] + xor_out[73][20][4] + xor_out[74][20][4];
assign sum_out[15][20][4] = xor_out[75][20][4] + xor_out[76][20][4] + xor_out[77][20][4] + xor_out[78][20][4] + xor_out[79][20][4];
assign sum_out[16][20][4] = xor_out[80][20][4] + xor_out[81][20][4] + xor_out[82][20][4] + xor_out[83][20][4] + xor_out[84][20][4];
assign sum_out[17][20][4] = xor_out[85][20][4] + xor_out[86][20][4] + xor_out[87][20][4] + xor_out[88][20][4] + xor_out[89][20][4];
assign sum_out[18][20][4] = xor_out[90][20][4] + xor_out[91][20][4] + xor_out[92][20][4] + xor_out[93][20][4] + xor_out[94][20][4];
assign sum_out[19][20][4] = xor_out[95][20][4] + xor_out[96][20][4] + xor_out[97][20][4] + xor_out[98][20][4] + xor_out[99][20][4];

assign sum_out[0][20][5] = xor_out[0][20][5] + xor_out[1][20][5] + xor_out[2][20][5] + xor_out[3][20][5] + xor_out[4][20][5];
assign sum_out[1][20][5] = xor_out[5][20][5] + xor_out[6][20][5] + xor_out[7][20][5] + xor_out[8][20][5] + xor_out[9][20][5];
assign sum_out[2][20][5] = xor_out[10][20][5] + xor_out[11][20][5] + xor_out[12][20][5] + xor_out[13][20][5] + xor_out[14][20][5];
assign sum_out[3][20][5] = xor_out[15][20][5] + xor_out[16][20][5] + xor_out[17][20][5] + xor_out[18][20][5] + xor_out[19][20][5];
assign sum_out[4][20][5] = xor_out[20][20][5] + xor_out[21][20][5] + xor_out[22][20][5] + xor_out[23][20][5] + xor_out[24][20][5];
assign sum_out[5][20][5] = xor_out[25][20][5] + xor_out[26][20][5] + xor_out[27][20][5] + xor_out[28][20][5] + xor_out[29][20][5];
assign sum_out[6][20][5] = xor_out[30][20][5] + xor_out[31][20][5] + xor_out[32][20][5] + xor_out[33][20][5] + xor_out[34][20][5];
assign sum_out[7][20][5] = xor_out[35][20][5] + xor_out[36][20][5] + xor_out[37][20][5] + xor_out[38][20][5] + xor_out[39][20][5];
assign sum_out[8][20][5] = xor_out[40][20][5] + xor_out[41][20][5] + xor_out[42][20][5] + xor_out[43][20][5] + xor_out[44][20][5];
assign sum_out[9][20][5] = xor_out[45][20][5] + xor_out[46][20][5] + xor_out[47][20][5] + xor_out[48][20][5] + xor_out[49][20][5];
assign sum_out[10][20][5] = xor_out[50][20][5] + xor_out[51][20][5] + xor_out[52][20][5] + xor_out[53][20][5] + xor_out[54][20][5];
assign sum_out[11][20][5] = xor_out[55][20][5] + xor_out[56][20][5] + xor_out[57][20][5] + xor_out[58][20][5] + xor_out[59][20][5];
assign sum_out[12][20][5] = xor_out[60][20][5] + xor_out[61][20][5] + xor_out[62][20][5] + xor_out[63][20][5] + xor_out[64][20][5];
assign sum_out[13][20][5] = xor_out[65][20][5] + xor_out[66][20][5] + xor_out[67][20][5] + xor_out[68][20][5] + xor_out[69][20][5];
assign sum_out[14][20][5] = xor_out[70][20][5] + xor_out[71][20][5] + xor_out[72][20][5] + xor_out[73][20][5] + xor_out[74][20][5];
assign sum_out[15][20][5] = xor_out[75][20][5] + xor_out[76][20][5] + xor_out[77][20][5] + xor_out[78][20][5] + xor_out[79][20][5];
assign sum_out[16][20][5] = xor_out[80][20][5] + xor_out[81][20][5] + xor_out[82][20][5] + xor_out[83][20][5] + xor_out[84][20][5];
assign sum_out[17][20][5] = xor_out[85][20][5] + xor_out[86][20][5] + xor_out[87][20][5] + xor_out[88][20][5] + xor_out[89][20][5];
assign sum_out[18][20][5] = xor_out[90][20][5] + xor_out[91][20][5] + xor_out[92][20][5] + xor_out[93][20][5] + xor_out[94][20][5];
assign sum_out[19][20][5] = xor_out[95][20][5] + xor_out[96][20][5] + xor_out[97][20][5] + xor_out[98][20][5] + xor_out[99][20][5];

assign sum_out[0][20][6] = xor_out[0][20][6] + xor_out[1][20][6] + xor_out[2][20][6] + xor_out[3][20][6] + xor_out[4][20][6];
assign sum_out[1][20][6] = xor_out[5][20][6] + xor_out[6][20][6] + xor_out[7][20][6] + xor_out[8][20][6] + xor_out[9][20][6];
assign sum_out[2][20][6] = xor_out[10][20][6] + xor_out[11][20][6] + xor_out[12][20][6] + xor_out[13][20][6] + xor_out[14][20][6];
assign sum_out[3][20][6] = xor_out[15][20][6] + xor_out[16][20][6] + xor_out[17][20][6] + xor_out[18][20][6] + xor_out[19][20][6];
assign sum_out[4][20][6] = xor_out[20][20][6] + xor_out[21][20][6] + xor_out[22][20][6] + xor_out[23][20][6] + xor_out[24][20][6];
assign sum_out[5][20][6] = xor_out[25][20][6] + xor_out[26][20][6] + xor_out[27][20][6] + xor_out[28][20][6] + xor_out[29][20][6];
assign sum_out[6][20][6] = xor_out[30][20][6] + xor_out[31][20][6] + xor_out[32][20][6] + xor_out[33][20][6] + xor_out[34][20][6];
assign sum_out[7][20][6] = xor_out[35][20][6] + xor_out[36][20][6] + xor_out[37][20][6] + xor_out[38][20][6] + xor_out[39][20][6];
assign sum_out[8][20][6] = xor_out[40][20][6] + xor_out[41][20][6] + xor_out[42][20][6] + xor_out[43][20][6] + xor_out[44][20][6];
assign sum_out[9][20][6] = xor_out[45][20][6] + xor_out[46][20][6] + xor_out[47][20][6] + xor_out[48][20][6] + xor_out[49][20][6];
assign sum_out[10][20][6] = xor_out[50][20][6] + xor_out[51][20][6] + xor_out[52][20][6] + xor_out[53][20][6] + xor_out[54][20][6];
assign sum_out[11][20][6] = xor_out[55][20][6] + xor_out[56][20][6] + xor_out[57][20][6] + xor_out[58][20][6] + xor_out[59][20][6];
assign sum_out[12][20][6] = xor_out[60][20][6] + xor_out[61][20][6] + xor_out[62][20][6] + xor_out[63][20][6] + xor_out[64][20][6];
assign sum_out[13][20][6] = xor_out[65][20][6] + xor_out[66][20][6] + xor_out[67][20][6] + xor_out[68][20][6] + xor_out[69][20][6];
assign sum_out[14][20][6] = xor_out[70][20][6] + xor_out[71][20][6] + xor_out[72][20][6] + xor_out[73][20][6] + xor_out[74][20][6];
assign sum_out[15][20][6] = xor_out[75][20][6] + xor_out[76][20][6] + xor_out[77][20][6] + xor_out[78][20][6] + xor_out[79][20][6];
assign sum_out[16][20][6] = xor_out[80][20][6] + xor_out[81][20][6] + xor_out[82][20][6] + xor_out[83][20][6] + xor_out[84][20][6];
assign sum_out[17][20][6] = xor_out[85][20][6] + xor_out[86][20][6] + xor_out[87][20][6] + xor_out[88][20][6] + xor_out[89][20][6];
assign sum_out[18][20][6] = xor_out[90][20][6] + xor_out[91][20][6] + xor_out[92][20][6] + xor_out[93][20][6] + xor_out[94][20][6];
assign sum_out[19][20][6] = xor_out[95][20][6] + xor_out[96][20][6] + xor_out[97][20][6] + xor_out[98][20][6] + xor_out[99][20][6];

assign sum_out[0][20][7] = xor_out[0][20][7] + xor_out[1][20][7] + xor_out[2][20][7] + xor_out[3][20][7] + xor_out[4][20][7];
assign sum_out[1][20][7] = xor_out[5][20][7] + xor_out[6][20][7] + xor_out[7][20][7] + xor_out[8][20][7] + xor_out[9][20][7];
assign sum_out[2][20][7] = xor_out[10][20][7] + xor_out[11][20][7] + xor_out[12][20][7] + xor_out[13][20][7] + xor_out[14][20][7];
assign sum_out[3][20][7] = xor_out[15][20][7] + xor_out[16][20][7] + xor_out[17][20][7] + xor_out[18][20][7] + xor_out[19][20][7];
assign sum_out[4][20][7] = xor_out[20][20][7] + xor_out[21][20][7] + xor_out[22][20][7] + xor_out[23][20][7] + xor_out[24][20][7];
assign sum_out[5][20][7] = xor_out[25][20][7] + xor_out[26][20][7] + xor_out[27][20][7] + xor_out[28][20][7] + xor_out[29][20][7];
assign sum_out[6][20][7] = xor_out[30][20][7] + xor_out[31][20][7] + xor_out[32][20][7] + xor_out[33][20][7] + xor_out[34][20][7];
assign sum_out[7][20][7] = xor_out[35][20][7] + xor_out[36][20][7] + xor_out[37][20][7] + xor_out[38][20][7] + xor_out[39][20][7];
assign sum_out[8][20][7] = xor_out[40][20][7] + xor_out[41][20][7] + xor_out[42][20][7] + xor_out[43][20][7] + xor_out[44][20][7];
assign sum_out[9][20][7] = xor_out[45][20][7] + xor_out[46][20][7] + xor_out[47][20][7] + xor_out[48][20][7] + xor_out[49][20][7];
assign sum_out[10][20][7] = xor_out[50][20][7] + xor_out[51][20][7] + xor_out[52][20][7] + xor_out[53][20][7] + xor_out[54][20][7];
assign sum_out[11][20][7] = xor_out[55][20][7] + xor_out[56][20][7] + xor_out[57][20][7] + xor_out[58][20][7] + xor_out[59][20][7];
assign sum_out[12][20][7] = xor_out[60][20][7] + xor_out[61][20][7] + xor_out[62][20][7] + xor_out[63][20][7] + xor_out[64][20][7];
assign sum_out[13][20][7] = xor_out[65][20][7] + xor_out[66][20][7] + xor_out[67][20][7] + xor_out[68][20][7] + xor_out[69][20][7];
assign sum_out[14][20][7] = xor_out[70][20][7] + xor_out[71][20][7] + xor_out[72][20][7] + xor_out[73][20][7] + xor_out[74][20][7];
assign sum_out[15][20][7] = xor_out[75][20][7] + xor_out[76][20][7] + xor_out[77][20][7] + xor_out[78][20][7] + xor_out[79][20][7];
assign sum_out[16][20][7] = xor_out[80][20][7] + xor_out[81][20][7] + xor_out[82][20][7] + xor_out[83][20][7] + xor_out[84][20][7];
assign sum_out[17][20][7] = xor_out[85][20][7] + xor_out[86][20][7] + xor_out[87][20][7] + xor_out[88][20][7] + xor_out[89][20][7];
assign sum_out[18][20][7] = xor_out[90][20][7] + xor_out[91][20][7] + xor_out[92][20][7] + xor_out[93][20][7] + xor_out[94][20][7];
assign sum_out[19][20][7] = xor_out[95][20][7] + xor_out[96][20][7] + xor_out[97][20][7] + xor_out[98][20][7] + xor_out[99][20][7];

assign sum_out[0][20][8] = xor_out[0][20][8] + xor_out[1][20][8] + xor_out[2][20][8] + xor_out[3][20][8] + xor_out[4][20][8];
assign sum_out[1][20][8] = xor_out[5][20][8] + xor_out[6][20][8] + xor_out[7][20][8] + xor_out[8][20][8] + xor_out[9][20][8];
assign sum_out[2][20][8] = xor_out[10][20][8] + xor_out[11][20][8] + xor_out[12][20][8] + xor_out[13][20][8] + xor_out[14][20][8];
assign sum_out[3][20][8] = xor_out[15][20][8] + xor_out[16][20][8] + xor_out[17][20][8] + xor_out[18][20][8] + xor_out[19][20][8];
assign sum_out[4][20][8] = xor_out[20][20][8] + xor_out[21][20][8] + xor_out[22][20][8] + xor_out[23][20][8] + xor_out[24][20][8];
assign sum_out[5][20][8] = xor_out[25][20][8] + xor_out[26][20][8] + xor_out[27][20][8] + xor_out[28][20][8] + xor_out[29][20][8];
assign sum_out[6][20][8] = xor_out[30][20][8] + xor_out[31][20][8] + xor_out[32][20][8] + xor_out[33][20][8] + xor_out[34][20][8];
assign sum_out[7][20][8] = xor_out[35][20][8] + xor_out[36][20][8] + xor_out[37][20][8] + xor_out[38][20][8] + xor_out[39][20][8];
assign sum_out[8][20][8] = xor_out[40][20][8] + xor_out[41][20][8] + xor_out[42][20][8] + xor_out[43][20][8] + xor_out[44][20][8];
assign sum_out[9][20][8] = xor_out[45][20][8] + xor_out[46][20][8] + xor_out[47][20][8] + xor_out[48][20][8] + xor_out[49][20][8];
assign sum_out[10][20][8] = xor_out[50][20][8] + xor_out[51][20][8] + xor_out[52][20][8] + xor_out[53][20][8] + xor_out[54][20][8];
assign sum_out[11][20][8] = xor_out[55][20][8] + xor_out[56][20][8] + xor_out[57][20][8] + xor_out[58][20][8] + xor_out[59][20][8];
assign sum_out[12][20][8] = xor_out[60][20][8] + xor_out[61][20][8] + xor_out[62][20][8] + xor_out[63][20][8] + xor_out[64][20][8];
assign sum_out[13][20][8] = xor_out[65][20][8] + xor_out[66][20][8] + xor_out[67][20][8] + xor_out[68][20][8] + xor_out[69][20][8];
assign sum_out[14][20][8] = xor_out[70][20][8] + xor_out[71][20][8] + xor_out[72][20][8] + xor_out[73][20][8] + xor_out[74][20][8];
assign sum_out[15][20][8] = xor_out[75][20][8] + xor_out[76][20][8] + xor_out[77][20][8] + xor_out[78][20][8] + xor_out[79][20][8];
assign sum_out[16][20][8] = xor_out[80][20][8] + xor_out[81][20][8] + xor_out[82][20][8] + xor_out[83][20][8] + xor_out[84][20][8];
assign sum_out[17][20][8] = xor_out[85][20][8] + xor_out[86][20][8] + xor_out[87][20][8] + xor_out[88][20][8] + xor_out[89][20][8];
assign sum_out[18][20][8] = xor_out[90][20][8] + xor_out[91][20][8] + xor_out[92][20][8] + xor_out[93][20][8] + xor_out[94][20][8];
assign sum_out[19][20][8] = xor_out[95][20][8] + xor_out[96][20][8] + xor_out[97][20][8] + xor_out[98][20][8] + xor_out[99][20][8];

assign sum_out[0][20][9] = xor_out[0][20][9] + xor_out[1][20][9] + xor_out[2][20][9] + xor_out[3][20][9] + xor_out[4][20][9];
assign sum_out[1][20][9] = xor_out[5][20][9] + xor_out[6][20][9] + xor_out[7][20][9] + xor_out[8][20][9] + xor_out[9][20][9];
assign sum_out[2][20][9] = xor_out[10][20][9] + xor_out[11][20][9] + xor_out[12][20][9] + xor_out[13][20][9] + xor_out[14][20][9];
assign sum_out[3][20][9] = xor_out[15][20][9] + xor_out[16][20][9] + xor_out[17][20][9] + xor_out[18][20][9] + xor_out[19][20][9];
assign sum_out[4][20][9] = xor_out[20][20][9] + xor_out[21][20][9] + xor_out[22][20][9] + xor_out[23][20][9] + xor_out[24][20][9];
assign sum_out[5][20][9] = xor_out[25][20][9] + xor_out[26][20][9] + xor_out[27][20][9] + xor_out[28][20][9] + xor_out[29][20][9];
assign sum_out[6][20][9] = xor_out[30][20][9] + xor_out[31][20][9] + xor_out[32][20][9] + xor_out[33][20][9] + xor_out[34][20][9];
assign sum_out[7][20][9] = xor_out[35][20][9] + xor_out[36][20][9] + xor_out[37][20][9] + xor_out[38][20][9] + xor_out[39][20][9];
assign sum_out[8][20][9] = xor_out[40][20][9] + xor_out[41][20][9] + xor_out[42][20][9] + xor_out[43][20][9] + xor_out[44][20][9];
assign sum_out[9][20][9] = xor_out[45][20][9] + xor_out[46][20][9] + xor_out[47][20][9] + xor_out[48][20][9] + xor_out[49][20][9];
assign sum_out[10][20][9] = xor_out[50][20][9] + xor_out[51][20][9] + xor_out[52][20][9] + xor_out[53][20][9] + xor_out[54][20][9];
assign sum_out[11][20][9] = xor_out[55][20][9] + xor_out[56][20][9] + xor_out[57][20][9] + xor_out[58][20][9] + xor_out[59][20][9];
assign sum_out[12][20][9] = xor_out[60][20][9] + xor_out[61][20][9] + xor_out[62][20][9] + xor_out[63][20][9] + xor_out[64][20][9];
assign sum_out[13][20][9] = xor_out[65][20][9] + xor_out[66][20][9] + xor_out[67][20][9] + xor_out[68][20][9] + xor_out[69][20][9];
assign sum_out[14][20][9] = xor_out[70][20][9] + xor_out[71][20][9] + xor_out[72][20][9] + xor_out[73][20][9] + xor_out[74][20][9];
assign sum_out[15][20][9] = xor_out[75][20][9] + xor_out[76][20][9] + xor_out[77][20][9] + xor_out[78][20][9] + xor_out[79][20][9];
assign sum_out[16][20][9] = xor_out[80][20][9] + xor_out[81][20][9] + xor_out[82][20][9] + xor_out[83][20][9] + xor_out[84][20][9];
assign sum_out[17][20][9] = xor_out[85][20][9] + xor_out[86][20][9] + xor_out[87][20][9] + xor_out[88][20][9] + xor_out[89][20][9];
assign sum_out[18][20][9] = xor_out[90][20][9] + xor_out[91][20][9] + xor_out[92][20][9] + xor_out[93][20][9] + xor_out[94][20][9];
assign sum_out[19][20][9] = xor_out[95][20][9] + xor_out[96][20][9] + xor_out[97][20][9] + xor_out[98][20][9] + xor_out[99][20][9];

assign sum_out[0][20][10] = xor_out[0][20][10] + xor_out[1][20][10] + xor_out[2][20][10] + xor_out[3][20][10] + xor_out[4][20][10];
assign sum_out[1][20][10] = xor_out[5][20][10] + xor_out[6][20][10] + xor_out[7][20][10] + xor_out[8][20][10] + xor_out[9][20][10];
assign sum_out[2][20][10] = xor_out[10][20][10] + xor_out[11][20][10] + xor_out[12][20][10] + xor_out[13][20][10] + xor_out[14][20][10];
assign sum_out[3][20][10] = xor_out[15][20][10] + xor_out[16][20][10] + xor_out[17][20][10] + xor_out[18][20][10] + xor_out[19][20][10];
assign sum_out[4][20][10] = xor_out[20][20][10] + xor_out[21][20][10] + xor_out[22][20][10] + xor_out[23][20][10] + xor_out[24][20][10];
assign sum_out[5][20][10] = xor_out[25][20][10] + xor_out[26][20][10] + xor_out[27][20][10] + xor_out[28][20][10] + xor_out[29][20][10];
assign sum_out[6][20][10] = xor_out[30][20][10] + xor_out[31][20][10] + xor_out[32][20][10] + xor_out[33][20][10] + xor_out[34][20][10];
assign sum_out[7][20][10] = xor_out[35][20][10] + xor_out[36][20][10] + xor_out[37][20][10] + xor_out[38][20][10] + xor_out[39][20][10];
assign sum_out[8][20][10] = xor_out[40][20][10] + xor_out[41][20][10] + xor_out[42][20][10] + xor_out[43][20][10] + xor_out[44][20][10];
assign sum_out[9][20][10] = xor_out[45][20][10] + xor_out[46][20][10] + xor_out[47][20][10] + xor_out[48][20][10] + xor_out[49][20][10];
assign sum_out[10][20][10] = xor_out[50][20][10] + xor_out[51][20][10] + xor_out[52][20][10] + xor_out[53][20][10] + xor_out[54][20][10];
assign sum_out[11][20][10] = xor_out[55][20][10] + xor_out[56][20][10] + xor_out[57][20][10] + xor_out[58][20][10] + xor_out[59][20][10];
assign sum_out[12][20][10] = xor_out[60][20][10] + xor_out[61][20][10] + xor_out[62][20][10] + xor_out[63][20][10] + xor_out[64][20][10];
assign sum_out[13][20][10] = xor_out[65][20][10] + xor_out[66][20][10] + xor_out[67][20][10] + xor_out[68][20][10] + xor_out[69][20][10];
assign sum_out[14][20][10] = xor_out[70][20][10] + xor_out[71][20][10] + xor_out[72][20][10] + xor_out[73][20][10] + xor_out[74][20][10];
assign sum_out[15][20][10] = xor_out[75][20][10] + xor_out[76][20][10] + xor_out[77][20][10] + xor_out[78][20][10] + xor_out[79][20][10];
assign sum_out[16][20][10] = xor_out[80][20][10] + xor_out[81][20][10] + xor_out[82][20][10] + xor_out[83][20][10] + xor_out[84][20][10];
assign sum_out[17][20][10] = xor_out[85][20][10] + xor_out[86][20][10] + xor_out[87][20][10] + xor_out[88][20][10] + xor_out[89][20][10];
assign sum_out[18][20][10] = xor_out[90][20][10] + xor_out[91][20][10] + xor_out[92][20][10] + xor_out[93][20][10] + xor_out[94][20][10];
assign sum_out[19][20][10] = xor_out[95][20][10] + xor_out[96][20][10] + xor_out[97][20][10] + xor_out[98][20][10] + xor_out[99][20][10];

assign sum_out[0][20][11] = xor_out[0][20][11] + xor_out[1][20][11] + xor_out[2][20][11] + xor_out[3][20][11] + xor_out[4][20][11];
assign sum_out[1][20][11] = xor_out[5][20][11] + xor_out[6][20][11] + xor_out[7][20][11] + xor_out[8][20][11] + xor_out[9][20][11];
assign sum_out[2][20][11] = xor_out[10][20][11] + xor_out[11][20][11] + xor_out[12][20][11] + xor_out[13][20][11] + xor_out[14][20][11];
assign sum_out[3][20][11] = xor_out[15][20][11] + xor_out[16][20][11] + xor_out[17][20][11] + xor_out[18][20][11] + xor_out[19][20][11];
assign sum_out[4][20][11] = xor_out[20][20][11] + xor_out[21][20][11] + xor_out[22][20][11] + xor_out[23][20][11] + xor_out[24][20][11];
assign sum_out[5][20][11] = xor_out[25][20][11] + xor_out[26][20][11] + xor_out[27][20][11] + xor_out[28][20][11] + xor_out[29][20][11];
assign sum_out[6][20][11] = xor_out[30][20][11] + xor_out[31][20][11] + xor_out[32][20][11] + xor_out[33][20][11] + xor_out[34][20][11];
assign sum_out[7][20][11] = xor_out[35][20][11] + xor_out[36][20][11] + xor_out[37][20][11] + xor_out[38][20][11] + xor_out[39][20][11];
assign sum_out[8][20][11] = xor_out[40][20][11] + xor_out[41][20][11] + xor_out[42][20][11] + xor_out[43][20][11] + xor_out[44][20][11];
assign sum_out[9][20][11] = xor_out[45][20][11] + xor_out[46][20][11] + xor_out[47][20][11] + xor_out[48][20][11] + xor_out[49][20][11];
assign sum_out[10][20][11] = xor_out[50][20][11] + xor_out[51][20][11] + xor_out[52][20][11] + xor_out[53][20][11] + xor_out[54][20][11];
assign sum_out[11][20][11] = xor_out[55][20][11] + xor_out[56][20][11] + xor_out[57][20][11] + xor_out[58][20][11] + xor_out[59][20][11];
assign sum_out[12][20][11] = xor_out[60][20][11] + xor_out[61][20][11] + xor_out[62][20][11] + xor_out[63][20][11] + xor_out[64][20][11];
assign sum_out[13][20][11] = xor_out[65][20][11] + xor_out[66][20][11] + xor_out[67][20][11] + xor_out[68][20][11] + xor_out[69][20][11];
assign sum_out[14][20][11] = xor_out[70][20][11] + xor_out[71][20][11] + xor_out[72][20][11] + xor_out[73][20][11] + xor_out[74][20][11];
assign sum_out[15][20][11] = xor_out[75][20][11] + xor_out[76][20][11] + xor_out[77][20][11] + xor_out[78][20][11] + xor_out[79][20][11];
assign sum_out[16][20][11] = xor_out[80][20][11] + xor_out[81][20][11] + xor_out[82][20][11] + xor_out[83][20][11] + xor_out[84][20][11];
assign sum_out[17][20][11] = xor_out[85][20][11] + xor_out[86][20][11] + xor_out[87][20][11] + xor_out[88][20][11] + xor_out[89][20][11];
assign sum_out[18][20][11] = xor_out[90][20][11] + xor_out[91][20][11] + xor_out[92][20][11] + xor_out[93][20][11] + xor_out[94][20][11];
assign sum_out[19][20][11] = xor_out[95][20][11] + xor_out[96][20][11] + xor_out[97][20][11] + xor_out[98][20][11] + xor_out[99][20][11];

assign sum_out[0][20][12] = xor_out[0][20][12] + xor_out[1][20][12] + xor_out[2][20][12] + xor_out[3][20][12] + xor_out[4][20][12];
assign sum_out[1][20][12] = xor_out[5][20][12] + xor_out[6][20][12] + xor_out[7][20][12] + xor_out[8][20][12] + xor_out[9][20][12];
assign sum_out[2][20][12] = xor_out[10][20][12] + xor_out[11][20][12] + xor_out[12][20][12] + xor_out[13][20][12] + xor_out[14][20][12];
assign sum_out[3][20][12] = xor_out[15][20][12] + xor_out[16][20][12] + xor_out[17][20][12] + xor_out[18][20][12] + xor_out[19][20][12];
assign sum_out[4][20][12] = xor_out[20][20][12] + xor_out[21][20][12] + xor_out[22][20][12] + xor_out[23][20][12] + xor_out[24][20][12];
assign sum_out[5][20][12] = xor_out[25][20][12] + xor_out[26][20][12] + xor_out[27][20][12] + xor_out[28][20][12] + xor_out[29][20][12];
assign sum_out[6][20][12] = xor_out[30][20][12] + xor_out[31][20][12] + xor_out[32][20][12] + xor_out[33][20][12] + xor_out[34][20][12];
assign sum_out[7][20][12] = xor_out[35][20][12] + xor_out[36][20][12] + xor_out[37][20][12] + xor_out[38][20][12] + xor_out[39][20][12];
assign sum_out[8][20][12] = xor_out[40][20][12] + xor_out[41][20][12] + xor_out[42][20][12] + xor_out[43][20][12] + xor_out[44][20][12];
assign sum_out[9][20][12] = xor_out[45][20][12] + xor_out[46][20][12] + xor_out[47][20][12] + xor_out[48][20][12] + xor_out[49][20][12];
assign sum_out[10][20][12] = xor_out[50][20][12] + xor_out[51][20][12] + xor_out[52][20][12] + xor_out[53][20][12] + xor_out[54][20][12];
assign sum_out[11][20][12] = xor_out[55][20][12] + xor_out[56][20][12] + xor_out[57][20][12] + xor_out[58][20][12] + xor_out[59][20][12];
assign sum_out[12][20][12] = xor_out[60][20][12] + xor_out[61][20][12] + xor_out[62][20][12] + xor_out[63][20][12] + xor_out[64][20][12];
assign sum_out[13][20][12] = xor_out[65][20][12] + xor_out[66][20][12] + xor_out[67][20][12] + xor_out[68][20][12] + xor_out[69][20][12];
assign sum_out[14][20][12] = xor_out[70][20][12] + xor_out[71][20][12] + xor_out[72][20][12] + xor_out[73][20][12] + xor_out[74][20][12];
assign sum_out[15][20][12] = xor_out[75][20][12] + xor_out[76][20][12] + xor_out[77][20][12] + xor_out[78][20][12] + xor_out[79][20][12];
assign sum_out[16][20][12] = xor_out[80][20][12] + xor_out[81][20][12] + xor_out[82][20][12] + xor_out[83][20][12] + xor_out[84][20][12];
assign sum_out[17][20][12] = xor_out[85][20][12] + xor_out[86][20][12] + xor_out[87][20][12] + xor_out[88][20][12] + xor_out[89][20][12];
assign sum_out[18][20][12] = xor_out[90][20][12] + xor_out[91][20][12] + xor_out[92][20][12] + xor_out[93][20][12] + xor_out[94][20][12];
assign sum_out[19][20][12] = xor_out[95][20][12] + xor_out[96][20][12] + xor_out[97][20][12] + xor_out[98][20][12] + xor_out[99][20][12];

assign sum_out[0][20][13] = xor_out[0][20][13] + xor_out[1][20][13] + xor_out[2][20][13] + xor_out[3][20][13] + xor_out[4][20][13];
assign sum_out[1][20][13] = xor_out[5][20][13] + xor_out[6][20][13] + xor_out[7][20][13] + xor_out[8][20][13] + xor_out[9][20][13];
assign sum_out[2][20][13] = xor_out[10][20][13] + xor_out[11][20][13] + xor_out[12][20][13] + xor_out[13][20][13] + xor_out[14][20][13];
assign sum_out[3][20][13] = xor_out[15][20][13] + xor_out[16][20][13] + xor_out[17][20][13] + xor_out[18][20][13] + xor_out[19][20][13];
assign sum_out[4][20][13] = xor_out[20][20][13] + xor_out[21][20][13] + xor_out[22][20][13] + xor_out[23][20][13] + xor_out[24][20][13];
assign sum_out[5][20][13] = xor_out[25][20][13] + xor_out[26][20][13] + xor_out[27][20][13] + xor_out[28][20][13] + xor_out[29][20][13];
assign sum_out[6][20][13] = xor_out[30][20][13] + xor_out[31][20][13] + xor_out[32][20][13] + xor_out[33][20][13] + xor_out[34][20][13];
assign sum_out[7][20][13] = xor_out[35][20][13] + xor_out[36][20][13] + xor_out[37][20][13] + xor_out[38][20][13] + xor_out[39][20][13];
assign sum_out[8][20][13] = xor_out[40][20][13] + xor_out[41][20][13] + xor_out[42][20][13] + xor_out[43][20][13] + xor_out[44][20][13];
assign sum_out[9][20][13] = xor_out[45][20][13] + xor_out[46][20][13] + xor_out[47][20][13] + xor_out[48][20][13] + xor_out[49][20][13];
assign sum_out[10][20][13] = xor_out[50][20][13] + xor_out[51][20][13] + xor_out[52][20][13] + xor_out[53][20][13] + xor_out[54][20][13];
assign sum_out[11][20][13] = xor_out[55][20][13] + xor_out[56][20][13] + xor_out[57][20][13] + xor_out[58][20][13] + xor_out[59][20][13];
assign sum_out[12][20][13] = xor_out[60][20][13] + xor_out[61][20][13] + xor_out[62][20][13] + xor_out[63][20][13] + xor_out[64][20][13];
assign sum_out[13][20][13] = xor_out[65][20][13] + xor_out[66][20][13] + xor_out[67][20][13] + xor_out[68][20][13] + xor_out[69][20][13];
assign sum_out[14][20][13] = xor_out[70][20][13] + xor_out[71][20][13] + xor_out[72][20][13] + xor_out[73][20][13] + xor_out[74][20][13];
assign sum_out[15][20][13] = xor_out[75][20][13] + xor_out[76][20][13] + xor_out[77][20][13] + xor_out[78][20][13] + xor_out[79][20][13];
assign sum_out[16][20][13] = xor_out[80][20][13] + xor_out[81][20][13] + xor_out[82][20][13] + xor_out[83][20][13] + xor_out[84][20][13];
assign sum_out[17][20][13] = xor_out[85][20][13] + xor_out[86][20][13] + xor_out[87][20][13] + xor_out[88][20][13] + xor_out[89][20][13];
assign sum_out[18][20][13] = xor_out[90][20][13] + xor_out[91][20][13] + xor_out[92][20][13] + xor_out[93][20][13] + xor_out[94][20][13];
assign sum_out[19][20][13] = xor_out[95][20][13] + xor_out[96][20][13] + xor_out[97][20][13] + xor_out[98][20][13] + xor_out[99][20][13];

assign sum_out[0][20][14] = xor_out[0][20][14] + xor_out[1][20][14] + xor_out[2][20][14] + xor_out[3][20][14] + xor_out[4][20][14];
assign sum_out[1][20][14] = xor_out[5][20][14] + xor_out[6][20][14] + xor_out[7][20][14] + xor_out[8][20][14] + xor_out[9][20][14];
assign sum_out[2][20][14] = xor_out[10][20][14] + xor_out[11][20][14] + xor_out[12][20][14] + xor_out[13][20][14] + xor_out[14][20][14];
assign sum_out[3][20][14] = xor_out[15][20][14] + xor_out[16][20][14] + xor_out[17][20][14] + xor_out[18][20][14] + xor_out[19][20][14];
assign sum_out[4][20][14] = xor_out[20][20][14] + xor_out[21][20][14] + xor_out[22][20][14] + xor_out[23][20][14] + xor_out[24][20][14];
assign sum_out[5][20][14] = xor_out[25][20][14] + xor_out[26][20][14] + xor_out[27][20][14] + xor_out[28][20][14] + xor_out[29][20][14];
assign sum_out[6][20][14] = xor_out[30][20][14] + xor_out[31][20][14] + xor_out[32][20][14] + xor_out[33][20][14] + xor_out[34][20][14];
assign sum_out[7][20][14] = xor_out[35][20][14] + xor_out[36][20][14] + xor_out[37][20][14] + xor_out[38][20][14] + xor_out[39][20][14];
assign sum_out[8][20][14] = xor_out[40][20][14] + xor_out[41][20][14] + xor_out[42][20][14] + xor_out[43][20][14] + xor_out[44][20][14];
assign sum_out[9][20][14] = xor_out[45][20][14] + xor_out[46][20][14] + xor_out[47][20][14] + xor_out[48][20][14] + xor_out[49][20][14];
assign sum_out[10][20][14] = xor_out[50][20][14] + xor_out[51][20][14] + xor_out[52][20][14] + xor_out[53][20][14] + xor_out[54][20][14];
assign sum_out[11][20][14] = xor_out[55][20][14] + xor_out[56][20][14] + xor_out[57][20][14] + xor_out[58][20][14] + xor_out[59][20][14];
assign sum_out[12][20][14] = xor_out[60][20][14] + xor_out[61][20][14] + xor_out[62][20][14] + xor_out[63][20][14] + xor_out[64][20][14];
assign sum_out[13][20][14] = xor_out[65][20][14] + xor_out[66][20][14] + xor_out[67][20][14] + xor_out[68][20][14] + xor_out[69][20][14];
assign sum_out[14][20][14] = xor_out[70][20][14] + xor_out[71][20][14] + xor_out[72][20][14] + xor_out[73][20][14] + xor_out[74][20][14];
assign sum_out[15][20][14] = xor_out[75][20][14] + xor_out[76][20][14] + xor_out[77][20][14] + xor_out[78][20][14] + xor_out[79][20][14];
assign sum_out[16][20][14] = xor_out[80][20][14] + xor_out[81][20][14] + xor_out[82][20][14] + xor_out[83][20][14] + xor_out[84][20][14];
assign sum_out[17][20][14] = xor_out[85][20][14] + xor_out[86][20][14] + xor_out[87][20][14] + xor_out[88][20][14] + xor_out[89][20][14];
assign sum_out[18][20][14] = xor_out[90][20][14] + xor_out[91][20][14] + xor_out[92][20][14] + xor_out[93][20][14] + xor_out[94][20][14];
assign sum_out[19][20][14] = xor_out[95][20][14] + xor_out[96][20][14] + xor_out[97][20][14] + xor_out[98][20][14] + xor_out[99][20][14];

assign sum_out[0][20][15] = xor_out[0][20][15] + xor_out[1][20][15] + xor_out[2][20][15] + xor_out[3][20][15] + xor_out[4][20][15];
assign sum_out[1][20][15] = xor_out[5][20][15] + xor_out[6][20][15] + xor_out[7][20][15] + xor_out[8][20][15] + xor_out[9][20][15];
assign sum_out[2][20][15] = xor_out[10][20][15] + xor_out[11][20][15] + xor_out[12][20][15] + xor_out[13][20][15] + xor_out[14][20][15];
assign sum_out[3][20][15] = xor_out[15][20][15] + xor_out[16][20][15] + xor_out[17][20][15] + xor_out[18][20][15] + xor_out[19][20][15];
assign sum_out[4][20][15] = xor_out[20][20][15] + xor_out[21][20][15] + xor_out[22][20][15] + xor_out[23][20][15] + xor_out[24][20][15];
assign sum_out[5][20][15] = xor_out[25][20][15] + xor_out[26][20][15] + xor_out[27][20][15] + xor_out[28][20][15] + xor_out[29][20][15];
assign sum_out[6][20][15] = xor_out[30][20][15] + xor_out[31][20][15] + xor_out[32][20][15] + xor_out[33][20][15] + xor_out[34][20][15];
assign sum_out[7][20][15] = xor_out[35][20][15] + xor_out[36][20][15] + xor_out[37][20][15] + xor_out[38][20][15] + xor_out[39][20][15];
assign sum_out[8][20][15] = xor_out[40][20][15] + xor_out[41][20][15] + xor_out[42][20][15] + xor_out[43][20][15] + xor_out[44][20][15];
assign sum_out[9][20][15] = xor_out[45][20][15] + xor_out[46][20][15] + xor_out[47][20][15] + xor_out[48][20][15] + xor_out[49][20][15];
assign sum_out[10][20][15] = xor_out[50][20][15] + xor_out[51][20][15] + xor_out[52][20][15] + xor_out[53][20][15] + xor_out[54][20][15];
assign sum_out[11][20][15] = xor_out[55][20][15] + xor_out[56][20][15] + xor_out[57][20][15] + xor_out[58][20][15] + xor_out[59][20][15];
assign sum_out[12][20][15] = xor_out[60][20][15] + xor_out[61][20][15] + xor_out[62][20][15] + xor_out[63][20][15] + xor_out[64][20][15];
assign sum_out[13][20][15] = xor_out[65][20][15] + xor_out[66][20][15] + xor_out[67][20][15] + xor_out[68][20][15] + xor_out[69][20][15];
assign sum_out[14][20][15] = xor_out[70][20][15] + xor_out[71][20][15] + xor_out[72][20][15] + xor_out[73][20][15] + xor_out[74][20][15];
assign sum_out[15][20][15] = xor_out[75][20][15] + xor_out[76][20][15] + xor_out[77][20][15] + xor_out[78][20][15] + xor_out[79][20][15];
assign sum_out[16][20][15] = xor_out[80][20][15] + xor_out[81][20][15] + xor_out[82][20][15] + xor_out[83][20][15] + xor_out[84][20][15];
assign sum_out[17][20][15] = xor_out[85][20][15] + xor_out[86][20][15] + xor_out[87][20][15] + xor_out[88][20][15] + xor_out[89][20][15];
assign sum_out[18][20][15] = xor_out[90][20][15] + xor_out[91][20][15] + xor_out[92][20][15] + xor_out[93][20][15] + xor_out[94][20][15];
assign sum_out[19][20][15] = xor_out[95][20][15] + xor_out[96][20][15] + xor_out[97][20][15] + xor_out[98][20][15] + xor_out[99][20][15];

assign sum_out[0][20][16] = xor_out[0][20][16] + xor_out[1][20][16] + xor_out[2][20][16] + xor_out[3][20][16] + xor_out[4][20][16];
assign sum_out[1][20][16] = xor_out[5][20][16] + xor_out[6][20][16] + xor_out[7][20][16] + xor_out[8][20][16] + xor_out[9][20][16];
assign sum_out[2][20][16] = xor_out[10][20][16] + xor_out[11][20][16] + xor_out[12][20][16] + xor_out[13][20][16] + xor_out[14][20][16];
assign sum_out[3][20][16] = xor_out[15][20][16] + xor_out[16][20][16] + xor_out[17][20][16] + xor_out[18][20][16] + xor_out[19][20][16];
assign sum_out[4][20][16] = xor_out[20][20][16] + xor_out[21][20][16] + xor_out[22][20][16] + xor_out[23][20][16] + xor_out[24][20][16];
assign sum_out[5][20][16] = xor_out[25][20][16] + xor_out[26][20][16] + xor_out[27][20][16] + xor_out[28][20][16] + xor_out[29][20][16];
assign sum_out[6][20][16] = xor_out[30][20][16] + xor_out[31][20][16] + xor_out[32][20][16] + xor_out[33][20][16] + xor_out[34][20][16];
assign sum_out[7][20][16] = xor_out[35][20][16] + xor_out[36][20][16] + xor_out[37][20][16] + xor_out[38][20][16] + xor_out[39][20][16];
assign sum_out[8][20][16] = xor_out[40][20][16] + xor_out[41][20][16] + xor_out[42][20][16] + xor_out[43][20][16] + xor_out[44][20][16];
assign sum_out[9][20][16] = xor_out[45][20][16] + xor_out[46][20][16] + xor_out[47][20][16] + xor_out[48][20][16] + xor_out[49][20][16];
assign sum_out[10][20][16] = xor_out[50][20][16] + xor_out[51][20][16] + xor_out[52][20][16] + xor_out[53][20][16] + xor_out[54][20][16];
assign sum_out[11][20][16] = xor_out[55][20][16] + xor_out[56][20][16] + xor_out[57][20][16] + xor_out[58][20][16] + xor_out[59][20][16];
assign sum_out[12][20][16] = xor_out[60][20][16] + xor_out[61][20][16] + xor_out[62][20][16] + xor_out[63][20][16] + xor_out[64][20][16];
assign sum_out[13][20][16] = xor_out[65][20][16] + xor_out[66][20][16] + xor_out[67][20][16] + xor_out[68][20][16] + xor_out[69][20][16];
assign sum_out[14][20][16] = xor_out[70][20][16] + xor_out[71][20][16] + xor_out[72][20][16] + xor_out[73][20][16] + xor_out[74][20][16];
assign sum_out[15][20][16] = xor_out[75][20][16] + xor_out[76][20][16] + xor_out[77][20][16] + xor_out[78][20][16] + xor_out[79][20][16];
assign sum_out[16][20][16] = xor_out[80][20][16] + xor_out[81][20][16] + xor_out[82][20][16] + xor_out[83][20][16] + xor_out[84][20][16];
assign sum_out[17][20][16] = xor_out[85][20][16] + xor_out[86][20][16] + xor_out[87][20][16] + xor_out[88][20][16] + xor_out[89][20][16];
assign sum_out[18][20][16] = xor_out[90][20][16] + xor_out[91][20][16] + xor_out[92][20][16] + xor_out[93][20][16] + xor_out[94][20][16];
assign sum_out[19][20][16] = xor_out[95][20][16] + xor_out[96][20][16] + xor_out[97][20][16] + xor_out[98][20][16] + xor_out[99][20][16];

assign sum_out[0][20][17] = xor_out[0][20][17] + xor_out[1][20][17] + xor_out[2][20][17] + xor_out[3][20][17] + xor_out[4][20][17];
assign sum_out[1][20][17] = xor_out[5][20][17] + xor_out[6][20][17] + xor_out[7][20][17] + xor_out[8][20][17] + xor_out[9][20][17];
assign sum_out[2][20][17] = xor_out[10][20][17] + xor_out[11][20][17] + xor_out[12][20][17] + xor_out[13][20][17] + xor_out[14][20][17];
assign sum_out[3][20][17] = xor_out[15][20][17] + xor_out[16][20][17] + xor_out[17][20][17] + xor_out[18][20][17] + xor_out[19][20][17];
assign sum_out[4][20][17] = xor_out[20][20][17] + xor_out[21][20][17] + xor_out[22][20][17] + xor_out[23][20][17] + xor_out[24][20][17];
assign sum_out[5][20][17] = xor_out[25][20][17] + xor_out[26][20][17] + xor_out[27][20][17] + xor_out[28][20][17] + xor_out[29][20][17];
assign sum_out[6][20][17] = xor_out[30][20][17] + xor_out[31][20][17] + xor_out[32][20][17] + xor_out[33][20][17] + xor_out[34][20][17];
assign sum_out[7][20][17] = xor_out[35][20][17] + xor_out[36][20][17] + xor_out[37][20][17] + xor_out[38][20][17] + xor_out[39][20][17];
assign sum_out[8][20][17] = xor_out[40][20][17] + xor_out[41][20][17] + xor_out[42][20][17] + xor_out[43][20][17] + xor_out[44][20][17];
assign sum_out[9][20][17] = xor_out[45][20][17] + xor_out[46][20][17] + xor_out[47][20][17] + xor_out[48][20][17] + xor_out[49][20][17];
assign sum_out[10][20][17] = xor_out[50][20][17] + xor_out[51][20][17] + xor_out[52][20][17] + xor_out[53][20][17] + xor_out[54][20][17];
assign sum_out[11][20][17] = xor_out[55][20][17] + xor_out[56][20][17] + xor_out[57][20][17] + xor_out[58][20][17] + xor_out[59][20][17];
assign sum_out[12][20][17] = xor_out[60][20][17] + xor_out[61][20][17] + xor_out[62][20][17] + xor_out[63][20][17] + xor_out[64][20][17];
assign sum_out[13][20][17] = xor_out[65][20][17] + xor_out[66][20][17] + xor_out[67][20][17] + xor_out[68][20][17] + xor_out[69][20][17];
assign sum_out[14][20][17] = xor_out[70][20][17] + xor_out[71][20][17] + xor_out[72][20][17] + xor_out[73][20][17] + xor_out[74][20][17];
assign sum_out[15][20][17] = xor_out[75][20][17] + xor_out[76][20][17] + xor_out[77][20][17] + xor_out[78][20][17] + xor_out[79][20][17];
assign sum_out[16][20][17] = xor_out[80][20][17] + xor_out[81][20][17] + xor_out[82][20][17] + xor_out[83][20][17] + xor_out[84][20][17];
assign sum_out[17][20][17] = xor_out[85][20][17] + xor_out[86][20][17] + xor_out[87][20][17] + xor_out[88][20][17] + xor_out[89][20][17];
assign sum_out[18][20][17] = xor_out[90][20][17] + xor_out[91][20][17] + xor_out[92][20][17] + xor_out[93][20][17] + xor_out[94][20][17];
assign sum_out[19][20][17] = xor_out[95][20][17] + xor_out[96][20][17] + xor_out[97][20][17] + xor_out[98][20][17] + xor_out[99][20][17];

assign sum_out[0][20][18] = xor_out[0][20][18] + xor_out[1][20][18] + xor_out[2][20][18] + xor_out[3][20][18] + xor_out[4][20][18];
assign sum_out[1][20][18] = xor_out[5][20][18] + xor_out[6][20][18] + xor_out[7][20][18] + xor_out[8][20][18] + xor_out[9][20][18];
assign sum_out[2][20][18] = xor_out[10][20][18] + xor_out[11][20][18] + xor_out[12][20][18] + xor_out[13][20][18] + xor_out[14][20][18];
assign sum_out[3][20][18] = xor_out[15][20][18] + xor_out[16][20][18] + xor_out[17][20][18] + xor_out[18][20][18] + xor_out[19][20][18];
assign sum_out[4][20][18] = xor_out[20][20][18] + xor_out[21][20][18] + xor_out[22][20][18] + xor_out[23][20][18] + xor_out[24][20][18];
assign sum_out[5][20][18] = xor_out[25][20][18] + xor_out[26][20][18] + xor_out[27][20][18] + xor_out[28][20][18] + xor_out[29][20][18];
assign sum_out[6][20][18] = xor_out[30][20][18] + xor_out[31][20][18] + xor_out[32][20][18] + xor_out[33][20][18] + xor_out[34][20][18];
assign sum_out[7][20][18] = xor_out[35][20][18] + xor_out[36][20][18] + xor_out[37][20][18] + xor_out[38][20][18] + xor_out[39][20][18];
assign sum_out[8][20][18] = xor_out[40][20][18] + xor_out[41][20][18] + xor_out[42][20][18] + xor_out[43][20][18] + xor_out[44][20][18];
assign sum_out[9][20][18] = xor_out[45][20][18] + xor_out[46][20][18] + xor_out[47][20][18] + xor_out[48][20][18] + xor_out[49][20][18];
assign sum_out[10][20][18] = xor_out[50][20][18] + xor_out[51][20][18] + xor_out[52][20][18] + xor_out[53][20][18] + xor_out[54][20][18];
assign sum_out[11][20][18] = xor_out[55][20][18] + xor_out[56][20][18] + xor_out[57][20][18] + xor_out[58][20][18] + xor_out[59][20][18];
assign sum_out[12][20][18] = xor_out[60][20][18] + xor_out[61][20][18] + xor_out[62][20][18] + xor_out[63][20][18] + xor_out[64][20][18];
assign sum_out[13][20][18] = xor_out[65][20][18] + xor_out[66][20][18] + xor_out[67][20][18] + xor_out[68][20][18] + xor_out[69][20][18];
assign sum_out[14][20][18] = xor_out[70][20][18] + xor_out[71][20][18] + xor_out[72][20][18] + xor_out[73][20][18] + xor_out[74][20][18];
assign sum_out[15][20][18] = xor_out[75][20][18] + xor_out[76][20][18] + xor_out[77][20][18] + xor_out[78][20][18] + xor_out[79][20][18];
assign sum_out[16][20][18] = xor_out[80][20][18] + xor_out[81][20][18] + xor_out[82][20][18] + xor_out[83][20][18] + xor_out[84][20][18];
assign sum_out[17][20][18] = xor_out[85][20][18] + xor_out[86][20][18] + xor_out[87][20][18] + xor_out[88][20][18] + xor_out[89][20][18];
assign sum_out[18][20][18] = xor_out[90][20][18] + xor_out[91][20][18] + xor_out[92][20][18] + xor_out[93][20][18] + xor_out[94][20][18];
assign sum_out[19][20][18] = xor_out[95][20][18] + xor_out[96][20][18] + xor_out[97][20][18] + xor_out[98][20][18] + xor_out[99][20][18];

assign sum_out[0][20][19] = xor_out[0][20][19] + xor_out[1][20][19] + xor_out[2][20][19] + xor_out[3][20][19] + xor_out[4][20][19];
assign sum_out[1][20][19] = xor_out[5][20][19] + xor_out[6][20][19] + xor_out[7][20][19] + xor_out[8][20][19] + xor_out[9][20][19];
assign sum_out[2][20][19] = xor_out[10][20][19] + xor_out[11][20][19] + xor_out[12][20][19] + xor_out[13][20][19] + xor_out[14][20][19];
assign sum_out[3][20][19] = xor_out[15][20][19] + xor_out[16][20][19] + xor_out[17][20][19] + xor_out[18][20][19] + xor_out[19][20][19];
assign sum_out[4][20][19] = xor_out[20][20][19] + xor_out[21][20][19] + xor_out[22][20][19] + xor_out[23][20][19] + xor_out[24][20][19];
assign sum_out[5][20][19] = xor_out[25][20][19] + xor_out[26][20][19] + xor_out[27][20][19] + xor_out[28][20][19] + xor_out[29][20][19];
assign sum_out[6][20][19] = xor_out[30][20][19] + xor_out[31][20][19] + xor_out[32][20][19] + xor_out[33][20][19] + xor_out[34][20][19];
assign sum_out[7][20][19] = xor_out[35][20][19] + xor_out[36][20][19] + xor_out[37][20][19] + xor_out[38][20][19] + xor_out[39][20][19];
assign sum_out[8][20][19] = xor_out[40][20][19] + xor_out[41][20][19] + xor_out[42][20][19] + xor_out[43][20][19] + xor_out[44][20][19];
assign sum_out[9][20][19] = xor_out[45][20][19] + xor_out[46][20][19] + xor_out[47][20][19] + xor_out[48][20][19] + xor_out[49][20][19];
assign sum_out[10][20][19] = xor_out[50][20][19] + xor_out[51][20][19] + xor_out[52][20][19] + xor_out[53][20][19] + xor_out[54][20][19];
assign sum_out[11][20][19] = xor_out[55][20][19] + xor_out[56][20][19] + xor_out[57][20][19] + xor_out[58][20][19] + xor_out[59][20][19];
assign sum_out[12][20][19] = xor_out[60][20][19] + xor_out[61][20][19] + xor_out[62][20][19] + xor_out[63][20][19] + xor_out[64][20][19];
assign sum_out[13][20][19] = xor_out[65][20][19] + xor_out[66][20][19] + xor_out[67][20][19] + xor_out[68][20][19] + xor_out[69][20][19];
assign sum_out[14][20][19] = xor_out[70][20][19] + xor_out[71][20][19] + xor_out[72][20][19] + xor_out[73][20][19] + xor_out[74][20][19];
assign sum_out[15][20][19] = xor_out[75][20][19] + xor_out[76][20][19] + xor_out[77][20][19] + xor_out[78][20][19] + xor_out[79][20][19];
assign sum_out[16][20][19] = xor_out[80][20][19] + xor_out[81][20][19] + xor_out[82][20][19] + xor_out[83][20][19] + xor_out[84][20][19];
assign sum_out[17][20][19] = xor_out[85][20][19] + xor_out[86][20][19] + xor_out[87][20][19] + xor_out[88][20][19] + xor_out[89][20][19];
assign sum_out[18][20][19] = xor_out[90][20][19] + xor_out[91][20][19] + xor_out[92][20][19] + xor_out[93][20][19] + xor_out[94][20][19];
assign sum_out[19][20][19] = xor_out[95][20][19] + xor_out[96][20][19] + xor_out[97][20][19] + xor_out[98][20][19] + xor_out[99][20][19];

assign sum_out[0][20][20] = xor_out[0][20][20] + xor_out[1][20][20] + xor_out[2][20][20] + xor_out[3][20][20] + xor_out[4][20][20];
assign sum_out[1][20][20] = xor_out[5][20][20] + xor_out[6][20][20] + xor_out[7][20][20] + xor_out[8][20][20] + xor_out[9][20][20];
assign sum_out[2][20][20] = xor_out[10][20][20] + xor_out[11][20][20] + xor_out[12][20][20] + xor_out[13][20][20] + xor_out[14][20][20];
assign sum_out[3][20][20] = xor_out[15][20][20] + xor_out[16][20][20] + xor_out[17][20][20] + xor_out[18][20][20] + xor_out[19][20][20];
assign sum_out[4][20][20] = xor_out[20][20][20] + xor_out[21][20][20] + xor_out[22][20][20] + xor_out[23][20][20] + xor_out[24][20][20];
assign sum_out[5][20][20] = xor_out[25][20][20] + xor_out[26][20][20] + xor_out[27][20][20] + xor_out[28][20][20] + xor_out[29][20][20];
assign sum_out[6][20][20] = xor_out[30][20][20] + xor_out[31][20][20] + xor_out[32][20][20] + xor_out[33][20][20] + xor_out[34][20][20];
assign sum_out[7][20][20] = xor_out[35][20][20] + xor_out[36][20][20] + xor_out[37][20][20] + xor_out[38][20][20] + xor_out[39][20][20];
assign sum_out[8][20][20] = xor_out[40][20][20] + xor_out[41][20][20] + xor_out[42][20][20] + xor_out[43][20][20] + xor_out[44][20][20];
assign sum_out[9][20][20] = xor_out[45][20][20] + xor_out[46][20][20] + xor_out[47][20][20] + xor_out[48][20][20] + xor_out[49][20][20];
assign sum_out[10][20][20] = xor_out[50][20][20] + xor_out[51][20][20] + xor_out[52][20][20] + xor_out[53][20][20] + xor_out[54][20][20];
assign sum_out[11][20][20] = xor_out[55][20][20] + xor_out[56][20][20] + xor_out[57][20][20] + xor_out[58][20][20] + xor_out[59][20][20];
assign sum_out[12][20][20] = xor_out[60][20][20] + xor_out[61][20][20] + xor_out[62][20][20] + xor_out[63][20][20] + xor_out[64][20][20];
assign sum_out[13][20][20] = xor_out[65][20][20] + xor_out[66][20][20] + xor_out[67][20][20] + xor_out[68][20][20] + xor_out[69][20][20];
assign sum_out[14][20][20] = xor_out[70][20][20] + xor_out[71][20][20] + xor_out[72][20][20] + xor_out[73][20][20] + xor_out[74][20][20];
assign sum_out[15][20][20] = xor_out[75][20][20] + xor_out[76][20][20] + xor_out[77][20][20] + xor_out[78][20][20] + xor_out[79][20][20];
assign sum_out[16][20][20] = xor_out[80][20][20] + xor_out[81][20][20] + xor_out[82][20][20] + xor_out[83][20][20] + xor_out[84][20][20];
assign sum_out[17][20][20] = xor_out[85][20][20] + xor_out[86][20][20] + xor_out[87][20][20] + xor_out[88][20][20] + xor_out[89][20][20];
assign sum_out[18][20][20] = xor_out[90][20][20] + xor_out[91][20][20] + xor_out[92][20][20] + xor_out[93][20][20] + xor_out[94][20][20];
assign sum_out[19][20][20] = xor_out[95][20][20] + xor_out[96][20][20] + xor_out[97][20][20] + xor_out[98][20][20] + xor_out[99][20][20];

assign sum_out[0][20][21] = xor_out[0][20][21] + xor_out[1][20][21] + xor_out[2][20][21] + xor_out[3][20][21] + xor_out[4][20][21];
assign sum_out[1][20][21] = xor_out[5][20][21] + xor_out[6][20][21] + xor_out[7][20][21] + xor_out[8][20][21] + xor_out[9][20][21];
assign sum_out[2][20][21] = xor_out[10][20][21] + xor_out[11][20][21] + xor_out[12][20][21] + xor_out[13][20][21] + xor_out[14][20][21];
assign sum_out[3][20][21] = xor_out[15][20][21] + xor_out[16][20][21] + xor_out[17][20][21] + xor_out[18][20][21] + xor_out[19][20][21];
assign sum_out[4][20][21] = xor_out[20][20][21] + xor_out[21][20][21] + xor_out[22][20][21] + xor_out[23][20][21] + xor_out[24][20][21];
assign sum_out[5][20][21] = xor_out[25][20][21] + xor_out[26][20][21] + xor_out[27][20][21] + xor_out[28][20][21] + xor_out[29][20][21];
assign sum_out[6][20][21] = xor_out[30][20][21] + xor_out[31][20][21] + xor_out[32][20][21] + xor_out[33][20][21] + xor_out[34][20][21];
assign sum_out[7][20][21] = xor_out[35][20][21] + xor_out[36][20][21] + xor_out[37][20][21] + xor_out[38][20][21] + xor_out[39][20][21];
assign sum_out[8][20][21] = xor_out[40][20][21] + xor_out[41][20][21] + xor_out[42][20][21] + xor_out[43][20][21] + xor_out[44][20][21];
assign sum_out[9][20][21] = xor_out[45][20][21] + xor_out[46][20][21] + xor_out[47][20][21] + xor_out[48][20][21] + xor_out[49][20][21];
assign sum_out[10][20][21] = xor_out[50][20][21] + xor_out[51][20][21] + xor_out[52][20][21] + xor_out[53][20][21] + xor_out[54][20][21];
assign sum_out[11][20][21] = xor_out[55][20][21] + xor_out[56][20][21] + xor_out[57][20][21] + xor_out[58][20][21] + xor_out[59][20][21];
assign sum_out[12][20][21] = xor_out[60][20][21] + xor_out[61][20][21] + xor_out[62][20][21] + xor_out[63][20][21] + xor_out[64][20][21];
assign sum_out[13][20][21] = xor_out[65][20][21] + xor_out[66][20][21] + xor_out[67][20][21] + xor_out[68][20][21] + xor_out[69][20][21];
assign sum_out[14][20][21] = xor_out[70][20][21] + xor_out[71][20][21] + xor_out[72][20][21] + xor_out[73][20][21] + xor_out[74][20][21];
assign sum_out[15][20][21] = xor_out[75][20][21] + xor_out[76][20][21] + xor_out[77][20][21] + xor_out[78][20][21] + xor_out[79][20][21];
assign sum_out[16][20][21] = xor_out[80][20][21] + xor_out[81][20][21] + xor_out[82][20][21] + xor_out[83][20][21] + xor_out[84][20][21];
assign sum_out[17][20][21] = xor_out[85][20][21] + xor_out[86][20][21] + xor_out[87][20][21] + xor_out[88][20][21] + xor_out[89][20][21];
assign sum_out[18][20][21] = xor_out[90][20][21] + xor_out[91][20][21] + xor_out[92][20][21] + xor_out[93][20][21] + xor_out[94][20][21];
assign sum_out[19][20][21] = xor_out[95][20][21] + xor_out[96][20][21] + xor_out[97][20][21] + xor_out[98][20][21] + xor_out[99][20][21];

assign sum_out[0][20][22] = xor_out[0][20][22] + xor_out[1][20][22] + xor_out[2][20][22] + xor_out[3][20][22] + xor_out[4][20][22];
assign sum_out[1][20][22] = xor_out[5][20][22] + xor_out[6][20][22] + xor_out[7][20][22] + xor_out[8][20][22] + xor_out[9][20][22];
assign sum_out[2][20][22] = xor_out[10][20][22] + xor_out[11][20][22] + xor_out[12][20][22] + xor_out[13][20][22] + xor_out[14][20][22];
assign sum_out[3][20][22] = xor_out[15][20][22] + xor_out[16][20][22] + xor_out[17][20][22] + xor_out[18][20][22] + xor_out[19][20][22];
assign sum_out[4][20][22] = xor_out[20][20][22] + xor_out[21][20][22] + xor_out[22][20][22] + xor_out[23][20][22] + xor_out[24][20][22];
assign sum_out[5][20][22] = xor_out[25][20][22] + xor_out[26][20][22] + xor_out[27][20][22] + xor_out[28][20][22] + xor_out[29][20][22];
assign sum_out[6][20][22] = xor_out[30][20][22] + xor_out[31][20][22] + xor_out[32][20][22] + xor_out[33][20][22] + xor_out[34][20][22];
assign sum_out[7][20][22] = xor_out[35][20][22] + xor_out[36][20][22] + xor_out[37][20][22] + xor_out[38][20][22] + xor_out[39][20][22];
assign sum_out[8][20][22] = xor_out[40][20][22] + xor_out[41][20][22] + xor_out[42][20][22] + xor_out[43][20][22] + xor_out[44][20][22];
assign sum_out[9][20][22] = xor_out[45][20][22] + xor_out[46][20][22] + xor_out[47][20][22] + xor_out[48][20][22] + xor_out[49][20][22];
assign sum_out[10][20][22] = xor_out[50][20][22] + xor_out[51][20][22] + xor_out[52][20][22] + xor_out[53][20][22] + xor_out[54][20][22];
assign sum_out[11][20][22] = xor_out[55][20][22] + xor_out[56][20][22] + xor_out[57][20][22] + xor_out[58][20][22] + xor_out[59][20][22];
assign sum_out[12][20][22] = xor_out[60][20][22] + xor_out[61][20][22] + xor_out[62][20][22] + xor_out[63][20][22] + xor_out[64][20][22];
assign sum_out[13][20][22] = xor_out[65][20][22] + xor_out[66][20][22] + xor_out[67][20][22] + xor_out[68][20][22] + xor_out[69][20][22];
assign sum_out[14][20][22] = xor_out[70][20][22] + xor_out[71][20][22] + xor_out[72][20][22] + xor_out[73][20][22] + xor_out[74][20][22];
assign sum_out[15][20][22] = xor_out[75][20][22] + xor_out[76][20][22] + xor_out[77][20][22] + xor_out[78][20][22] + xor_out[79][20][22];
assign sum_out[16][20][22] = xor_out[80][20][22] + xor_out[81][20][22] + xor_out[82][20][22] + xor_out[83][20][22] + xor_out[84][20][22];
assign sum_out[17][20][22] = xor_out[85][20][22] + xor_out[86][20][22] + xor_out[87][20][22] + xor_out[88][20][22] + xor_out[89][20][22];
assign sum_out[18][20][22] = xor_out[90][20][22] + xor_out[91][20][22] + xor_out[92][20][22] + xor_out[93][20][22] + xor_out[94][20][22];
assign sum_out[19][20][22] = xor_out[95][20][22] + xor_out[96][20][22] + xor_out[97][20][22] + xor_out[98][20][22] + xor_out[99][20][22];

assign sum_out[0][20][23] = xor_out[0][20][23] + xor_out[1][20][23] + xor_out[2][20][23] + xor_out[3][20][23] + xor_out[4][20][23];
assign sum_out[1][20][23] = xor_out[5][20][23] + xor_out[6][20][23] + xor_out[7][20][23] + xor_out[8][20][23] + xor_out[9][20][23];
assign sum_out[2][20][23] = xor_out[10][20][23] + xor_out[11][20][23] + xor_out[12][20][23] + xor_out[13][20][23] + xor_out[14][20][23];
assign sum_out[3][20][23] = xor_out[15][20][23] + xor_out[16][20][23] + xor_out[17][20][23] + xor_out[18][20][23] + xor_out[19][20][23];
assign sum_out[4][20][23] = xor_out[20][20][23] + xor_out[21][20][23] + xor_out[22][20][23] + xor_out[23][20][23] + xor_out[24][20][23];
assign sum_out[5][20][23] = xor_out[25][20][23] + xor_out[26][20][23] + xor_out[27][20][23] + xor_out[28][20][23] + xor_out[29][20][23];
assign sum_out[6][20][23] = xor_out[30][20][23] + xor_out[31][20][23] + xor_out[32][20][23] + xor_out[33][20][23] + xor_out[34][20][23];
assign sum_out[7][20][23] = xor_out[35][20][23] + xor_out[36][20][23] + xor_out[37][20][23] + xor_out[38][20][23] + xor_out[39][20][23];
assign sum_out[8][20][23] = xor_out[40][20][23] + xor_out[41][20][23] + xor_out[42][20][23] + xor_out[43][20][23] + xor_out[44][20][23];
assign sum_out[9][20][23] = xor_out[45][20][23] + xor_out[46][20][23] + xor_out[47][20][23] + xor_out[48][20][23] + xor_out[49][20][23];
assign sum_out[10][20][23] = xor_out[50][20][23] + xor_out[51][20][23] + xor_out[52][20][23] + xor_out[53][20][23] + xor_out[54][20][23];
assign sum_out[11][20][23] = xor_out[55][20][23] + xor_out[56][20][23] + xor_out[57][20][23] + xor_out[58][20][23] + xor_out[59][20][23];
assign sum_out[12][20][23] = xor_out[60][20][23] + xor_out[61][20][23] + xor_out[62][20][23] + xor_out[63][20][23] + xor_out[64][20][23];
assign sum_out[13][20][23] = xor_out[65][20][23] + xor_out[66][20][23] + xor_out[67][20][23] + xor_out[68][20][23] + xor_out[69][20][23];
assign sum_out[14][20][23] = xor_out[70][20][23] + xor_out[71][20][23] + xor_out[72][20][23] + xor_out[73][20][23] + xor_out[74][20][23];
assign sum_out[15][20][23] = xor_out[75][20][23] + xor_out[76][20][23] + xor_out[77][20][23] + xor_out[78][20][23] + xor_out[79][20][23];
assign sum_out[16][20][23] = xor_out[80][20][23] + xor_out[81][20][23] + xor_out[82][20][23] + xor_out[83][20][23] + xor_out[84][20][23];
assign sum_out[17][20][23] = xor_out[85][20][23] + xor_out[86][20][23] + xor_out[87][20][23] + xor_out[88][20][23] + xor_out[89][20][23];
assign sum_out[18][20][23] = xor_out[90][20][23] + xor_out[91][20][23] + xor_out[92][20][23] + xor_out[93][20][23] + xor_out[94][20][23];
assign sum_out[19][20][23] = xor_out[95][20][23] + xor_out[96][20][23] + xor_out[97][20][23] + xor_out[98][20][23] + xor_out[99][20][23];

assign sum_out[0][21][0] = xor_out[0][21][0] + xor_out[1][21][0] + xor_out[2][21][0] + xor_out[3][21][0] + xor_out[4][21][0];
assign sum_out[1][21][0] = xor_out[5][21][0] + xor_out[6][21][0] + xor_out[7][21][0] + xor_out[8][21][0] + xor_out[9][21][0];
assign sum_out[2][21][0] = xor_out[10][21][0] + xor_out[11][21][0] + xor_out[12][21][0] + xor_out[13][21][0] + xor_out[14][21][0];
assign sum_out[3][21][0] = xor_out[15][21][0] + xor_out[16][21][0] + xor_out[17][21][0] + xor_out[18][21][0] + xor_out[19][21][0];
assign sum_out[4][21][0] = xor_out[20][21][0] + xor_out[21][21][0] + xor_out[22][21][0] + xor_out[23][21][0] + xor_out[24][21][0];
assign sum_out[5][21][0] = xor_out[25][21][0] + xor_out[26][21][0] + xor_out[27][21][0] + xor_out[28][21][0] + xor_out[29][21][0];
assign sum_out[6][21][0] = xor_out[30][21][0] + xor_out[31][21][0] + xor_out[32][21][0] + xor_out[33][21][0] + xor_out[34][21][0];
assign sum_out[7][21][0] = xor_out[35][21][0] + xor_out[36][21][0] + xor_out[37][21][0] + xor_out[38][21][0] + xor_out[39][21][0];
assign sum_out[8][21][0] = xor_out[40][21][0] + xor_out[41][21][0] + xor_out[42][21][0] + xor_out[43][21][0] + xor_out[44][21][0];
assign sum_out[9][21][0] = xor_out[45][21][0] + xor_out[46][21][0] + xor_out[47][21][0] + xor_out[48][21][0] + xor_out[49][21][0];
assign sum_out[10][21][0] = xor_out[50][21][0] + xor_out[51][21][0] + xor_out[52][21][0] + xor_out[53][21][0] + xor_out[54][21][0];
assign sum_out[11][21][0] = xor_out[55][21][0] + xor_out[56][21][0] + xor_out[57][21][0] + xor_out[58][21][0] + xor_out[59][21][0];
assign sum_out[12][21][0] = xor_out[60][21][0] + xor_out[61][21][0] + xor_out[62][21][0] + xor_out[63][21][0] + xor_out[64][21][0];
assign sum_out[13][21][0] = xor_out[65][21][0] + xor_out[66][21][0] + xor_out[67][21][0] + xor_out[68][21][0] + xor_out[69][21][0];
assign sum_out[14][21][0] = xor_out[70][21][0] + xor_out[71][21][0] + xor_out[72][21][0] + xor_out[73][21][0] + xor_out[74][21][0];
assign sum_out[15][21][0] = xor_out[75][21][0] + xor_out[76][21][0] + xor_out[77][21][0] + xor_out[78][21][0] + xor_out[79][21][0];
assign sum_out[16][21][0] = xor_out[80][21][0] + xor_out[81][21][0] + xor_out[82][21][0] + xor_out[83][21][0] + xor_out[84][21][0];
assign sum_out[17][21][0] = xor_out[85][21][0] + xor_out[86][21][0] + xor_out[87][21][0] + xor_out[88][21][0] + xor_out[89][21][0];
assign sum_out[18][21][0] = xor_out[90][21][0] + xor_out[91][21][0] + xor_out[92][21][0] + xor_out[93][21][0] + xor_out[94][21][0];
assign sum_out[19][21][0] = xor_out[95][21][0] + xor_out[96][21][0] + xor_out[97][21][0] + xor_out[98][21][0] + xor_out[99][21][0];

assign sum_out[0][21][1] = xor_out[0][21][1] + xor_out[1][21][1] + xor_out[2][21][1] + xor_out[3][21][1] + xor_out[4][21][1];
assign sum_out[1][21][1] = xor_out[5][21][1] + xor_out[6][21][1] + xor_out[7][21][1] + xor_out[8][21][1] + xor_out[9][21][1];
assign sum_out[2][21][1] = xor_out[10][21][1] + xor_out[11][21][1] + xor_out[12][21][1] + xor_out[13][21][1] + xor_out[14][21][1];
assign sum_out[3][21][1] = xor_out[15][21][1] + xor_out[16][21][1] + xor_out[17][21][1] + xor_out[18][21][1] + xor_out[19][21][1];
assign sum_out[4][21][1] = xor_out[20][21][1] + xor_out[21][21][1] + xor_out[22][21][1] + xor_out[23][21][1] + xor_out[24][21][1];
assign sum_out[5][21][1] = xor_out[25][21][1] + xor_out[26][21][1] + xor_out[27][21][1] + xor_out[28][21][1] + xor_out[29][21][1];
assign sum_out[6][21][1] = xor_out[30][21][1] + xor_out[31][21][1] + xor_out[32][21][1] + xor_out[33][21][1] + xor_out[34][21][1];
assign sum_out[7][21][1] = xor_out[35][21][1] + xor_out[36][21][1] + xor_out[37][21][1] + xor_out[38][21][1] + xor_out[39][21][1];
assign sum_out[8][21][1] = xor_out[40][21][1] + xor_out[41][21][1] + xor_out[42][21][1] + xor_out[43][21][1] + xor_out[44][21][1];
assign sum_out[9][21][1] = xor_out[45][21][1] + xor_out[46][21][1] + xor_out[47][21][1] + xor_out[48][21][1] + xor_out[49][21][1];
assign sum_out[10][21][1] = xor_out[50][21][1] + xor_out[51][21][1] + xor_out[52][21][1] + xor_out[53][21][1] + xor_out[54][21][1];
assign sum_out[11][21][1] = xor_out[55][21][1] + xor_out[56][21][1] + xor_out[57][21][1] + xor_out[58][21][1] + xor_out[59][21][1];
assign sum_out[12][21][1] = xor_out[60][21][1] + xor_out[61][21][1] + xor_out[62][21][1] + xor_out[63][21][1] + xor_out[64][21][1];
assign sum_out[13][21][1] = xor_out[65][21][1] + xor_out[66][21][1] + xor_out[67][21][1] + xor_out[68][21][1] + xor_out[69][21][1];
assign sum_out[14][21][1] = xor_out[70][21][1] + xor_out[71][21][1] + xor_out[72][21][1] + xor_out[73][21][1] + xor_out[74][21][1];
assign sum_out[15][21][1] = xor_out[75][21][1] + xor_out[76][21][1] + xor_out[77][21][1] + xor_out[78][21][1] + xor_out[79][21][1];
assign sum_out[16][21][1] = xor_out[80][21][1] + xor_out[81][21][1] + xor_out[82][21][1] + xor_out[83][21][1] + xor_out[84][21][1];
assign sum_out[17][21][1] = xor_out[85][21][1] + xor_out[86][21][1] + xor_out[87][21][1] + xor_out[88][21][1] + xor_out[89][21][1];
assign sum_out[18][21][1] = xor_out[90][21][1] + xor_out[91][21][1] + xor_out[92][21][1] + xor_out[93][21][1] + xor_out[94][21][1];
assign sum_out[19][21][1] = xor_out[95][21][1] + xor_out[96][21][1] + xor_out[97][21][1] + xor_out[98][21][1] + xor_out[99][21][1];

assign sum_out[0][21][2] = xor_out[0][21][2] + xor_out[1][21][2] + xor_out[2][21][2] + xor_out[3][21][2] + xor_out[4][21][2];
assign sum_out[1][21][2] = xor_out[5][21][2] + xor_out[6][21][2] + xor_out[7][21][2] + xor_out[8][21][2] + xor_out[9][21][2];
assign sum_out[2][21][2] = xor_out[10][21][2] + xor_out[11][21][2] + xor_out[12][21][2] + xor_out[13][21][2] + xor_out[14][21][2];
assign sum_out[3][21][2] = xor_out[15][21][2] + xor_out[16][21][2] + xor_out[17][21][2] + xor_out[18][21][2] + xor_out[19][21][2];
assign sum_out[4][21][2] = xor_out[20][21][2] + xor_out[21][21][2] + xor_out[22][21][2] + xor_out[23][21][2] + xor_out[24][21][2];
assign sum_out[5][21][2] = xor_out[25][21][2] + xor_out[26][21][2] + xor_out[27][21][2] + xor_out[28][21][2] + xor_out[29][21][2];
assign sum_out[6][21][2] = xor_out[30][21][2] + xor_out[31][21][2] + xor_out[32][21][2] + xor_out[33][21][2] + xor_out[34][21][2];
assign sum_out[7][21][2] = xor_out[35][21][2] + xor_out[36][21][2] + xor_out[37][21][2] + xor_out[38][21][2] + xor_out[39][21][2];
assign sum_out[8][21][2] = xor_out[40][21][2] + xor_out[41][21][2] + xor_out[42][21][2] + xor_out[43][21][2] + xor_out[44][21][2];
assign sum_out[9][21][2] = xor_out[45][21][2] + xor_out[46][21][2] + xor_out[47][21][2] + xor_out[48][21][2] + xor_out[49][21][2];
assign sum_out[10][21][2] = xor_out[50][21][2] + xor_out[51][21][2] + xor_out[52][21][2] + xor_out[53][21][2] + xor_out[54][21][2];
assign sum_out[11][21][2] = xor_out[55][21][2] + xor_out[56][21][2] + xor_out[57][21][2] + xor_out[58][21][2] + xor_out[59][21][2];
assign sum_out[12][21][2] = xor_out[60][21][2] + xor_out[61][21][2] + xor_out[62][21][2] + xor_out[63][21][2] + xor_out[64][21][2];
assign sum_out[13][21][2] = xor_out[65][21][2] + xor_out[66][21][2] + xor_out[67][21][2] + xor_out[68][21][2] + xor_out[69][21][2];
assign sum_out[14][21][2] = xor_out[70][21][2] + xor_out[71][21][2] + xor_out[72][21][2] + xor_out[73][21][2] + xor_out[74][21][2];
assign sum_out[15][21][2] = xor_out[75][21][2] + xor_out[76][21][2] + xor_out[77][21][2] + xor_out[78][21][2] + xor_out[79][21][2];
assign sum_out[16][21][2] = xor_out[80][21][2] + xor_out[81][21][2] + xor_out[82][21][2] + xor_out[83][21][2] + xor_out[84][21][2];
assign sum_out[17][21][2] = xor_out[85][21][2] + xor_out[86][21][2] + xor_out[87][21][2] + xor_out[88][21][2] + xor_out[89][21][2];
assign sum_out[18][21][2] = xor_out[90][21][2] + xor_out[91][21][2] + xor_out[92][21][2] + xor_out[93][21][2] + xor_out[94][21][2];
assign sum_out[19][21][2] = xor_out[95][21][2] + xor_out[96][21][2] + xor_out[97][21][2] + xor_out[98][21][2] + xor_out[99][21][2];

assign sum_out[0][21][3] = xor_out[0][21][3] + xor_out[1][21][3] + xor_out[2][21][3] + xor_out[3][21][3] + xor_out[4][21][3];
assign sum_out[1][21][3] = xor_out[5][21][3] + xor_out[6][21][3] + xor_out[7][21][3] + xor_out[8][21][3] + xor_out[9][21][3];
assign sum_out[2][21][3] = xor_out[10][21][3] + xor_out[11][21][3] + xor_out[12][21][3] + xor_out[13][21][3] + xor_out[14][21][3];
assign sum_out[3][21][3] = xor_out[15][21][3] + xor_out[16][21][3] + xor_out[17][21][3] + xor_out[18][21][3] + xor_out[19][21][3];
assign sum_out[4][21][3] = xor_out[20][21][3] + xor_out[21][21][3] + xor_out[22][21][3] + xor_out[23][21][3] + xor_out[24][21][3];
assign sum_out[5][21][3] = xor_out[25][21][3] + xor_out[26][21][3] + xor_out[27][21][3] + xor_out[28][21][3] + xor_out[29][21][3];
assign sum_out[6][21][3] = xor_out[30][21][3] + xor_out[31][21][3] + xor_out[32][21][3] + xor_out[33][21][3] + xor_out[34][21][3];
assign sum_out[7][21][3] = xor_out[35][21][3] + xor_out[36][21][3] + xor_out[37][21][3] + xor_out[38][21][3] + xor_out[39][21][3];
assign sum_out[8][21][3] = xor_out[40][21][3] + xor_out[41][21][3] + xor_out[42][21][3] + xor_out[43][21][3] + xor_out[44][21][3];
assign sum_out[9][21][3] = xor_out[45][21][3] + xor_out[46][21][3] + xor_out[47][21][3] + xor_out[48][21][3] + xor_out[49][21][3];
assign sum_out[10][21][3] = xor_out[50][21][3] + xor_out[51][21][3] + xor_out[52][21][3] + xor_out[53][21][3] + xor_out[54][21][3];
assign sum_out[11][21][3] = xor_out[55][21][3] + xor_out[56][21][3] + xor_out[57][21][3] + xor_out[58][21][3] + xor_out[59][21][3];
assign sum_out[12][21][3] = xor_out[60][21][3] + xor_out[61][21][3] + xor_out[62][21][3] + xor_out[63][21][3] + xor_out[64][21][3];
assign sum_out[13][21][3] = xor_out[65][21][3] + xor_out[66][21][3] + xor_out[67][21][3] + xor_out[68][21][3] + xor_out[69][21][3];
assign sum_out[14][21][3] = xor_out[70][21][3] + xor_out[71][21][3] + xor_out[72][21][3] + xor_out[73][21][3] + xor_out[74][21][3];
assign sum_out[15][21][3] = xor_out[75][21][3] + xor_out[76][21][3] + xor_out[77][21][3] + xor_out[78][21][3] + xor_out[79][21][3];
assign sum_out[16][21][3] = xor_out[80][21][3] + xor_out[81][21][3] + xor_out[82][21][3] + xor_out[83][21][3] + xor_out[84][21][3];
assign sum_out[17][21][3] = xor_out[85][21][3] + xor_out[86][21][3] + xor_out[87][21][3] + xor_out[88][21][3] + xor_out[89][21][3];
assign sum_out[18][21][3] = xor_out[90][21][3] + xor_out[91][21][3] + xor_out[92][21][3] + xor_out[93][21][3] + xor_out[94][21][3];
assign sum_out[19][21][3] = xor_out[95][21][3] + xor_out[96][21][3] + xor_out[97][21][3] + xor_out[98][21][3] + xor_out[99][21][3];

assign sum_out[0][21][4] = xor_out[0][21][4] + xor_out[1][21][4] + xor_out[2][21][4] + xor_out[3][21][4] + xor_out[4][21][4];
assign sum_out[1][21][4] = xor_out[5][21][4] + xor_out[6][21][4] + xor_out[7][21][4] + xor_out[8][21][4] + xor_out[9][21][4];
assign sum_out[2][21][4] = xor_out[10][21][4] + xor_out[11][21][4] + xor_out[12][21][4] + xor_out[13][21][4] + xor_out[14][21][4];
assign sum_out[3][21][4] = xor_out[15][21][4] + xor_out[16][21][4] + xor_out[17][21][4] + xor_out[18][21][4] + xor_out[19][21][4];
assign sum_out[4][21][4] = xor_out[20][21][4] + xor_out[21][21][4] + xor_out[22][21][4] + xor_out[23][21][4] + xor_out[24][21][4];
assign sum_out[5][21][4] = xor_out[25][21][4] + xor_out[26][21][4] + xor_out[27][21][4] + xor_out[28][21][4] + xor_out[29][21][4];
assign sum_out[6][21][4] = xor_out[30][21][4] + xor_out[31][21][4] + xor_out[32][21][4] + xor_out[33][21][4] + xor_out[34][21][4];
assign sum_out[7][21][4] = xor_out[35][21][4] + xor_out[36][21][4] + xor_out[37][21][4] + xor_out[38][21][4] + xor_out[39][21][4];
assign sum_out[8][21][4] = xor_out[40][21][4] + xor_out[41][21][4] + xor_out[42][21][4] + xor_out[43][21][4] + xor_out[44][21][4];
assign sum_out[9][21][4] = xor_out[45][21][4] + xor_out[46][21][4] + xor_out[47][21][4] + xor_out[48][21][4] + xor_out[49][21][4];
assign sum_out[10][21][4] = xor_out[50][21][4] + xor_out[51][21][4] + xor_out[52][21][4] + xor_out[53][21][4] + xor_out[54][21][4];
assign sum_out[11][21][4] = xor_out[55][21][4] + xor_out[56][21][4] + xor_out[57][21][4] + xor_out[58][21][4] + xor_out[59][21][4];
assign sum_out[12][21][4] = xor_out[60][21][4] + xor_out[61][21][4] + xor_out[62][21][4] + xor_out[63][21][4] + xor_out[64][21][4];
assign sum_out[13][21][4] = xor_out[65][21][4] + xor_out[66][21][4] + xor_out[67][21][4] + xor_out[68][21][4] + xor_out[69][21][4];
assign sum_out[14][21][4] = xor_out[70][21][4] + xor_out[71][21][4] + xor_out[72][21][4] + xor_out[73][21][4] + xor_out[74][21][4];
assign sum_out[15][21][4] = xor_out[75][21][4] + xor_out[76][21][4] + xor_out[77][21][4] + xor_out[78][21][4] + xor_out[79][21][4];
assign sum_out[16][21][4] = xor_out[80][21][4] + xor_out[81][21][4] + xor_out[82][21][4] + xor_out[83][21][4] + xor_out[84][21][4];
assign sum_out[17][21][4] = xor_out[85][21][4] + xor_out[86][21][4] + xor_out[87][21][4] + xor_out[88][21][4] + xor_out[89][21][4];
assign sum_out[18][21][4] = xor_out[90][21][4] + xor_out[91][21][4] + xor_out[92][21][4] + xor_out[93][21][4] + xor_out[94][21][4];
assign sum_out[19][21][4] = xor_out[95][21][4] + xor_out[96][21][4] + xor_out[97][21][4] + xor_out[98][21][4] + xor_out[99][21][4];

assign sum_out[0][21][5] = xor_out[0][21][5] + xor_out[1][21][5] + xor_out[2][21][5] + xor_out[3][21][5] + xor_out[4][21][5];
assign sum_out[1][21][5] = xor_out[5][21][5] + xor_out[6][21][5] + xor_out[7][21][5] + xor_out[8][21][5] + xor_out[9][21][5];
assign sum_out[2][21][5] = xor_out[10][21][5] + xor_out[11][21][5] + xor_out[12][21][5] + xor_out[13][21][5] + xor_out[14][21][5];
assign sum_out[3][21][5] = xor_out[15][21][5] + xor_out[16][21][5] + xor_out[17][21][5] + xor_out[18][21][5] + xor_out[19][21][5];
assign sum_out[4][21][5] = xor_out[20][21][5] + xor_out[21][21][5] + xor_out[22][21][5] + xor_out[23][21][5] + xor_out[24][21][5];
assign sum_out[5][21][5] = xor_out[25][21][5] + xor_out[26][21][5] + xor_out[27][21][5] + xor_out[28][21][5] + xor_out[29][21][5];
assign sum_out[6][21][5] = xor_out[30][21][5] + xor_out[31][21][5] + xor_out[32][21][5] + xor_out[33][21][5] + xor_out[34][21][5];
assign sum_out[7][21][5] = xor_out[35][21][5] + xor_out[36][21][5] + xor_out[37][21][5] + xor_out[38][21][5] + xor_out[39][21][5];
assign sum_out[8][21][5] = xor_out[40][21][5] + xor_out[41][21][5] + xor_out[42][21][5] + xor_out[43][21][5] + xor_out[44][21][5];
assign sum_out[9][21][5] = xor_out[45][21][5] + xor_out[46][21][5] + xor_out[47][21][5] + xor_out[48][21][5] + xor_out[49][21][5];
assign sum_out[10][21][5] = xor_out[50][21][5] + xor_out[51][21][5] + xor_out[52][21][5] + xor_out[53][21][5] + xor_out[54][21][5];
assign sum_out[11][21][5] = xor_out[55][21][5] + xor_out[56][21][5] + xor_out[57][21][5] + xor_out[58][21][5] + xor_out[59][21][5];
assign sum_out[12][21][5] = xor_out[60][21][5] + xor_out[61][21][5] + xor_out[62][21][5] + xor_out[63][21][5] + xor_out[64][21][5];
assign sum_out[13][21][5] = xor_out[65][21][5] + xor_out[66][21][5] + xor_out[67][21][5] + xor_out[68][21][5] + xor_out[69][21][5];
assign sum_out[14][21][5] = xor_out[70][21][5] + xor_out[71][21][5] + xor_out[72][21][5] + xor_out[73][21][5] + xor_out[74][21][5];
assign sum_out[15][21][5] = xor_out[75][21][5] + xor_out[76][21][5] + xor_out[77][21][5] + xor_out[78][21][5] + xor_out[79][21][5];
assign sum_out[16][21][5] = xor_out[80][21][5] + xor_out[81][21][5] + xor_out[82][21][5] + xor_out[83][21][5] + xor_out[84][21][5];
assign sum_out[17][21][5] = xor_out[85][21][5] + xor_out[86][21][5] + xor_out[87][21][5] + xor_out[88][21][5] + xor_out[89][21][5];
assign sum_out[18][21][5] = xor_out[90][21][5] + xor_out[91][21][5] + xor_out[92][21][5] + xor_out[93][21][5] + xor_out[94][21][5];
assign sum_out[19][21][5] = xor_out[95][21][5] + xor_out[96][21][5] + xor_out[97][21][5] + xor_out[98][21][5] + xor_out[99][21][5];

assign sum_out[0][21][6] = xor_out[0][21][6] + xor_out[1][21][6] + xor_out[2][21][6] + xor_out[3][21][6] + xor_out[4][21][6];
assign sum_out[1][21][6] = xor_out[5][21][6] + xor_out[6][21][6] + xor_out[7][21][6] + xor_out[8][21][6] + xor_out[9][21][6];
assign sum_out[2][21][6] = xor_out[10][21][6] + xor_out[11][21][6] + xor_out[12][21][6] + xor_out[13][21][6] + xor_out[14][21][6];
assign sum_out[3][21][6] = xor_out[15][21][6] + xor_out[16][21][6] + xor_out[17][21][6] + xor_out[18][21][6] + xor_out[19][21][6];
assign sum_out[4][21][6] = xor_out[20][21][6] + xor_out[21][21][6] + xor_out[22][21][6] + xor_out[23][21][6] + xor_out[24][21][6];
assign sum_out[5][21][6] = xor_out[25][21][6] + xor_out[26][21][6] + xor_out[27][21][6] + xor_out[28][21][6] + xor_out[29][21][6];
assign sum_out[6][21][6] = xor_out[30][21][6] + xor_out[31][21][6] + xor_out[32][21][6] + xor_out[33][21][6] + xor_out[34][21][6];
assign sum_out[7][21][6] = xor_out[35][21][6] + xor_out[36][21][6] + xor_out[37][21][6] + xor_out[38][21][6] + xor_out[39][21][6];
assign sum_out[8][21][6] = xor_out[40][21][6] + xor_out[41][21][6] + xor_out[42][21][6] + xor_out[43][21][6] + xor_out[44][21][6];
assign sum_out[9][21][6] = xor_out[45][21][6] + xor_out[46][21][6] + xor_out[47][21][6] + xor_out[48][21][6] + xor_out[49][21][6];
assign sum_out[10][21][6] = xor_out[50][21][6] + xor_out[51][21][6] + xor_out[52][21][6] + xor_out[53][21][6] + xor_out[54][21][6];
assign sum_out[11][21][6] = xor_out[55][21][6] + xor_out[56][21][6] + xor_out[57][21][6] + xor_out[58][21][6] + xor_out[59][21][6];
assign sum_out[12][21][6] = xor_out[60][21][6] + xor_out[61][21][6] + xor_out[62][21][6] + xor_out[63][21][6] + xor_out[64][21][6];
assign sum_out[13][21][6] = xor_out[65][21][6] + xor_out[66][21][6] + xor_out[67][21][6] + xor_out[68][21][6] + xor_out[69][21][6];
assign sum_out[14][21][6] = xor_out[70][21][6] + xor_out[71][21][6] + xor_out[72][21][6] + xor_out[73][21][6] + xor_out[74][21][6];
assign sum_out[15][21][6] = xor_out[75][21][6] + xor_out[76][21][6] + xor_out[77][21][6] + xor_out[78][21][6] + xor_out[79][21][6];
assign sum_out[16][21][6] = xor_out[80][21][6] + xor_out[81][21][6] + xor_out[82][21][6] + xor_out[83][21][6] + xor_out[84][21][6];
assign sum_out[17][21][6] = xor_out[85][21][6] + xor_out[86][21][6] + xor_out[87][21][6] + xor_out[88][21][6] + xor_out[89][21][6];
assign sum_out[18][21][6] = xor_out[90][21][6] + xor_out[91][21][6] + xor_out[92][21][6] + xor_out[93][21][6] + xor_out[94][21][6];
assign sum_out[19][21][6] = xor_out[95][21][6] + xor_out[96][21][6] + xor_out[97][21][6] + xor_out[98][21][6] + xor_out[99][21][6];

assign sum_out[0][21][7] = xor_out[0][21][7] + xor_out[1][21][7] + xor_out[2][21][7] + xor_out[3][21][7] + xor_out[4][21][7];
assign sum_out[1][21][7] = xor_out[5][21][7] + xor_out[6][21][7] + xor_out[7][21][7] + xor_out[8][21][7] + xor_out[9][21][7];
assign sum_out[2][21][7] = xor_out[10][21][7] + xor_out[11][21][7] + xor_out[12][21][7] + xor_out[13][21][7] + xor_out[14][21][7];
assign sum_out[3][21][7] = xor_out[15][21][7] + xor_out[16][21][7] + xor_out[17][21][7] + xor_out[18][21][7] + xor_out[19][21][7];
assign sum_out[4][21][7] = xor_out[20][21][7] + xor_out[21][21][7] + xor_out[22][21][7] + xor_out[23][21][7] + xor_out[24][21][7];
assign sum_out[5][21][7] = xor_out[25][21][7] + xor_out[26][21][7] + xor_out[27][21][7] + xor_out[28][21][7] + xor_out[29][21][7];
assign sum_out[6][21][7] = xor_out[30][21][7] + xor_out[31][21][7] + xor_out[32][21][7] + xor_out[33][21][7] + xor_out[34][21][7];
assign sum_out[7][21][7] = xor_out[35][21][7] + xor_out[36][21][7] + xor_out[37][21][7] + xor_out[38][21][7] + xor_out[39][21][7];
assign sum_out[8][21][7] = xor_out[40][21][7] + xor_out[41][21][7] + xor_out[42][21][7] + xor_out[43][21][7] + xor_out[44][21][7];
assign sum_out[9][21][7] = xor_out[45][21][7] + xor_out[46][21][7] + xor_out[47][21][7] + xor_out[48][21][7] + xor_out[49][21][7];
assign sum_out[10][21][7] = xor_out[50][21][7] + xor_out[51][21][7] + xor_out[52][21][7] + xor_out[53][21][7] + xor_out[54][21][7];
assign sum_out[11][21][7] = xor_out[55][21][7] + xor_out[56][21][7] + xor_out[57][21][7] + xor_out[58][21][7] + xor_out[59][21][7];
assign sum_out[12][21][7] = xor_out[60][21][7] + xor_out[61][21][7] + xor_out[62][21][7] + xor_out[63][21][7] + xor_out[64][21][7];
assign sum_out[13][21][7] = xor_out[65][21][7] + xor_out[66][21][7] + xor_out[67][21][7] + xor_out[68][21][7] + xor_out[69][21][7];
assign sum_out[14][21][7] = xor_out[70][21][7] + xor_out[71][21][7] + xor_out[72][21][7] + xor_out[73][21][7] + xor_out[74][21][7];
assign sum_out[15][21][7] = xor_out[75][21][7] + xor_out[76][21][7] + xor_out[77][21][7] + xor_out[78][21][7] + xor_out[79][21][7];
assign sum_out[16][21][7] = xor_out[80][21][7] + xor_out[81][21][7] + xor_out[82][21][7] + xor_out[83][21][7] + xor_out[84][21][7];
assign sum_out[17][21][7] = xor_out[85][21][7] + xor_out[86][21][7] + xor_out[87][21][7] + xor_out[88][21][7] + xor_out[89][21][7];
assign sum_out[18][21][7] = xor_out[90][21][7] + xor_out[91][21][7] + xor_out[92][21][7] + xor_out[93][21][7] + xor_out[94][21][7];
assign sum_out[19][21][7] = xor_out[95][21][7] + xor_out[96][21][7] + xor_out[97][21][7] + xor_out[98][21][7] + xor_out[99][21][7];

assign sum_out[0][21][8] = xor_out[0][21][8] + xor_out[1][21][8] + xor_out[2][21][8] + xor_out[3][21][8] + xor_out[4][21][8];
assign sum_out[1][21][8] = xor_out[5][21][8] + xor_out[6][21][8] + xor_out[7][21][8] + xor_out[8][21][8] + xor_out[9][21][8];
assign sum_out[2][21][8] = xor_out[10][21][8] + xor_out[11][21][8] + xor_out[12][21][8] + xor_out[13][21][8] + xor_out[14][21][8];
assign sum_out[3][21][8] = xor_out[15][21][8] + xor_out[16][21][8] + xor_out[17][21][8] + xor_out[18][21][8] + xor_out[19][21][8];
assign sum_out[4][21][8] = xor_out[20][21][8] + xor_out[21][21][8] + xor_out[22][21][8] + xor_out[23][21][8] + xor_out[24][21][8];
assign sum_out[5][21][8] = xor_out[25][21][8] + xor_out[26][21][8] + xor_out[27][21][8] + xor_out[28][21][8] + xor_out[29][21][8];
assign sum_out[6][21][8] = xor_out[30][21][8] + xor_out[31][21][8] + xor_out[32][21][8] + xor_out[33][21][8] + xor_out[34][21][8];
assign sum_out[7][21][8] = xor_out[35][21][8] + xor_out[36][21][8] + xor_out[37][21][8] + xor_out[38][21][8] + xor_out[39][21][8];
assign sum_out[8][21][8] = xor_out[40][21][8] + xor_out[41][21][8] + xor_out[42][21][8] + xor_out[43][21][8] + xor_out[44][21][8];
assign sum_out[9][21][8] = xor_out[45][21][8] + xor_out[46][21][8] + xor_out[47][21][8] + xor_out[48][21][8] + xor_out[49][21][8];
assign sum_out[10][21][8] = xor_out[50][21][8] + xor_out[51][21][8] + xor_out[52][21][8] + xor_out[53][21][8] + xor_out[54][21][8];
assign sum_out[11][21][8] = xor_out[55][21][8] + xor_out[56][21][8] + xor_out[57][21][8] + xor_out[58][21][8] + xor_out[59][21][8];
assign sum_out[12][21][8] = xor_out[60][21][8] + xor_out[61][21][8] + xor_out[62][21][8] + xor_out[63][21][8] + xor_out[64][21][8];
assign sum_out[13][21][8] = xor_out[65][21][8] + xor_out[66][21][8] + xor_out[67][21][8] + xor_out[68][21][8] + xor_out[69][21][8];
assign sum_out[14][21][8] = xor_out[70][21][8] + xor_out[71][21][8] + xor_out[72][21][8] + xor_out[73][21][8] + xor_out[74][21][8];
assign sum_out[15][21][8] = xor_out[75][21][8] + xor_out[76][21][8] + xor_out[77][21][8] + xor_out[78][21][8] + xor_out[79][21][8];
assign sum_out[16][21][8] = xor_out[80][21][8] + xor_out[81][21][8] + xor_out[82][21][8] + xor_out[83][21][8] + xor_out[84][21][8];
assign sum_out[17][21][8] = xor_out[85][21][8] + xor_out[86][21][8] + xor_out[87][21][8] + xor_out[88][21][8] + xor_out[89][21][8];
assign sum_out[18][21][8] = xor_out[90][21][8] + xor_out[91][21][8] + xor_out[92][21][8] + xor_out[93][21][8] + xor_out[94][21][8];
assign sum_out[19][21][8] = xor_out[95][21][8] + xor_out[96][21][8] + xor_out[97][21][8] + xor_out[98][21][8] + xor_out[99][21][8];

assign sum_out[0][21][9] = xor_out[0][21][9] + xor_out[1][21][9] + xor_out[2][21][9] + xor_out[3][21][9] + xor_out[4][21][9];
assign sum_out[1][21][9] = xor_out[5][21][9] + xor_out[6][21][9] + xor_out[7][21][9] + xor_out[8][21][9] + xor_out[9][21][9];
assign sum_out[2][21][9] = xor_out[10][21][9] + xor_out[11][21][9] + xor_out[12][21][9] + xor_out[13][21][9] + xor_out[14][21][9];
assign sum_out[3][21][9] = xor_out[15][21][9] + xor_out[16][21][9] + xor_out[17][21][9] + xor_out[18][21][9] + xor_out[19][21][9];
assign sum_out[4][21][9] = xor_out[20][21][9] + xor_out[21][21][9] + xor_out[22][21][9] + xor_out[23][21][9] + xor_out[24][21][9];
assign sum_out[5][21][9] = xor_out[25][21][9] + xor_out[26][21][9] + xor_out[27][21][9] + xor_out[28][21][9] + xor_out[29][21][9];
assign sum_out[6][21][9] = xor_out[30][21][9] + xor_out[31][21][9] + xor_out[32][21][9] + xor_out[33][21][9] + xor_out[34][21][9];
assign sum_out[7][21][9] = xor_out[35][21][9] + xor_out[36][21][9] + xor_out[37][21][9] + xor_out[38][21][9] + xor_out[39][21][9];
assign sum_out[8][21][9] = xor_out[40][21][9] + xor_out[41][21][9] + xor_out[42][21][9] + xor_out[43][21][9] + xor_out[44][21][9];
assign sum_out[9][21][9] = xor_out[45][21][9] + xor_out[46][21][9] + xor_out[47][21][9] + xor_out[48][21][9] + xor_out[49][21][9];
assign sum_out[10][21][9] = xor_out[50][21][9] + xor_out[51][21][9] + xor_out[52][21][9] + xor_out[53][21][9] + xor_out[54][21][9];
assign sum_out[11][21][9] = xor_out[55][21][9] + xor_out[56][21][9] + xor_out[57][21][9] + xor_out[58][21][9] + xor_out[59][21][9];
assign sum_out[12][21][9] = xor_out[60][21][9] + xor_out[61][21][9] + xor_out[62][21][9] + xor_out[63][21][9] + xor_out[64][21][9];
assign sum_out[13][21][9] = xor_out[65][21][9] + xor_out[66][21][9] + xor_out[67][21][9] + xor_out[68][21][9] + xor_out[69][21][9];
assign sum_out[14][21][9] = xor_out[70][21][9] + xor_out[71][21][9] + xor_out[72][21][9] + xor_out[73][21][9] + xor_out[74][21][9];
assign sum_out[15][21][9] = xor_out[75][21][9] + xor_out[76][21][9] + xor_out[77][21][9] + xor_out[78][21][9] + xor_out[79][21][9];
assign sum_out[16][21][9] = xor_out[80][21][9] + xor_out[81][21][9] + xor_out[82][21][9] + xor_out[83][21][9] + xor_out[84][21][9];
assign sum_out[17][21][9] = xor_out[85][21][9] + xor_out[86][21][9] + xor_out[87][21][9] + xor_out[88][21][9] + xor_out[89][21][9];
assign sum_out[18][21][9] = xor_out[90][21][9] + xor_out[91][21][9] + xor_out[92][21][9] + xor_out[93][21][9] + xor_out[94][21][9];
assign sum_out[19][21][9] = xor_out[95][21][9] + xor_out[96][21][9] + xor_out[97][21][9] + xor_out[98][21][9] + xor_out[99][21][9];

assign sum_out[0][21][10] = xor_out[0][21][10] + xor_out[1][21][10] + xor_out[2][21][10] + xor_out[3][21][10] + xor_out[4][21][10];
assign sum_out[1][21][10] = xor_out[5][21][10] + xor_out[6][21][10] + xor_out[7][21][10] + xor_out[8][21][10] + xor_out[9][21][10];
assign sum_out[2][21][10] = xor_out[10][21][10] + xor_out[11][21][10] + xor_out[12][21][10] + xor_out[13][21][10] + xor_out[14][21][10];
assign sum_out[3][21][10] = xor_out[15][21][10] + xor_out[16][21][10] + xor_out[17][21][10] + xor_out[18][21][10] + xor_out[19][21][10];
assign sum_out[4][21][10] = xor_out[20][21][10] + xor_out[21][21][10] + xor_out[22][21][10] + xor_out[23][21][10] + xor_out[24][21][10];
assign sum_out[5][21][10] = xor_out[25][21][10] + xor_out[26][21][10] + xor_out[27][21][10] + xor_out[28][21][10] + xor_out[29][21][10];
assign sum_out[6][21][10] = xor_out[30][21][10] + xor_out[31][21][10] + xor_out[32][21][10] + xor_out[33][21][10] + xor_out[34][21][10];
assign sum_out[7][21][10] = xor_out[35][21][10] + xor_out[36][21][10] + xor_out[37][21][10] + xor_out[38][21][10] + xor_out[39][21][10];
assign sum_out[8][21][10] = xor_out[40][21][10] + xor_out[41][21][10] + xor_out[42][21][10] + xor_out[43][21][10] + xor_out[44][21][10];
assign sum_out[9][21][10] = xor_out[45][21][10] + xor_out[46][21][10] + xor_out[47][21][10] + xor_out[48][21][10] + xor_out[49][21][10];
assign sum_out[10][21][10] = xor_out[50][21][10] + xor_out[51][21][10] + xor_out[52][21][10] + xor_out[53][21][10] + xor_out[54][21][10];
assign sum_out[11][21][10] = xor_out[55][21][10] + xor_out[56][21][10] + xor_out[57][21][10] + xor_out[58][21][10] + xor_out[59][21][10];
assign sum_out[12][21][10] = xor_out[60][21][10] + xor_out[61][21][10] + xor_out[62][21][10] + xor_out[63][21][10] + xor_out[64][21][10];
assign sum_out[13][21][10] = xor_out[65][21][10] + xor_out[66][21][10] + xor_out[67][21][10] + xor_out[68][21][10] + xor_out[69][21][10];
assign sum_out[14][21][10] = xor_out[70][21][10] + xor_out[71][21][10] + xor_out[72][21][10] + xor_out[73][21][10] + xor_out[74][21][10];
assign sum_out[15][21][10] = xor_out[75][21][10] + xor_out[76][21][10] + xor_out[77][21][10] + xor_out[78][21][10] + xor_out[79][21][10];
assign sum_out[16][21][10] = xor_out[80][21][10] + xor_out[81][21][10] + xor_out[82][21][10] + xor_out[83][21][10] + xor_out[84][21][10];
assign sum_out[17][21][10] = xor_out[85][21][10] + xor_out[86][21][10] + xor_out[87][21][10] + xor_out[88][21][10] + xor_out[89][21][10];
assign sum_out[18][21][10] = xor_out[90][21][10] + xor_out[91][21][10] + xor_out[92][21][10] + xor_out[93][21][10] + xor_out[94][21][10];
assign sum_out[19][21][10] = xor_out[95][21][10] + xor_out[96][21][10] + xor_out[97][21][10] + xor_out[98][21][10] + xor_out[99][21][10];

assign sum_out[0][21][11] = xor_out[0][21][11] + xor_out[1][21][11] + xor_out[2][21][11] + xor_out[3][21][11] + xor_out[4][21][11];
assign sum_out[1][21][11] = xor_out[5][21][11] + xor_out[6][21][11] + xor_out[7][21][11] + xor_out[8][21][11] + xor_out[9][21][11];
assign sum_out[2][21][11] = xor_out[10][21][11] + xor_out[11][21][11] + xor_out[12][21][11] + xor_out[13][21][11] + xor_out[14][21][11];
assign sum_out[3][21][11] = xor_out[15][21][11] + xor_out[16][21][11] + xor_out[17][21][11] + xor_out[18][21][11] + xor_out[19][21][11];
assign sum_out[4][21][11] = xor_out[20][21][11] + xor_out[21][21][11] + xor_out[22][21][11] + xor_out[23][21][11] + xor_out[24][21][11];
assign sum_out[5][21][11] = xor_out[25][21][11] + xor_out[26][21][11] + xor_out[27][21][11] + xor_out[28][21][11] + xor_out[29][21][11];
assign sum_out[6][21][11] = xor_out[30][21][11] + xor_out[31][21][11] + xor_out[32][21][11] + xor_out[33][21][11] + xor_out[34][21][11];
assign sum_out[7][21][11] = xor_out[35][21][11] + xor_out[36][21][11] + xor_out[37][21][11] + xor_out[38][21][11] + xor_out[39][21][11];
assign sum_out[8][21][11] = xor_out[40][21][11] + xor_out[41][21][11] + xor_out[42][21][11] + xor_out[43][21][11] + xor_out[44][21][11];
assign sum_out[9][21][11] = xor_out[45][21][11] + xor_out[46][21][11] + xor_out[47][21][11] + xor_out[48][21][11] + xor_out[49][21][11];
assign sum_out[10][21][11] = xor_out[50][21][11] + xor_out[51][21][11] + xor_out[52][21][11] + xor_out[53][21][11] + xor_out[54][21][11];
assign sum_out[11][21][11] = xor_out[55][21][11] + xor_out[56][21][11] + xor_out[57][21][11] + xor_out[58][21][11] + xor_out[59][21][11];
assign sum_out[12][21][11] = xor_out[60][21][11] + xor_out[61][21][11] + xor_out[62][21][11] + xor_out[63][21][11] + xor_out[64][21][11];
assign sum_out[13][21][11] = xor_out[65][21][11] + xor_out[66][21][11] + xor_out[67][21][11] + xor_out[68][21][11] + xor_out[69][21][11];
assign sum_out[14][21][11] = xor_out[70][21][11] + xor_out[71][21][11] + xor_out[72][21][11] + xor_out[73][21][11] + xor_out[74][21][11];
assign sum_out[15][21][11] = xor_out[75][21][11] + xor_out[76][21][11] + xor_out[77][21][11] + xor_out[78][21][11] + xor_out[79][21][11];
assign sum_out[16][21][11] = xor_out[80][21][11] + xor_out[81][21][11] + xor_out[82][21][11] + xor_out[83][21][11] + xor_out[84][21][11];
assign sum_out[17][21][11] = xor_out[85][21][11] + xor_out[86][21][11] + xor_out[87][21][11] + xor_out[88][21][11] + xor_out[89][21][11];
assign sum_out[18][21][11] = xor_out[90][21][11] + xor_out[91][21][11] + xor_out[92][21][11] + xor_out[93][21][11] + xor_out[94][21][11];
assign sum_out[19][21][11] = xor_out[95][21][11] + xor_out[96][21][11] + xor_out[97][21][11] + xor_out[98][21][11] + xor_out[99][21][11];

assign sum_out[0][21][12] = xor_out[0][21][12] + xor_out[1][21][12] + xor_out[2][21][12] + xor_out[3][21][12] + xor_out[4][21][12];
assign sum_out[1][21][12] = xor_out[5][21][12] + xor_out[6][21][12] + xor_out[7][21][12] + xor_out[8][21][12] + xor_out[9][21][12];
assign sum_out[2][21][12] = xor_out[10][21][12] + xor_out[11][21][12] + xor_out[12][21][12] + xor_out[13][21][12] + xor_out[14][21][12];
assign sum_out[3][21][12] = xor_out[15][21][12] + xor_out[16][21][12] + xor_out[17][21][12] + xor_out[18][21][12] + xor_out[19][21][12];
assign sum_out[4][21][12] = xor_out[20][21][12] + xor_out[21][21][12] + xor_out[22][21][12] + xor_out[23][21][12] + xor_out[24][21][12];
assign sum_out[5][21][12] = xor_out[25][21][12] + xor_out[26][21][12] + xor_out[27][21][12] + xor_out[28][21][12] + xor_out[29][21][12];
assign sum_out[6][21][12] = xor_out[30][21][12] + xor_out[31][21][12] + xor_out[32][21][12] + xor_out[33][21][12] + xor_out[34][21][12];
assign sum_out[7][21][12] = xor_out[35][21][12] + xor_out[36][21][12] + xor_out[37][21][12] + xor_out[38][21][12] + xor_out[39][21][12];
assign sum_out[8][21][12] = xor_out[40][21][12] + xor_out[41][21][12] + xor_out[42][21][12] + xor_out[43][21][12] + xor_out[44][21][12];
assign sum_out[9][21][12] = xor_out[45][21][12] + xor_out[46][21][12] + xor_out[47][21][12] + xor_out[48][21][12] + xor_out[49][21][12];
assign sum_out[10][21][12] = xor_out[50][21][12] + xor_out[51][21][12] + xor_out[52][21][12] + xor_out[53][21][12] + xor_out[54][21][12];
assign sum_out[11][21][12] = xor_out[55][21][12] + xor_out[56][21][12] + xor_out[57][21][12] + xor_out[58][21][12] + xor_out[59][21][12];
assign sum_out[12][21][12] = xor_out[60][21][12] + xor_out[61][21][12] + xor_out[62][21][12] + xor_out[63][21][12] + xor_out[64][21][12];
assign sum_out[13][21][12] = xor_out[65][21][12] + xor_out[66][21][12] + xor_out[67][21][12] + xor_out[68][21][12] + xor_out[69][21][12];
assign sum_out[14][21][12] = xor_out[70][21][12] + xor_out[71][21][12] + xor_out[72][21][12] + xor_out[73][21][12] + xor_out[74][21][12];
assign sum_out[15][21][12] = xor_out[75][21][12] + xor_out[76][21][12] + xor_out[77][21][12] + xor_out[78][21][12] + xor_out[79][21][12];
assign sum_out[16][21][12] = xor_out[80][21][12] + xor_out[81][21][12] + xor_out[82][21][12] + xor_out[83][21][12] + xor_out[84][21][12];
assign sum_out[17][21][12] = xor_out[85][21][12] + xor_out[86][21][12] + xor_out[87][21][12] + xor_out[88][21][12] + xor_out[89][21][12];
assign sum_out[18][21][12] = xor_out[90][21][12] + xor_out[91][21][12] + xor_out[92][21][12] + xor_out[93][21][12] + xor_out[94][21][12];
assign sum_out[19][21][12] = xor_out[95][21][12] + xor_out[96][21][12] + xor_out[97][21][12] + xor_out[98][21][12] + xor_out[99][21][12];

assign sum_out[0][21][13] = xor_out[0][21][13] + xor_out[1][21][13] + xor_out[2][21][13] + xor_out[3][21][13] + xor_out[4][21][13];
assign sum_out[1][21][13] = xor_out[5][21][13] + xor_out[6][21][13] + xor_out[7][21][13] + xor_out[8][21][13] + xor_out[9][21][13];
assign sum_out[2][21][13] = xor_out[10][21][13] + xor_out[11][21][13] + xor_out[12][21][13] + xor_out[13][21][13] + xor_out[14][21][13];
assign sum_out[3][21][13] = xor_out[15][21][13] + xor_out[16][21][13] + xor_out[17][21][13] + xor_out[18][21][13] + xor_out[19][21][13];
assign sum_out[4][21][13] = xor_out[20][21][13] + xor_out[21][21][13] + xor_out[22][21][13] + xor_out[23][21][13] + xor_out[24][21][13];
assign sum_out[5][21][13] = xor_out[25][21][13] + xor_out[26][21][13] + xor_out[27][21][13] + xor_out[28][21][13] + xor_out[29][21][13];
assign sum_out[6][21][13] = xor_out[30][21][13] + xor_out[31][21][13] + xor_out[32][21][13] + xor_out[33][21][13] + xor_out[34][21][13];
assign sum_out[7][21][13] = xor_out[35][21][13] + xor_out[36][21][13] + xor_out[37][21][13] + xor_out[38][21][13] + xor_out[39][21][13];
assign sum_out[8][21][13] = xor_out[40][21][13] + xor_out[41][21][13] + xor_out[42][21][13] + xor_out[43][21][13] + xor_out[44][21][13];
assign sum_out[9][21][13] = xor_out[45][21][13] + xor_out[46][21][13] + xor_out[47][21][13] + xor_out[48][21][13] + xor_out[49][21][13];
assign sum_out[10][21][13] = xor_out[50][21][13] + xor_out[51][21][13] + xor_out[52][21][13] + xor_out[53][21][13] + xor_out[54][21][13];
assign sum_out[11][21][13] = xor_out[55][21][13] + xor_out[56][21][13] + xor_out[57][21][13] + xor_out[58][21][13] + xor_out[59][21][13];
assign sum_out[12][21][13] = xor_out[60][21][13] + xor_out[61][21][13] + xor_out[62][21][13] + xor_out[63][21][13] + xor_out[64][21][13];
assign sum_out[13][21][13] = xor_out[65][21][13] + xor_out[66][21][13] + xor_out[67][21][13] + xor_out[68][21][13] + xor_out[69][21][13];
assign sum_out[14][21][13] = xor_out[70][21][13] + xor_out[71][21][13] + xor_out[72][21][13] + xor_out[73][21][13] + xor_out[74][21][13];
assign sum_out[15][21][13] = xor_out[75][21][13] + xor_out[76][21][13] + xor_out[77][21][13] + xor_out[78][21][13] + xor_out[79][21][13];
assign sum_out[16][21][13] = xor_out[80][21][13] + xor_out[81][21][13] + xor_out[82][21][13] + xor_out[83][21][13] + xor_out[84][21][13];
assign sum_out[17][21][13] = xor_out[85][21][13] + xor_out[86][21][13] + xor_out[87][21][13] + xor_out[88][21][13] + xor_out[89][21][13];
assign sum_out[18][21][13] = xor_out[90][21][13] + xor_out[91][21][13] + xor_out[92][21][13] + xor_out[93][21][13] + xor_out[94][21][13];
assign sum_out[19][21][13] = xor_out[95][21][13] + xor_out[96][21][13] + xor_out[97][21][13] + xor_out[98][21][13] + xor_out[99][21][13];

assign sum_out[0][21][14] = xor_out[0][21][14] + xor_out[1][21][14] + xor_out[2][21][14] + xor_out[3][21][14] + xor_out[4][21][14];
assign sum_out[1][21][14] = xor_out[5][21][14] + xor_out[6][21][14] + xor_out[7][21][14] + xor_out[8][21][14] + xor_out[9][21][14];
assign sum_out[2][21][14] = xor_out[10][21][14] + xor_out[11][21][14] + xor_out[12][21][14] + xor_out[13][21][14] + xor_out[14][21][14];
assign sum_out[3][21][14] = xor_out[15][21][14] + xor_out[16][21][14] + xor_out[17][21][14] + xor_out[18][21][14] + xor_out[19][21][14];
assign sum_out[4][21][14] = xor_out[20][21][14] + xor_out[21][21][14] + xor_out[22][21][14] + xor_out[23][21][14] + xor_out[24][21][14];
assign sum_out[5][21][14] = xor_out[25][21][14] + xor_out[26][21][14] + xor_out[27][21][14] + xor_out[28][21][14] + xor_out[29][21][14];
assign sum_out[6][21][14] = xor_out[30][21][14] + xor_out[31][21][14] + xor_out[32][21][14] + xor_out[33][21][14] + xor_out[34][21][14];
assign sum_out[7][21][14] = xor_out[35][21][14] + xor_out[36][21][14] + xor_out[37][21][14] + xor_out[38][21][14] + xor_out[39][21][14];
assign sum_out[8][21][14] = xor_out[40][21][14] + xor_out[41][21][14] + xor_out[42][21][14] + xor_out[43][21][14] + xor_out[44][21][14];
assign sum_out[9][21][14] = xor_out[45][21][14] + xor_out[46][21][14] + xor_out[47][21][14] + xor_out[48][21][14] + xor_out[49][21][14];
assign sum_out[10][21][14] = xor_out[50][21][14] + xor_out[51][21][14] + xor_out[52][21][14] + xor_out[53][21][14] + xor_out[54][21][14];
assign sum_out[11][21][14] = xor_out[55][21][14] + xor_out[56][21][14] + xor_out[57][21][14] + xor_out[58][21][14] + xor_out[59][21][14];
assign sum_out[12][21][14] = xor_out[60][21][14] + xor_out[61][21][14] + xor_out[62][21][14] + xor_out[63][21][14] + xor_out[64][21][14];
assign sum_out[13][21][14] = xor_out[65][21][14] + xor_out[66][21][14] + xor_out[67][21][14] + xor_out[68][21][14] + xor_out[69][21][14];
assign sum_out[14][21][14] = xor_out[70][21][14] + xor_out[71][21][14] + xor_out[72][21][14] + xor_out[73][21][14] + xor_out[74][21][14];
assign sum_out[15][21][14] = xor_out[75][21][14] + xor_out[76][21][14] + xor_out[77][21][14] + xor_out[78][21][14] + xor_out[79][21][14];
assign sum_out[16][21][14] = xor_out[80][21][14] + xor_out[81][21][14] + xor_out[82][21][14] + xor_out[83][21][14] + xor_out[84][21][14];
assign sum_out[17][21][14] = xor_out[85][21][14] + xor_out[86][21][14] + xor_out[87][21][14] + xor_out[88][21][14] + xor_out[89][21][14];
assign sum_out[18][21][14] = xor_out[90][21][14] + xor_out[91][21][14] + xor_out[92][21][14] + xor_out[93][21][14] + xor_out[94][21][14];
assign sum_out[19][21][14] = xor_out[95][21][14] + xor_out[96][21][14] + xor_out[97][21][14] + xor_out[98][21][14] + xor_out[99][21][14];

assign sum_out[0][21][15] = xor_out[0][21][15] + xor_out[1][21][15] + xor_out[2][21][15] + xor_out[3][21][15] + xor_out[4][21][15];
assign sum_out[1][21][15] = xor_out[5][21][15] + xor_out[6][21][15] + xor_out[7][21][15] + xor_out[8][21][15] + xor_out[9][21][15];
assign sum_out[2][21][15] = xor_out[10][21][15] + xor_out[11][21][15] + xor_out[12][21][15] + xor_out[13][21][15] + xor_out[14][21][15];
assign sum_out[3][21][15] = xor_out[15][21][15] + xor_out[16][21][15] + xor_out[17][21][15] + xor_out[18][21][15] + xor_out[19][21][15];
assign sum_out[4][21][15] = xor_out[20][21][15] + xor_out[21][21][15] + xor_out[22][21][15] + xor_out[23][21][15] + xor_out[24][21][15];
assign sum_out[5][21][15] = xor_out[25][21][15] + xor_out[26][21][15] + xor_out[27][21][15] + xor_out[28][21][15] + xor_out[29][21][15];
assign sum_out[6][21][15] = xor_out[30][21][15] + xor_out[31][21][15] + xor_out[32][21][15] + xor_out[33][21][15] + xor_out[34][21][15];
assign sum_out[7][21][15] = xor_out[35][21][15] + xor_out[36][21][15] + xor_out[37][21][15] + xor_out[38][21][15] + xor_out[39][21][15];
assign sum_out[8][21][15] = xor_out[40][21][15] + xor_out[41][21][15] + xor_out[42][21][15] + xor_out[43][21][15] + xor_out[44][21][15];
assign sum_out[9][21][15] = xor_out[45][21][15] + xor_out[46][21][15] + xor_out[47][21][15] + xor_out[48][21][15] + xor_out[49][21][15];
assign sum_out[10][21][15] = xor_out[50][21][15] + xor_out[51][21][15] + xor_out[52][21][15] + xor_out[53][21][15] + xor_out[54][21][15];
assign sum_out[11][21][15] = xor_out[55][21][15] + xor_out[56][21][15] + xor_out[57][21][15] + xor_out[58][21][15] + xor_out[59][21][15];
assign sum_out[12][21][15] = xor_out[60][21][15] + xor_out[61][21][15] + xor_out[62][21][15] + xor_out[63][21][15] + xor_out[64][21][15];
assign sum_out[13][21][15] = xor_out[65][21][15] + xor_out[66][21][15] + xor_out[67][21][15] + xor_out[68][21][15] + xor_out[69][21][15];
assign sum_out[14][21][15] = xor_out[70][21][15] + xor_out[71][21][15] + xor_out[72][21][15] + xor_out[73][21][15] + xor_out[74][21][15];
assign sum_out[15][21][15] = xor_out[75][21][15] + xor_out[76][21][15] + xor_out[77][21][15] + xor_out[78][21][15] + xor_out[79][21][15];
assign sum_out[16][21][15] = xor_out[80][21][15] + xor_out[81][21][15] + xor_out[82][21][15] + xor_out[83][21][15] + xor_out[84][21][15];
assign sum_out[17][21][15] = xor_out[85][21][15] + xor_out[86][21][15] + xor_out[87][21][15] + xor_out[88][21][15] + xor_out[89][21][15];
assign sum_out[18][21][15] = xor_out[90][21][15] + xor_out[91][21][15] + xor_out[92][21][15] + xor_out[93][21][15] + xor_out[94][21][15];
assign sum_out[19][21][15] = xor_out[95][21][15] + xor_out[96][21][15] + xor_out[97][21][15] + xor_out[98][21][15] + xor_out[99][21][15];

assign sum_out[0][21][16] = xor_out[0][21][16] + xor_out[1][21][16] + xor_out[2][21][16] + xor_out[3][21][16] + xor_out[4][21][16];
assign sum_out[1][21][16] = xor_out[5][21][16] + xor_out[6][21][16] + xor_out[7][21][16] + xor_out[8][21][16] + xor_out[9][21][16];
assign sum_out[2][21][16] = xor_out[10][21][16] + xor_out[11][21][16] + xor_out[12][21][16] + xor_out[13][21][16] + xor_out[14][21][16];
assign sum_out[3][21][16] = xor_out[15][21][16] + xor_out[16][21][16] + xor_out[17][21][16] + xor_out[18][21][16] + xor_out[19][21][16];
assign sum_out[4][21][16] = xor_out[20][21][16] + xor_out[21][21][16] + xor_out[22][21][16] + xor_out[23][21][16] + xor_out[24][21][16];
assign sum_out[5][21][16] = xor_out[25][21][16] + xor_out[26][21][16] + xor_out[27][21][16] + xor_out[28][21][16] + xor_out[29][21][16];
assign sum_out[6][21][16] = xor_out[30][21][16] + xor_out[31][21][16] + xor_out[32][21][16] + xor_out[33][21][16] + xor_out[34][21][16];
assign sum_out[7][21][16] = xor_out[35][21][16] + xor_out[36][21][16] + xor_out[37][21][16] + xor_out[38][21][16] + xor_out[39][21][16];
assign sum_out[8][21][16] = xor_out[40][21][16] + xor_out[41][21][16] + xor_out[42][21][16] + xor_out[43][21][16] + xor_out[44][21][16];
assign sum_out[9][21][16] = xor_out[45][21][16] + xor_out[46][21][16] + xor_out[47][21][16] + xor_out[48][21][16] + xor_out[49][21][16];
assign sum_out[10][21][16] = xor_out[50][21][16] + xor_out[51][21][16] + xor_out[52][21][16] + xor_out[53][21][16] + xor_out[54][21][16];
assign sum_out[11][21][16] = xor_out[55][21][16] + xor_out[56][21][16] + xor_out[57][21][16] + xor_out[58][21][16] + xor_out[59][21][16];
assign sum_out[12][21][16] = xor_out[60][21][16] + xor_out[61][21][16] + xor_out[62][21][16] + xor_out[63][21][16] + xor_out[64][21][16];
assign sum_out[13][21][16] = xor_out[65][21][16] + xor_out[66][21][16] + xor_out[67][21][16] + xor_out[68][21][16] + xor_out[69][21][16];
assign sum_out[14][21][16] = xor_out[70][21][16] + xor_out[71][21][16] + xor_out[72][21][16] + xor_out[73][21][16] + xor_out[74][21][16];
assign sum_out[15][21][16] = xor_out[75][21][16] + xor_out[76][21][16] + xor_out[77][21][16] + xor_out[78][21][16] + xor_out[79][21][16];
assign sum_out[16][21][16] = xor_out[80][21][16] + xor_out[81][21][16] + xor_out[82][21][16] + xor_out[83][21][16] + xor_out[84][21][16];
assign sum_out[17][21][16] = xor_out[85][21][16] + xor_out[86][21][16] + xor_out[87][21][16] + xor_out[88][21][16] + xor_out[89][21][16];
assign sum_out[18][21][16] = xor_out[90][21][16] + xor_out[91][21][16] + xor_out[92][21][16] + xor_out[93][21][16] + xor_out[94][21][16];
assign sum_out[19][21][16] = xor_out[95][21][16] + xor_out[96][21][16] + xor_out[97][21][16] + xor_out[98][21][16] + xor_out[99][21][16];

assign sum_out[0][21][17] = xor_out[0][21][17] + xor_out[1][21][17] + xor_out[2][21][17] + xor_out[3][21][17] + xor_out[4][21][17];
assign sum_out[1][21][17] = xor_out[5][21][17] + xor_out[6][21][17] + xor_out[7][21][17] + xor_out[8][21][17] + xor_out[9][21][17];
assign sum_out[2][21][17] = xor_out[10][21][17] + xor_out[11][21][17] + xor_out[12][21][17] + xor_out[13][21][17] + xor_out[14][21][17];
assign sum_out[3][21][17] = xor_out[15][21][17] + xor_out[16][21][17] + xor_out[17][21][17] + xor_out[18][21][17] + xor_out[19][21][17];
assign sum_out[4][21][17] = xor_out[20][21][17] + xor_out[21][21][17] + xor_out[22][21][17] + xor_out[23][21][17] + xor_out[24][21][17];
assign sum_out[5][21][17] = xor_out[25][21][17] + xor_out[26][21][17] + xor_out[27][21][17] + xor_out[28][21][17] + xor_out[29][21][17];
assign sum_out[6][21][17] = xor_out[30][21][17] + xor_out[31][21][17] + xor_out[32][21][17] + xor_out[33][21][17] + xor_out[34][21][17];
assign sum_out[7][21][17] = xor_out[35][21][17] + xor_out[36][21][17] + xor_out[37][21][17] + xor_out[38][21][17] + xor_out[39][21][17];
assign sum_out[8][21][17] = xor_out[40][21][17] + xor_out[41][21][17] + xor_out[42][21][17] + xor_out[43][21][17] + xor_out[44][21][17];
assign sum_out[9][21][17] = xor_out[45][21][17] + xor_out[46][21][17] + xor_out[47][21][17] + xor_out[48][21][17] + xor_out[49][21][17];
assign sum_out[10][21][17] = xor_out[50][21][17] + xor_out[51][21][17] + xor_out[52][21][17] + xor_out[53][21][17] + xor_out[54][21][17];
assign sum_out[11][21][17] = xor_out[55][21][17] + xor_out[56][21][17] + xor_out[57][21][17] + xor_out[58][21][17] + xor_out[59][21][17];
assign sum_out[12][21][17] = xor_out[60][21][17] + xor_out[61][21][17] + xor_out[62][21][17] + xor_out[63][21][17] + xor_out[64][21][17];
assign sum_out[13][21][17] = xor_out[65][21][17] + xor_out[66][21][17] + xor_out[67][21][17] + xor_out[68][21][17] + xor_out[69][21][17];
assign sum_out[14][21][17] = xor_out[70][21][17] + xor_out[71][21][17] + xor_out[72][21][17] + xor_out[73][21][17] + xor_out[74][21][17];
assign sum_out[15][21][17] = xor_out[75][21][17] + xor_out[76][21][17] + xor_out[77][21][17] + xor_out[78][21][17] + xor_out[79][21][17];
assign sum_out[16][21][17] = xor_out[80][21][17] + xor_out[81][21][17] + xor_out[82][21][17] + xor_out[83][21][17] + xor_out[84][21][17];
assign sum_out[17][21][17] = xor_out[85][21][17] + xor_out[86][21][17] + xor_out[87][21][17] + xor_out[88][21][17] + xor_out[89][21][17];
assign sum_out[18][21][17] = xor_out[90][21][17] + xor_out[91][21][17] + xor_out[92][21][17] + xor_out[93][21][17] + xor_out[94][21][17];
assign sum_out[19][21][17] = xor_out[95][21][17] + xor_out[96][21][17] + xor_out[97][21][17] + xor_out[98][21][17] + xor_out[99][21][17];

assign sum_out[0][21][18] = xor_out[0][21][18] + xor_out[1][21][18] + xor_out[2][21][18] + xor_out[3][21][18] + xor_out[4][21][18];
assign sum_out[1][21][18] = xor_out[5][21][18] + xor_out[6][21][18] + xor_out[7][21][18] + xor_out[8][21][18] + xor_out[9][21][18];
assign sum_out[2][21][18] = xor_out[10][21][18] + xor_out[11][21][18] + xor_out[12][21][18] + xor_out[13][21][18] + xor_out[14][21][18];
assign sum_out[3][21][18] = xor_out[15][21][18] + xor_out[16][21][18] + xor_out[17][21][18] + xor_out[18][21][18] + xor_out[19][21][18];
assign sum_out[4][21][18] = xor_out[20][21][18] + xor_out[21][21][18] + xor_out[22][21][18] + xor_out[23][21][18] + xor_out[24][21][18];
assign sum_out[5][21][18] = xor_out[25][21][18] + xor_out[26][21][18] + xor_out[27][21][18] + xor_out[28][21][18] + xor_out[29][21][18];
assign sum_out[6][21][18] = xor_out[30][21][18] + xor_out[31][21][18] + xor_out[32][21][18] + xor_out[33][21][18] + xor_out[34][21][18];
assign sum_out[7][21][18] = xor_out[35][21][18] + xor_out[36][21][18] + xor_out[37][21][18] + xor_out[38][21][18] + xor_out[39][21][18];
assign sum_out[8][21][18] = xor_out[40][21][18] + xor_out[41][21][18] + xor_out[42][21][18] + xor_out[43][21][18] + xor_out[44][21][18];
assign sum_out[9][21][18] = xor_out[45][21][18] + xor_out[46][21][18] + xor_out[47][21][18] + xor_out[48][21][18] + xor_out[49][21][18];
assign sum_out[10][21][18] = xor_out[50][21][18] + xor_out[51][21][18] + xor_out[52][21][18] + xor_out[53][21][18] + xor_out[54][21][18];
assign sum_out[11][21][18] = xor_out[55][21][18] + xor_out[56][21][18] + xor_out[57][21][18] + xor_out[58][21][18] + xor_out[59][21][18];
assign sum_out[12][21][18] = xor_out[60][21][18] + xor_out[61][21][18] + xor_out[62][21][18] + xor_out[63][21][18] + xor_out[64][21][18];
assign sum_out[13][21][18] = xor_out[65][21][18] + xor_out[66][21][18] + xor_out[67][21][18] + xor_out[68][21][18] + xor_out[69][21][18];
assign sum_out[14][21][18] = xor_out[70][21][18] + xor_out[71][21][18] + xor_out[72][21][18] + xor_out[73][21][18] + xor_out[74][21][18];
assign sum_out[15][21][18] = xor_out[75][21][18] + xor_out[76][21][18] + xor_out[77][21][18] + xor_out[78][21][18] + xor_out[79][21][18];
assign sum_out[16][21][18] = xor_out[80][21][18] + xor_out[81][21][18] + xor_out[82][21][18] + xor_out[83][21][18] + xor_out[84][21][18];
assign sum_out[17][21][18] = xor_out[85][21][18] + xor_out[86][21][18] + xor_out[87][21][18] + xor_out[88][21][18] + xor_out[89][21][18];
assign sum_out[18][21][18] = xor_out[90][21][18] + xor_out[91][21][18] + xor_out[92][21][18] + xor_out[93][21][18] + xor_out[94][21][18];
assign sum_out[19][21][18] = xor_out[95][21][18] + xor_out[96][21][18] + xor_out[97][21][18] + xor_out[98][21][18] + xor_out[99][21][18];

assign sum_out[0][21][19] = xor_out[0][21][19] + xor_out[1][21][19] + xor_out[2][21][19] + xor_out[3][21][19] + xor_out[4][21][19];
assign sum_out[1][21][19] = xor_out[5][21][19] + xor_out[6][21][19] + xor_out[7][21][19] + xor_out[8][21][19] + xor_out[9][21][19];
assign sum_out[2][21][19] = xor_out[10][21][19] + xor_out[11][21][19] + xor_out[12][21][19] + xor_out[13][21][19] + xor_out[14][21][19];
assign sum_out[3][21][19] = xor_out[15][21][19] + xor_out[16][21][19] + xor_out[17][21][19] + xor_out[18][21][19] + xor_out[19][21][19];
assign sum_out[4][21][19] = xor_out[20][21][19] + xor_out[21][21][19] + xor_out[22][21][19] + xor_out[23][21][19] + xor_out[24][21][19];
assign sum_out[5][21][19] = xor_out[25][21][19] + xor_out[26][21][19] + xor_out[27][21][19] + xor_out[28][21][19] + xor_out[29][21][19];
assign sum_out[6][21][19] = xor_out[30][21][19] + xor_out[31][21][19] + xor_out[32][21][19] + xor_out[33][21][19] + xor_out[34][21][19];
assign sum_out[7][21][19] = xor_out[35][21][19] + xor_out[36][21][19] + xor_out[37][21][19] + xor_out[38][21][19] + xor_out[39][21][19];
assign sum_out[8][21][19] = xor_out[40][21][19] + xor_out[41][21][19] + xor_out[42][21][19] + xor_out[43][21][19] + xor_out[44][21][19];
assign sum_out[9][21][19] = xor_out[45][21][19] + xor_out[46][21][19] + xor_out[47][21][19] + xor_out[48][21][19] + xor_out[49][21][19];
assign sum_out[10][21][19] = xor_out[50][21][19] + xor_out[51][21][19] + xor_out[52][21][19] + xor_out[53][21][19] + xor_out[54][21][19];
assign sum_out[11][21][19] = xor_out[55][21][19] + xor_out[56][21][19] + xor_out[57][21][19] + xor_out[58][21][19] + xor_out[59][21][19];
assign sum_out[12][21][19] = xor_out[60][21][19] + xor_out[61][21][19] + xor_out[62][21][19] + xor_out[63][21][19] + xor_out[64][21][19];
assign sum_out[13][21][19] = xor_out[65][21][19] + xor_out[66][21][19] + xor_out[67][21][19] + xor_out[68][21][19] + xor_out[69][21][19];
assign sum_out[14][21][19] = xor_out[70][21][19] + xor_out[71][21][19] + xor_out[72][21][19] + xor_out[73][21][19] + xor_out[74][21][19];
assign sum_out[15][21][19] = xor_out[75][21][19] + xor_out[76][21][19] + xor_out[77][21][19] + xor_out[78][21][19] + xor_out[79][21][19];
assign sum_out[16][21][19] = xor_out[80][21][19] + xor_out[81][21][19] + xor_out[82][21][19] + xor_out[83][21][19] + xor_out[84][21][19];
assign sum_out[17][21][19] = xor_out[85][21][19] + xor_out[86][21][19] + xor_out[87][21][19] + xor_out[88][21][19] + xor_out[89][21][19];
assign sum_out[18][21][19] = xor_out[90][21][19] + xor_out[91][21][19] + xor_out[92][21][19] + xor_out[93][21][19] + xor_out[94][21][19];
assign sum_out[19][21][19] = xor_out[95][21][19] + xor_out[96][21][19] + xor_out[97][21][19] + xor_out[98][21][19] + xor_out[99][21][19];

assign sum_out[0][21][20] = xor_out[0][21][20] + xor_out[1][21][20] + xor_out[2][21][20] + xor_out[3][21][20] + xor_out[4][21][20];
assign sum_out[1][21][20] = xor_out[5][21][20] + xor_out[6][21][20] + xor_out[7][21][20] + xor_out[8][21][20] + xor_out[9][21][20];
assign sum_out[2][21][20] = xor_out[10][21][20] + xor_out[11][21][20] + xor_out[12][21][20] + xor_out[13][21][20] + xor_out[14][21][20];
assign sum_out[3][21][20] = xor_out[15][21][20] + xor_out[16][21][20] + xor_out[17][21][20] + xor_out[18][21][20] + xor_out[19][21][20];
assign sum_out[4][21][20] = xor_out[20][21][20] + xor_out[21][21][20] + xor_out[22][21][20] + xor_out[23][21][20] + xor_out[24][21][20];
assign sum_out[5][21][20] = xor_out[25][21][20] + xor_out[26][21][20] + xor_out[27][21][20] + xor_out[28][21][20] + xor_out[29][21][20];
assign sum_out[6][21][20] = xor_out[30][21][20] + xor_out[31][21][20] + xor_out[32][21][20] + xor_out[33][21][20] + xor_out[34][21][20];
assign sum_out[7][21][20] = xor_out[35][21][20] + xor_out[36][21][20] + xor_out[37][21][20] + xor_out[38][21][20] + xor_out[39][21][20];
assign sum_out[8][21][20] = xor_out[40][21][20] + xor_out[41][21][20] + xor_out[42][21][20] + xor_out[43][21][20] + xor_out[44][21][20];
assign sum_out[9][21][20] = xor_out[45][21][20] + xor_out[46][21][20] + xor_out[47][21][20] + xor_out[48][21][20] + xor_out[49][21][20];
assign sum_out[10][21][20] = xor_out[50][21][20] + xor_out[51][21][20] + xor_out[52][21][20] + xor_out[53][21][20] + xor_out[54][21][20];
assign sum_out[11][21][20] = xor_out[55][21][20] + xor_out[56][21][20] + xor_out[57][21][20] + xor_out[58][21][20] + xor_out[59][21][20];
assign sum_out[12][21][20] = xor_out[60][21][20] + xor_out[61][21][20] + xor_out[62][21][20] + xor_out[63][21][20] + xor_out[64][21][20];
assign sum_out[13][21][20] = xor_out[65][21][20] + xor_out[66][21][20] + xor_out[67][21][20] + xor_out[68][21][20] + xor_out[69][21][20];
assign sum_out[14][21][20] = xor_out[70][21][20] + xor_out[71][21][20] + xor_out[72][21][20] + xor_out[73][21][20] + xor_out[74][21][20];
assign sum_out[15][21][20] = xor_out[75][21][20] + xor_out[76][21][20] + xor_out[77][21][20] + xor_out[78][21][20] + xor_out[79][21][20];
assign sum_out[16][21][20] = xor_out[80][21][20] + xor_out[81][21][20] + xor_out[82][21][20] + xor_out[83][21][20] + xor_out[84][21][20];
assign sum_out[17][21][20] = xor_out[85][21][20] + xor_out[86][21][20] + xor_out[87][21][20] + xor_out[88][21][20] + xor_out[89][21][20];
assign sum_out[18][21][20] = xor_out[90][21][20] + xor_out[91][21][20] + xor_out[92][21][20] + xor_out[93][21][20] + xor_out[94][21][20];
assign sum_out[19][21][20] = xor_out[95][21][20] + xor_out[96][21][20] + xor_out[97][21][20] + xor_out[98][21][20] + xor_out[99][21][20];

assign sum_out[0][21][21] = xor_out[0][21][21] + xor_out[1][21][21] + xor_out[2][21][21] + xor_out[3][21][21] + xor_out[4][21][21];
assign sum_out[1][21][21] = xor_out[5][21][21] + xor_out[6][21][21] + xor_out[7][21][21] + xor_out[8][21][21] + xor_out[9][21][21];
assign sum_out[2][21][21] = xor_out[10][21][21] + xor_out[11][21][21] + xor_out[12][21][21] + xor_out[13][21][21] + xor_out[14][21][21];
assign sum_out[3][21][21] = xor_out[15][21][21] + xor_out[16][21][21] + xor_out[17][21][21] + xor_out[18][21][21] + xor_out[19][21][21];
assign sum_out[4][21][21] = xor_out[20][21][21] + xor_out[21][21][21] + xor_out[22][21][21] + xor_out[23][21][21] + xor_out[24][21][21];
assign sum_out[5][21][21] = xor_out[25][21][21] + xor_out[26][21][21] + xor_out[27][21][21] + xor_out[28][21][21] + xor_out[29][21][21];
assign sum_out[6][21][21] = xor_out[30][21][21] + xor_out[31][21][21] + xor_out[32][21][21] + xor_out[33][21][21] + xor_out[34][21][21];
assign sum_out[7][21][21] = xor_out[35][21][21] + xor_out[36][21][21] + xor_out[37][21][21] + xor_out[38][21][21] + xor_out[39][21][21];
assign sum_out[8][21][21] = xor_out[40][21][21] + xor_out[41][21][21] + xor_out[42][21][21] + xor_out[43][21][21] + xor_out[44][21][21];
assign sum_out[9][21][21] = xor_out[45][21][21] + xor_out[46][21][21] + xor_out[47][21][21] + xor_out[48][21][21] + xor_out[49][21][21];
assign sum_out[10][21][21] = xor_out[50][21][21] + xor_out[51][21][21] + xor_out[52][21][21] + xor_out[53][21][21] + xor_out[54][21][21];
assign sum_out[11][21][21] = xor_out[55][21][21] + xor_out[56][21][21] + xor_out[57][21][21] + xor_out[58][21][21] + xor_out[59][21][21];
assign sum_out[12][21][21] = xor_out[60][21][21] + xor_out[61][21][21] + xor_out[62][21][21] + xor_out[63][21][21] + xor_out[64][21][21];
assign sum_out[13][21][21] = xor_out[65][21][21] + xor_out[66][21][21] + xor_out[67][21][21] + xor_out[68][21][21] + xor_out[69][21][21];
assign sum_out[14][21][21] = xor_out[70][21][21] + xor_out[71][21][21] + xor_out[72][21][21] + xor_out[73][21][21] + xor_out[74][21][21];
assign sum_out[15][21][21] = xor_out[75][21][21] + xor_out[76][21][21] + xor_out[77][21][21] + xor_out[78][21][21] + xor_out[79][21][21];
assign sum_out[16][21][21] = xor_out[80][21][21] + xor_out[81][21][21] + xor_out[82][21][21] + xor_out[83][21][21] + xor_out[84][21][21];
assign sum_out[17][21][21] = xor_out[85][21][21] + xor_out[86][21][21] + xor_out[87][21][21] + xor_out[88][21][21] + xor_out[89][21][21];
assign sum_out[18][21][21] = xor_out[90][21][21] + xor_out[91][21][21] + xor_out[92][21][21] + xor_out[93][21][21] + xor_out[94][21][21];
assign sum_out[19][21][21] = xor_out[95][21][21] + xor_out[96][21][21] + xor_out[97][21][21] + xor_out[98][21][21] + xor_out[99][21][21];

assign sum_out[0][21][22] = xor_out[0][21][22] + xor_out[1][21][22] + xor_out[2][21][22] + xor_out[3][21][22] + xor_out[4][21][22];
assign sum_out[1][21][22] = xor_out[5][21][22] + xor_out[6][21][22] + xor_out[7][21][22] + xor_out[8][21][22] + xor_out[9][21][22];
assign sum_out[2][21][22] = xor_out[10][21][22] + xor_out[11][21][22] + xor_out[12][21][22] + xor_out[13][21][22] + xor_out[14][21][22];
assign sum_out[3][21][22] = xor_out[15][21][22] + xor_out[16][21][22] + xor_out[17][21][22] + xor_out[18][21][22] + xor_out[19][21][22];
assign sum_out[4][21][22] = xor_out[20][21][22] + xor_out[21][21][22] + xor_out[22][21][22] + xor_out[23][21][22] + xor_out[24][21][22];
assign sum_out[5][21][22] = xor_out[25][21][22] + xor_out[26][21][22] + xor_out[27][21][22] + xor_out[28][21][22] + xor_out[29][21][22];
assign sum_out[6][21][22] = xor_out[30][21][22] + xor_out[31][21][22] + xor_out[32][21][22] + xor_out[33][21][22] + xor_out[34][21][22];
assign sum_out[7][21][22] = xor_out[35][21][22] + xor_out[36][21][22] + xor_out[37][21][22] + xor_out[38][21][22] + xor_out[39][21][22];
assign sum_out[8][21][22] = xor_out[40][21][22] + xor_out[41][21][22] + xor_out[42][21][22] + xor_out[43][21][22] + xor_out[44][21][22];
assign sum_out[9][21][22] = xor_out[45][21][22] + xor_out[46][21][22] + xor_out[47][21][22] + xor_out[48][21][22] + xor_out[49][21][22];
assign sum_out[10][21][22] = xor_out[50][21][22] + xor_out[51][21][22] + xor_out[52][21][22] + xor_out[53][21][22] + xor_out[54][21][22];
assign sum_out[11][21][22] = xor_out[55][21][22] + xor_out[56][21][22] + xor_out[57][21][22] + xor_out[58][21][22] + xor_out[59][21][22];
assign sum_out[12][21][22] = xor_out[60][21][22] + xor_out[61][21][22] + xor_out[62][21][22] + xor_out[63][21][22] + xor_out[64][21][22];
assign sum_out[13][21][22] = xor_out[65][21][22] + xor_out[66][21][22] + xor_out[67][21][22] + xor_out[68][21][22] + xor_out[69][21][22];
assign sum_out[14][21][22] = xor_out[70][21][22] + xor_out[71][21][22] + xor_out[72][21][22] + xor_out[73][21][22] + xor_out[74][21][22];
assign sum_out[15][21][22] = xor_out[75][21][22] + xor_out[76][21][22] + xor_out[77][21][22] + xor_out[78][21][22] + xor_out[79][21][22];
assign sum_out[16][21][22] = xor_out[80][21][22] + xor_out[81][21][22] + xor_out[82][21][22] + xor_out[83][21][22] + xor_out[84][21][22];
assign sum_out[17][21][22] = xor_out[85][21][22] + xor_out[86][21][22] + xor_out[87][21][22] + xor_out[88][21][22] + xor_out[89][21][22];
assign sum_out[18][21][22] = xor_out[90][21][22] + xor_out[91][21][22] + xor_out[92][21][22] + xor_out[93][21][22] + xor_out[94][21][22];
assign sum_out[19][21][22] = xor_out[95][21][22] + xor_out[96][21][22] + xor_out[97][21][22] + xor_out[98][21][22] + xor_out[99][21][22];

assign sum_out[0][21][23] = xor_out[0][21][23] + xor_out[1][21][23] + xor_out[2][21][23] + xor_out[3][21][23] + xor_out[4][21][23];
assign sum_out[1][21][23] = xor_out[5][21][23] + xor_out[6][21][23] + xor_out[7][21][23] + xor_out[8][21][23] + xor_out[9][21][23];
assign sum_out[2][21][23] = xor_out[10][21][23] + xor_out[11][21][23] + xor_out[12][21][23] + xor_out[13][21][23] + xor_out[14][21][23];
assign sum_out[3][21][23] = xor_out[15][21][23] + xor_out[16][21][23] + xor_out[17][21][23] + xor_out[18][21][23] + xor_out[19][21][23];
assign sum_out[4][21][23] = xor_out[20][21][23] + xor_out[21][21][23] + xor_out[22][21][23] + xor_out[23][21][23] + xor_out[24][21][23];
assign sum_out[5][21][23] = xor_out[25][21][23] + xor_out[26][21][23] + xor_out[27][21][23] + xor_out[28][21][23] + xor_out[29][21][23];
assign sum_out[6][21][23] = xor_out[30][21][23] + xor_out[31][21][23] + xor_out[32][21][23] + xor_out[33][21][23] + xor_out[34][21][23];
assign sum_out[7][21][23] = xor_out[35][21][23] + xor_out[36][21][23] + xor_out[37][21][23] + xor_out[38][21][23] + xor_out[39][21][23];
assign sum_out[8][21][23] = xor_out[40][21][23] + xor_out[41][21][23] + xor_out[42][21][23] + xor_out[43][21][23] + xor_out[44][21][23];
assign sum_out[9][21][23] = xor_out[45][21][23] + xor_out[46][21][23] + xor_out[47][21][23] + xor_out[48][21][23] + xor_out[49][21][23];
assign sum_out[10][21][23] = xor_out[50][21][23] + xor_out[51][21][23] + xor_out[52][21][23] + xor_out[53][21][23] + xor_out[54][21][23];
assign sum_out[11][21][23] = xor_out[55][21][23] + xor_out[56][21][23] + xor_out[57][21][23] + xor_out[58][21][23] + xor_out[59][21][23];
assign sum_out[12][21][23] = xor_out[60][21][23] + xor_out[61][21][23] + xor_out[62][21][23] + xor_out[63][21][23] + xor_out[64][21][23];
assign sum_out[13][21][23] = xor_out[65][21][23] + xor_out[66][21][23] + xor_out[67][21][23] + xor_out[68][21][23] + xor_out[69][21][23];
assign sum_out[14][21][23] = xor_out[70][21][23] + xor_out[71][21][23] + xor_out[72][21][23] + xor_out[73][21][23] + xor_out[74][21][23];
assign sum_out[15][21][23] = xor_out[75][21][23] + xor_out[76][21][23] + xor_out[77][21][23] + xor_out[78][21][23] + xor_out[79][21][23];
assign sum_out[16][21][23] = xor_out[80][21][23] + xor_out[81][21][23] + xor_out[82][21][23] + xor_out[83][21][23] + xor_out[84][21][23];
assign sum_out[17][21][23] = xor_out[85][21][23] + xor_out[86][21][23] + xor_out[87][21][23] + xor_out[88][21][23] + xor_out[89][21][23];
assign sum_out[18][21][23] = xor_out[90][21][23] + xor_out[91][21][23] + xor_out[92][21][23] + xor_out[93][21][23] + xor_out[94][21][23];
assign sum_out[19][21][23] = xor_out[95][21][23] + xor_out[96][21][23] + xor_out[97][21][23] + xor_out[98][21][23] + xor_out[99][21][23];

assign sum_out[0][22][0] = xor_out[0][22][0] + xor_out[1][22][0] + xor_out[2][22][0] + xor_out[3][22][0] + xor_out[4][22][0];
assign sum_out[1][22][0] = xor_out[5][22][0] + xor_out[6][22][0] + xor_out[7][22][0] + xor_out[8][22][0] + xor_out[9][22][0];
assign sum_out[2][22][0] = xor_out[10][22][0] + xor_out[11][22][0] + xor_out[12][22][0] + xor_out[13][22][0] + xor_out[14][22][0];
assign sum_out[3][22][0] = xor_out[15][22][0] + xor_out[16][22][0] + xor_out[17][22][0] + xor_out[18][22][0] + xor_out[19][22][0];
assign sum_out[4][22][0] = xor_out[20][22][0] + xor_out[21][22][0] + xor_out[22][22][0] + xor_out[23][22][0] + xor_out[24][22][0];
assign sum_out[5][22][0] = xor_out[25][22][0] + xor_out[26][22][0] + xor_out[27][22][0] + xor_out[28][22][0] + xor_out[29][22][0];
assign sum_out[6][22][0] = xor_out[30][22][0] + xor_out[31][22][0] + xor_out[32][22][0] + xor_out[33][22][0] + xor_out[34][22][0];
assign sum_out[7][22][0] = xor_out[35][22][0] + xor_out[36][22][0] + xor_out[37][22][0] + xor_out[38][22][0] + xor_out[39][22][0];
assign sum_out[8][22][0] = xor_out[40][22][0] + xor_out[41][22][0] + xor_out[42][22][0] + xor_out[43][22][0] + xor_out[44][22][0];
assign sum_out[9][22][0] = xor_out[45][22][0] + xor_out[46][22][0] + xor_out[47][22][0] + xor_out[48][22][0] + xor_out[49][22][0];
assign sum_out[10][22][0] = xor_out[50][22][0] + xor_out[51][22][0] + xor_out[52][22][0] + xor_out[53][22][0] + xor_out[54][22][0];
assign sum_out[11][22][0] = xor_out[55][22][0] + xor_out[56][22][0] + xor_out[57][22][0] + xor_out[58][22][0] + xor_out[59][22][0];
assign sum_out[12][22][0] = xor_out[60][22][0] + xor_out[61][22][0] + xor_out[62][22][0] + xor_out[63][22][0] + xor_out[64][22][0];
assign sum_out[13][22][0] = xor_out[65][22][0] + xor_out[66][22][0] + xor_out[67][22][0] + xor_out[68][22][0] + xor_out[69][22][0];
assign sum_out[14][22][0] = xor_out[70][22][0] + xor_out[71][22][0] + xor_out[72][22][0] + xor_out[73][22][0] + xor_out[74][22][0];
assign sum_out[15][22][0] = xor_out[75][22][0] + xor_out[76][22][0] + xor_out[77][22][0] + xor_out[78][22][0] + xor_out[79][22][0];
assign sum_out[16][22][0] = xor_out[80][22][0] + xor_out[81][22][0] + xor_out[82][22][0] + xor_out[83][22][0] + xor_out[84][22][0];
assign sum_out[17][22][0] = xor_out[85][22][0] + xor_out[86][22][0] + xor_out[87][22][0] + xor_out[88][22][0] + xor_out[89][22][0];
assign sum_out[18][22][0] = xor_out[90][22][0] + xor_out[91][22][0] + xor_out[92][22][0] + xor_out[93][22][0] + xor_out[94][22][0];
assign sum_out[19][22][0] = xor_out[95][22][0] + xor_out[96][22][0] + xor_out[97][22][0] + xor_out[98][22][0] + xor_out[99][22][0];

assign sum_out[0][22][1] = xor_out[0][22][1] + xor_out[1][22][1] + xor_out[2][22][1] + xor_out[3][22][1] + xor_out[4][22][1];
assign sum_out[1][22][1] = xor_out[5][22][1] + xor_out[6][22][1] + xor_out[7][22][1] + xor_out[8][22][1] + xor_out[9][22][1];
assign sum_out[2][22][1] = xor_out[10][22][1] + xor_out[11][22][1] + xor_out[12][22][1] + xor_out[13][22][1] + xor_out[14][22][1];
assign sum_out[3][22][1] = xor_out[15][22][1] + xor_out[16][22][1] + xor_out[17][22][1] + xor_out[18][22][1] + xor_out[19][22][1];
assign sum_out[4][22][1] = xor_out[20][22][1] + xor_out[21][22][1] + xor_out[22][22][1] + xor_out[23][22][1] + xor_out[24][22][1];
assign sum_out[5][22][1] = xor_out[25][22][1] + xor_out[26][22][1] + xor_out[27][22][1] + xor_out[28][22][1] + xor_out[29][22][1];
assign sum_out[6][22][1] = xor_out[30][22][1] + xor_out[31][22][1] + xor_out[32][22][1] + xor_out[33][22][1] + xor_out[34][22][1];
assign sum_out[7][22][1] = xor_out[35][22][1] + xor_out[36][22][1] + xor_out[37][22][1] + xor_out[38][22][1] + xor_out[39][22][1];
assign sum_out[8][22][1] = xor_out[40][22][1] + xor_out[41][22][1] + xor_out[42][22][1] + xor_out[43][22][1] + xor_out[44][22][1];
assign sum_out[9][22][1] = xor_out[45][22][1] + xor_out[46][22][1] + xor_out[47][22][1] + xor_out[48][22][1] + xor_out[49][22][1];
assign sum_out[10][22][1] = xor_out[50][22][1] + xor_out[51][22][1] + xor_out[52][22][1] + xor_out[53][22][1] + xor_out[54][22][1];
assign sum_out[11][22][1] = xor_out[55][22][1] + xor_out[56][22][1] + xor_out[57][22][1] + xor_out[58][22][1] + xor_out[59][22][1];
assign sum_out[12][22][1] = xor_out[60][22][1] + xor_out[61][22][1] + xor_out[62][22][1] + xor_out[63][22][1] + xor_out[64][22][1];
assign sum_out[13][22][1] = xor_out[65][22][1] + xor_out[66][22][1] + xor_out[67][22][1] + xor_out[68][22][1] + xor_out[69][22][1];
assign sum_out[14][22][1] = xor_out[70][22][1] + xor_out[71][22][1] + xor_out[72][22][1] + xor_out[73][22][1] + xor_out[74][22][1];
assign sum_out[15][22][1] = xor_out[75][22][1] + xor_out[76][22][1] + xor_out[77][22][1] + xor_out[78][22][1] + xor_out[79][22][1];
assign sum_out[16][22][1] = xor_out[80][22][1] + xor_out[81][22][1] + xor_out[82][22][1] + xor_out[83][22][1] + xor_out[84][22][1];
assign sum_out[17][22][1] = xor_out[85][22][1] + xor_out[86][22][1] + xor_out[87][22][1] + xor_out[88][22][1] + xor_out[89][22][1];
assign sum_out[18][22][1] = xor_out[90][22][1] + xor_out[91][22][1] + xor_out[92][22][1] + xor_out[93][22][1] + xor_out[94][22][1];
assign sum_out[19][22][1] = xor_out[95][22][1] + xor_out[96][22][1] + xor_out[97][22][1] + xor_out[98][22][1] + xor_out[99][22][1];

assign sum_out[0][22][2] = xor_out[0][22][2] + xor_out[1][22][2] + xor_out[2][22][2] + xor_out[3][22][2] + xor_out[4][22][2];
assign sum_out[1][22][2] = xor_out[5][22][2] + xor_out[6][22][2] + xor_out[7][22][2] + xor_out[8][22][2] + xor_out[9][22][2];
assign sum_out[2][22][2] = xor_out[10][22][2] + xor_out[11][22][2] + xor_out[12][22][2] + xor_out[13][22][2] + xor_out[14][22][2];
assign sum_out[3][22][2] = xor_out[15][22][2] + xor_out[16][22][2] + xor_out[17][22][2] + xor_out[18][22][2] + xor_out[19][22][2];
assign sum_out[4][22][2] = xor_out[20][22][2] + xor_out[21][22][2] + xor_out[22][22][2] + xor_out[23][22][2] + xor_out[24][22][2];
assign sum_out[5][22][2] = xor_out[25][22][2] + xor_out[26][22][2] + xor_out[27][22][2] + xor_out[28][22][2] + xor_out[29][22][2];
assign sum_out[6][22][2] = xor_out[30][22][2] + xor_out[31][22][2] + xor_out[32][22][2] + xor_out[33][22][2] + xor_out[34][22][2];
assign sum_out[7][22][2] = xor_out[35][22][2] + xor_out[36][22][2] + xor_out[37][22][2] + xor_out[38][22][2] + xor_out[39][22][2];
assign sum_out[8][22][2] = xor_out[40][22][2] + xor_out[41][22][2] + xor_out[42][22][2] + xor_out[43][22][2] + xor_out[44][22][2];
assign sum_out[9][22][2] = xor_out[45][22][2] + xor_out[46][22][2] + xor_out[47][22][2] + xor_out[48][22][2] + xor_out[49][22][2];
assign sum_out[10][22][2] = xor_out[50][22][2] + xor_out[51][22][2] + xor_out[52][22][2] + xor_out[53][22][2] + xor_out[54][22][2];
assign sum_out[11][22][2] = xor_out[55][22][2] + xor_out[56][22][2] + xor_out[57][22][2] + xor_out[58][22][2] + xor_out[59][22][2];
assign sum_out[12][22][2] = xor_out[60][22][2] + xor_out[61][22][2] + xor_out[62][22][2] + xor_out[63][22][2] + xor_out[64][22][2];
assign sum_out[13][22][2] = xor_out[65][22][2] + xor_out[66][22][2] + xor_out[67][22][2] + xor_out[68][22][2] + xor_out[69][22][2];
assign sum_out[14][22][2] = xor_out[70][22][2] + xor_out[71][22][2] + xor_out[72][22][2] + xor_out[73][22][2] + xor_out[74][22][2];
assign sum_out[15][22][2] = xor_out[75][22][2] + xor_out[76][22][2] + xor_out[77][22][2] + xor_out[78][22][2] + xor_out[79][22][2];
assign sum_out[16][22][2] = xor_out[80][22][2] + xor_out[81][22][2] + xor_out[82][22][2] + xor_out[83][22][2] + xor_out[84][22][2];
assign sum_out[17][22][2] = xor_out[85][22][2] + xor_out[86][22][2] + xor_out[87][22][2] + xor_out[88][22][2] + xor_out[89][22][2];
assign sum_out[18][22][2] = xor_out[90][22][2] + xor_out[91][22][2] + xor_out[92][22][2] + xor_out[93][22][2] + xor_out[94][22][2];
assign sum_out[19][22][2] = xor_out[95][22][2] + xor_out[96][22][2] + xor_out[97][22][2] + xor_out[98][22][2] + xor_out[99][22][2];

assign sum_out[0][22][3] = xor_out[0][22][3] + xor_out[1][22][3] + xor_out[2][22][3] + xor_out[3][22][3] + xor_out[4][22][3];
assign sum_out[1][22][3] = xor_out[5][22][3] + xor_out[6][22][3] + xor_out[7][22][3] + xor_out[8][22][3] + xor_out[9][22][3];
assign sum_out[2][22][3] = xor_out[10][22][3] + xor_out[11][22][3] + xor_out[12][22][3] + xor_out[13][22][3] + xor_out[14][22][3];
assign sum_out[3][22][3] = xor_out[15][22][3] + xor_out[16][22][3] + xor_out[17][22][3] + xor_out[18][22][3] + xor_out[19][22][3];
assign sum_out[4][22][3] = xor_out[20][22][3] + xor_out[21][22][3] + xor_out[22][22][3] + xor_out[23][22][3] + xor_out[24][22][3];
assign sum_out[5][22][3] = xor_out[25][22][3] + xor_out[26][22][3] + xor_out[27][22][3] + xor_out[28][22][3] + xor_out[29][22][3];
assign sum_out[6][22][3] = xor_out[30][22][3] + xor_out[31][22][3] + xor_out[32][22][3] + xor_out[33][22][3] + xor_out[34][22][3];
assign sum_out[7][22][3] = xor_out[35][22][3] + xor_out[36][22][3] + xor_out[37][22][3] + xor_out[38][22][3] + xor_out[39][22][3];
assign sum_out[8][22][3] = xor_out[40][22][3] + xor_out[41][22][3] + xor_out[42][22][3] + xor_out[43][22][3] + xor_out[44][22][3];
assign sum_out[9][22][3] = xor_out[45][22][3] + xor_out[46][22][3] + xor_out[47][22][3] + xor_out[48][22][3] + xor_out[49][22][3];
assign sum_out[10][22][3] = xor_out[50][22][3] + xor_out[51][22][3] + xor_out[52][22][3] + xor_out[53][22][3] + xor_out[54][22][3];
assign sum_out[11][22][3] = xor_out[55][22][3] + xor_out[56][22][3] + xor_out[57][22][3] + xor_out[58][22][3] + xor_out[59][22][3];
assign sum_out[12][22][3] = xor_out[60][22][3] + xor_out[61][22][3] + xor_out[62][22][3] + xor_out[63][22][3] + xor_out[64][22][3];
assign sum_out[13][22][3] = xor_out[65][22][3] + xor_out[66][22][3] + xor_out[67][22][3] + xor_out[68][22][3] + xor_out[69][22][3];
assign sum_out[14][22][3] = xor_out[70][22][3] + xor_out[71][22][3] + xor_out[72][22][3] + xor_out[73][22][3] + xor_out[74][22][3];
assign sum_out[15][22][3] = xor_out[75][22][3] + xor_out[76][22][3] + xor_out[77][22][3] + xor_out[78][22][3] + xor_out[79][22][3];
assign sum_out[16][22][3] = xor_out[80][22][3] + xor_out[81][22][3] + xor_out[82][22][3] + xor_out[83][22][3] + xor_out[84][22][3];
assign sum_out[17][22][3] = xor_out[85][22][3] + xor_out[86][22][3] + xor_out[87][22][3] + xor_out[88][22][3] + xor_out[89][22][3];
assign sum_out[18][22][3] = xor_out[90][22][3] + xor_out[91][22][3] + xor_out[92][22][3] + xor_out[93][22][3] + xor_out[94][22][3];
assign sum_out[19][22][3] = xor_out[95][22][3] + xor_out[96][22][3] + xor_out[97][22][3] + xor_out[98][22][3] + xor_out[99][22][3];

assign sum_out[0][22][4] = xor_out[0][22][4] + xor_out[1][22][4] + xor_out[2][22][4] + xor_out[3][22][4] + xor_out[4][22][4];
assign sum_out[1][22][4] = xor_out[5][22][4] + xor_out[6][22][4] + xor_out[7][22][4] + xor_out[8][22][4] + xor_out[9][22][4];
assign sum_out[2][22][4] = xor_out[10][22][4] + xor_out[11][22][4] + xor_out[12][22][4] + xor_out[13][22][4] + xor_out[14][22][4];
assign sum_out[3][22][4] = xor_out[15][22][4] + xor_out[16][22][4] + xor_out[17][22][4] + xor_out[18][22][4] + xor_out[19][22][4];
assign sum_out[4][22][4] = xor_out[20][22][4] + xor_out[21][22][4] + xor_out[22][22][4] + xor_out[23][22][4] + xor_out[24][22][4];
assign sum_out[5][22][4] = xor_out[25][22][4] + xor_out[26][22][4] + xor_out[27][22][4] + xor_out[28][22][4] + xor_out[29][22][4];
assign sum_out[6][22][4] = xor_out[30][22][4] + xor_out[31][22][4] + xor_out[32][22][4] + xor_out[33][22][4] + xor_out[34][22][4];
assign sum_out[7][22][4] = xor_out[35][22][4] + xor_out[36][22][4] + xor_out[37][22][4] + xor_out[38][22][4] + xor_out[39][22][4];
assign sum_out[8][22][4] = xor_out[40][22][4] + xor_out[41][22][4] + xor_out[42][22][4] + xor_out[43][22][4] + xor_out[44][22][4];
assign sum_out[9][22][4] = xor_out[45][22][4] + xor_out[46][22][4] + xor_out[47][22][4] + xor_out[48][22][4] + xor_out[49][22][4];
assign sum_out[10][22][4] = xor_out[50][22][4] + xor_out[51][22][4] + xor_out[52][22][4] + xor_out[53][22][4] + xor_out[54][22][4];
assign sum_out[11][22][4] = xor_out[55][22][4] + xor_out[56][22][4] + xor_out[57][22][4] + xor_out[58][22][4] + xor_out[59][22][4];
assign sum_out[12][22][4] = xor_out[60][22][4] + xor_out[61][22][4] + xor_out[62][22][4] + xor_out[63][22][4] + xor_out[64][22][4];
assign sum_out[13][22][4] = xor_out[65][22][4] + xor_out[66][22][4] + xor_out[67][22][4] + xor_out[68][22][4] + xor_out[69][22][4];
assign sum_out[14][22][4] = xor_out[70][22][4] + xor_out[71][22][4] + xor_out[72][22][4] + xor_out[73][22][4] + xor_out[74][22][4];
assign sum_out[15][22][4] = xor_out[75][22][4] + xor_out[76][22][4] + xor_out[77][22][4] + xor_out[78][22][4] + xor_out[79][22][4];
assign sum_out[16][22][4] = xor_out[80][22][4] + xor_out[81][22][4] + xor_out[82][22][4] + xor_out[83][22][4] + xor_out[84][22][4];
assign sum_out[17][22][4] = xor_out[85][22][4] + xor_out[86][22][4] + xor_out[87][22][4] + xor_out[88][22][4] + xor_out[89][22][4];
assign sum_out[18][22][4] = xor_out[90][22][4] + xor_out[91][22][4] + xor_out[92][22][4] + xor_out[93][22][4] + xor_out[94][22][4];
assign sum_out[19][22][4] = xor_out[95][22][4] + xor_out[96][22][4] + xor_out[97][22][4] + xor_out[98][22][4] + xor_out[99][22][4];

assign sum_out[0][22][5] = xor_out[0][22][5] + xor_out[1][22][5] + xor_out[2][22][5] + xor_out[3][22][5] + xor_out[4][22][5];
assign sum_out[1][22][5] = xor_out[5][22][5] + xor_out[6][22][5] + xor_out[7][22][5] + xor_out[8][22][5] + xor_out[9][22][5];
assign sum_out[2][22][5] = xor_out[10][22][5] + xor_out[11][22][5] + xor_out[12][22][5] + xor_out[13][22][5] + xor_out[14][22][5];
assign sum_out[3][22][5] = xor_out[15][22][5] + xor_out[16][22][5] + xor_out[17][22][5] + xor_out[18][22][5] + xor_out[19][22][5];
assign sum_out[4][22][5] = xor_out[20][22][5] + xor_out[21][22][5] + xor_out[22][22][5] + xor_out[23][22][5] + xor_out[24][22][5];
assign sum_out[5][22][5] = xor_out[25][22][5] + xor_out[26][22][5] + xor_out[27][22][5] + xor_out[28][22][5] + xor_out[29][22][5];
assign sum_out[6][22][5] = xor_out[30][22][5] + xor_out[31][22][5] + xor_out[32][22][5] + xor_out[33][22][5] + xor_out[34][22][5];
assign sum_out[7][22][5] = xor_out[35][22][5] + xor_out[36][22][5] + xor_out[37][22][5] + xor_out[38][22][5] + xor_out[39][22][5];
assign sum_out[8][22][5] = xor_out[40][22][5] + xor_out[41][22][5] + xor_out[42][22][5] + xor_out[43][22][5] + xor_out[44][22][5];
assign sum_out[9][22][5] = xor_out[45][22][5] + xor_out[46][22][5] + xor_out[47][22][5] + xor_out[48][22][5] + xor_out[49][22][5];
assign sum_out[10][22][5] = xor_out[50][22][5] + xor_out[51][22][5] + xor_out[52][22][5] + xor_out[53][22][5] + xor_out[54][22][5];
assign sum_out[11][22][5] = xor_out[55][22][5] + xor_out[56][22][5] + xor_out[57][22][5] + xor_out[58][22][5] + xor_out[59][22][5];
assign sum_out[12][22][5] = xor_out[60][22][5] + xor_out[61][22][5] + xor_out[62][22][5] + xor_out[63][22][5] + xor_out[64][22][5];
assign sum_out[13][22][5] = xor_out[65][22][5] + xor_out[66][22][5] + xor_out[67][22][5] + xor_out[68][22][5] + xor_out[69][22][5];
assign sum_out[14][22][5] = xor_out[70][22][5] + xor_out[71][22][5] + xor_out[72][22][5] + xor_out[73][22][5] + xor_out[74][22][5];
assign sum_out[15][22][5] = xor_out[75][22][5] + xor_out[76][22][5] + xor_out[77][22][5] + xor_out[78][22][5] + xor_out[79][22][5];
assign sum_out[16][22][5] = xor_out[80][22][5] + xor_out[81][22][5] + xor_out[82][22][5] + xor_out[83][22][5] + xor_out[84][22][5];
assign sum_out[17][22][5] = xor_out[85][22][5] + xor_out[86][22][5] + xor_out[87][22][5] + xor_out[88][22][5] + xor_out[89][22][5];
assign sum_out[18][22][5] = xor_out[90][22][5] + xor_out[91][22][5] + xor_out[92][22][5] + xor_out[93][22][5] + xor_out[94][22][5];
assign sum_out[19][22][5] = xor_out[95][22][5] + xor_out[96][22][5] + xor_out[97][22][5] + xor_out[98][22][5] + xor_out[99][22][5];

assign sum_out[0][22][6] = xor_out[0][22][6] + xor_out[1][22][6] + xor_out[2][22][6] + xor_out[3][22][6] + xor_out[4][22][6];
assign sum_out[1][22][6] = xor_out[5][22][6] + xor_out[6][22][6] + xor_out[7][22][6] + xor_out[8][22][6] + xor_out[9][22][6];
assign sum_out[2][22][6] = xor_out[10][22][6] + xor_out[11][22][6] + xor_out[12][22][6] + xor_out[13][22][6] + xor_out[14][22][6];
assign sum_out[3][22][6] = xor_out[15][22][6] + xor_out[16][22][6] + xor_out[17][22][6] + xor_out[18][22][6] + xor_out[19][22][6];
assign sum_out[4][22][6] = xor_out[20][22][6] + xor_out[21][22][6] + xor_out[22][22][6] + xor_out[23][22][6] + xor_out[24][22][6];
assign sum_out[5][22][6] = xor_out[25][22][6] + xor_out[26][22][6] + xor_out[27][22][6] + xor_out[28][22][6] + xor_out[29][22][6];
assign sum_out[6][22][6] = xor_out[30][22][6] + xor_out[31][22][6] + xor_out[32][22][6] + xor_out[33][22][6] + xor_out[34][22][6];
assign sum_out[7][22][6] = xor_out[35][22][6] + xor_out[36][22][6] + xor_out[37][22][6] + xor_out[38][22][6] + xor_out[39][22][6];
assign sum_out[8][22][6] = xor_out[40][22][6] + xor_out[41][22][6] + xor_out[42][22][6] + xor_out[43][22][6] + xor_out[44][22][6];
assign sum_out[9][22][6] = xor_out[45][22][6] + xor_out[46][22][6] + xor_out[47][22][6] + xor_out[48][22][6] + xor_out[49][22][6];
assign sum_out[10][22][6] = xor_out[50][22][6] + xor_out[51][22][6] + xor_out[52][22][6] + xor_out[53][22][6] + xor_out[54][22][6];
assign sum_out[11][22][6] = xor_out[55][22][6] + xor_out[56][22][6] + xor_out[57][22][6] + xor_out[58][22][6] + xor_out[59][22][6];
assign sum_out[12][22][6] = xor_out[60][22][6] + xor_out[61][22][6] + xor_out[62][22][6] + xor_out[63][22][6] + xor_out[64][22][6];
assign sum_out[13][22][6] = xor_out[65][22][6] + xor_out[66][22][6] + xor_out[67][22][6] + xor_out[68][22][6] + xor_out[69][22][6];
assign sum_out[14][22][6] = xor_out[70][22][6] + xor_out[71][22][6] + xor_out[72][22][6] + xor_out[73][22][6] + xor_out[74][22][6];
assign sum_out[15][22][6] = xor_out[75][22][6] + xor_out[76][22][6] + xor_out[77][22][6] + xor_out[78][22][6] + xor_out[79][22][6];
assign sum_out[16][22][6] = xor_out[80][22][6] + xor_out[81][22][6] + xor_out[82][22][6] + xor_out[83][22][6] + xor_out[84][22][6];
assign sum_out[17][22][6] = xor_out[85][22][6] + xor_out[86][22][6] + xor_out[87][22][6] + xor_out[88][22][6] + xor_out[89][22][6];
assign sum_out[18][22][6] = xor_out[90][22][6] + xor_out[91][22][6] + xor_out[92][22][6] + xor_out[93][22][6] + xor_out[94][22][6];
assign sum_out[19][22][6] = xor_out[95][22][6] + xor_out[96][22][6] + xor_out[97][22][6] + xor_out[98][22][6] + xor_out[99][22][6];

assign sum_out[0][22][7] = xor_out[0][22][7] + xor_out[1][22][7] + xor_out[2][22][7] + xor_out[3][22][7] + xor_out[4][22][7];
assign sum_out[1][22][7] = xor_out[5][22][7] + xor_out[6][22][7] + xor_out[7][22][7] + xor_out[8][22][7] + xor_out[9][22][7];
assign sum_out[2][22][7] = xor_out[10][22][7] + xor_out[11][22][7] + xor_out[12][22][7] + xor_out[13][22][7] + xor_out[14][22][7];
assign sum_out[3][22][7] = xor_out[15][22][7] + xor_out[16][22][7] + xor_out[17][22][7] + xor_out[18][22][7] + xor_out[19][22][7];
assign sum_out[4][22][7] = xor_out[20][22][7] + xor_out[21][22][7] + xor_out[22][22][7] + xor_out[23][22][7] + xor_out[24][22][7];
assign sum_out[5][22][7] = xor_out[25][22][7] + xor_out[26][22][7] + xor_out[27][22][7] + xor_out[28][22][7] + xor_out[29][22][7];
assign sum_out[6][22][7] = xor_out[30][22][7] + xor_out[31][22][7] + xor_out[32][22][7] + xor_out[33][22][7] + xor_out[34][22][7];
assign sum_out[7][22][7] = xor_out[35][22][7] + xor_out[36][22][7] + xor_out[37][22][7] + xor_out[38][22][7] + xor_out[39][22][7];
assign sum_out[8][22][7] = xor_out[40][22][7] + xor_out[41][22][7] + xor_out[42][22][7] + xor_out[43][22][7] + xor_out[44][22][7];
assign sum_out[9][22][7] = xor_out[45][22][7] + xor_out[46][22][7] + xor_out[47][22][7] + xor_out[48][22][7] + xor_out[49][22][7];
assign sum_out[10][22][7] = xor_out[50][22][7] + xor_out[51][22][7] + xor_out[52][22][7] + xor_out[53][22][7] + xor_out[54][22][7];
assign sum_out[11][22][7] = xor_out[55][22][7] + xor_out[56][22][7] + xor_out[57][22][7] + xor_out[58][22][7] + xor_out[59][22][7];
assign sum_out[12][22][7] = xor_out[60][22][7] + xor_out[61][22][7] + xor_out[62][22][7] + xor_out[63][22][7] + xor_out[64][22][7];
assign sum_out[13][22][7] = xor_out[65][22][7] + xor_out[66][22][7] + xor_out[67][22][7] + xor_out[68][22][7] + xor_out[69][22][7];
assign sum_out[14][22][7] = xor_out[70][22][7] + xor_out[71][22][7] + xor_out[72][22][7] + xor_out[73][22][7] + xor_out[74][22][7];
assign sum_out[15][22][7] = xor_out[75][22][7] + xor_out[76][22][7] + xor_out[77][22][7] + xor_out[78][22][7] + xor_out[79][22][7];
assign sum_out[16][22][7] = xor_out[80][22][7] + xor_out[81][22][7] + xor_out[82][22][7] + xor_out[83][22][7] + xor_out[84][22][7];
assign sum_out[17][22][7] = xor_out[85][22][7] + xor_out[86][22][7] + xor_out[87][22][7] + xor_out[88][22][7] + xor_out[89][22][7];
assign sum_out[18][22][7] = xor_out[90][22][7] + xor_out[91][22][7] + xor_out[92][22][7] + xor_out[93][22][7] + xor_out[94][22][7];
assign sum_out[19][22][7] = xor_out[95][22][7] + xor_out[96][22][7] + xor_out[97][22][7] + xor_out[98][22][7] + xor_out[99][22][7];

assign sum_out[0][22][8] = xor_out[0][22][8] + xor_out[1][22][8] + xor_out[2][22][8] + xor_out[3][22][8] + xor_out[4][22][8];
assign sum_out[1][22][8] = xor_out[5][22][8] + xor_out[6][22][8] + xor_out[7][22][8] + xor_out[8][22][8] + xor_out[9][22][8];
assign sum_out[2][22][8] = xor_out[10][22][8] + xor_out[11][22][8] + xor_out[12][22][8] + xor_out[13][22][8] + xor_out[14][22][8];
assign sum_out[3][22][8] = xor_out[15][22][8] + xor_out[16][22][8] + xor_out[17][22][8] + xor_out[18][22][8] + xor_out[19][22][8];
assign sum_out[4][22][8] = xor_out[20][22][8] + xor_out[21][22][8] + xor_out[22][22][8] + xor_out[23][22][8] + xor_out[24][22][8];
assign sum_out[5][22][8] = xor_out[25][22][8] + xor_out[26][22][8] + xor_out[27][22][8] + xor_out[28][22][8] + xor_out[29][22][8];
assign sum_out[6][22][8] = xor_out[30][22][8] + xor_out[31][22][8] + xor_out[32][22][8] + xor_out[33][22][8] + xor_out[34][22][8];
assign sum_out[7][22][8] = xor_out[35][22][8] + xor_out[36][22][8] + xor_out[37][22][8] + xor_out[38][22][8] + xor_out[39][22][8];
assign sum_out[8][22][8] = xor_out[40][22][8] + xor_out[41][22][8] + xor_out[42][22][8] + xor_out[43][22][8] + xor_out[44][22][8];
assign sum_out[9][22][8] = xor_out[45][22][8] + xor_out[46][22][8] + xor_out[47][22][8] + xor_out[48][22][8] + xor_out[49][22][8];
assign sum_out[10][22][8] = xor_out[50][22][8] + xor_out[51][22][8] + xor_out[52][22][8] + xor_out[53][22][8] + xor_out[54][22][8];
assign sum_out[11][22][8] = xor_out[55][22][8] + xor_out[56][22][8] + xor_out[57][22][8] + xor_out[58][22][8] + xor_out[59][22][8];
assign sum_out[12][22][8] = xor_out[60][22][8] + xor_out[61][22][8] + xor_out[62][22][8] + xor_out[63][22][8] + xor_out[64][22][8];
assign sum_out[13][22][8] = xor_out[65][22][8] + xor_out[66][22][8] + xor_out[67][22][8] + xor_out[68][22][8] + xor_out[69][22][8];
assign sum_out[14][22][8] = xor_out[70][22][8] + xor_out[71][22][8] + xor_out[72][22][8] + xor_out[73][22][8] + xor_out[74][22][8];
assign sum_out[15][22][8] = xor_out[75][22][8] + xor_out[76][22][8] + xor_out[77][22][8] + xor_out[78][22][8] + xor_out[79][22][8];
assign sum_out[16][22][8] = xor_out[80][22][8] + xor_out[81][22][8] + xor_out[82][22][8] + xor_out[83][22][8] + xor_out[84][22][8];
assign sum_out[17][22][8] = xor_out[85][22][8] + xor_out[86][22][8] + xor_out[87][22][8] + xor_out[88][22][8] + xor_out[89][22][8];
assign sum_out[18][22][8] = xor_out[90][22][8] + xor_out[91][22][8] + xor_out[92][22][8] + xor_out[93][22][8] + xor_out[94][22][8];
assign sum_out[19][22][8] = xor_out[95][22][8] + xor_out[96][22][8] + xor_out[97][22][8] + xor_out[98][22][8] + xor_out[99][22][8];

assign sum_out[0][22][9] = xor_out[0][22][9] + xor_out[1][22][9] + xor_out[2][22][9] + xor_out[3][22][9] + xor_out[4][22][9];
assign sum_out[1][22][9] = xor_out[5][22][9] + xor_out[6][22][9] + xor_out[7][22][9] + xor_out[8][22][9] + xor_out[9][22][9];
assign sum_out[2][22][9] = xor_out[10][22][9] + xor_out[11][22][9] + xor_out[12][22][9] + xor_out[13][22][9] + xor_out[14][22][9];
assign sum_out[3][22][9] = xor_out[15][22][9] + xor_out[16][22][9] + xor_out[17][22][9] + xor_out[18][22][9] + xor_out[19][22][9];
assign sum_out[4][22][9] = xor_out[20][22][9] + xor_out[21][22][9] + xor_out[22][22][9] + xor_out[23][22][9] + xor_out[24][22][9];
assign sum_out[5][22][9] = xor_out[25][22][9] + xor_out[26][22][9] + xor_out[27][22][9] + xor_out[28][22][9] + xor_out[29][22][9];
assign sum_out[6][22][9] = xor_out[30][22][9] + xor_out[31][22][9] + xor_out[32][22][9] + xor_out[33][22][9] + xor_out[34][22][9];
assign sum_out[7][22][9] = xor_out[35][22][9] + xor_out[36][22][9] + xor_out[37][22][9] + xor_out[38][22][9] + xor_out[39][22][9];
assign sum_out[8][22][9] = xor_out[40][22][9] + xor_out[41][22][9] + xor_out[42][22][9] + xor_out[43][22][9] + xor_out[44][22][9];
assign sum_out[9][22][9] = xor_out[45][22][9] + xor_out[46][22][9] + xor_out[47][22][9] + xor_out[48][22][9] + xor_out[49][22][9];
assign sum_out[10][22][9] = xor_out[50][22][9] + xor_out[51][22][9] + xor_out[52][22][9] + xor_out[53][22][9] + xor_out[54][22][9];
assign sum_out[11][22][9] = xor_out[55][22][9] + xor_out[56][22][9] + xor_out[57][22][9] + xor_out[58][22][9] + xor_out[59][22][9];
assign sum_out[12][22][9] = xor_out[60][22][9] + xor_out[61][22][9] + xor_out[62][22][9] + xor_out[63][22][9] + xor_out[64][22][9];
assign sum_out[13][22][9] = xor_out[65][22][9] + xor_out[66][22][9] + xor_out[67][22][9] + xor_out[68][22][9] + xor_out[69][22][9];
assign sum_out[14][22][9] = xor_out[70][22][9] + xor_out[71][22][9] + xor_out[72][22][9] + xor_out[73][22][9] + xor_out[74][22][9];
assign sum_out[15][22][9] = xor_out[75][22][9] + xor_out[76][22][9] + xor_out[77][22][9] + xor_out[78][22][9] + xor_out[79][22][9];
assign sum_out[16][22][9] = xor_out[80][22][9] + xor_out[81][22][9] + xor_out[82][22][9] + xor_out[83][22][9] + xor_out[84][22][9];
assign sum_out[17][22][9] = xor_out[85][22][9] + xor_out[86][22][9] + xor_out[87][22][9] + xor_out[88][22][9] + xor_out[89][22][9];
assign sum_out[18][22][9] = xor_out[90][22][9] + xor_out[91][22][9] + xor_out[92][22][9] + xor_out[93][22][9] + xor_out[94][22][9];
assign sum_out[19][22][9] = xor_out[95][22][9] + xor_out[96][22][9] + xor_out[97][22][9] + xor_out[98][22][9] + xor_out[99][22][9];

assign sum_out[0][22][10] = xor_out[0][22][10] + xor_out[1][22][10] + xor_out[2][22][10] + xor_out[3][22][10] + xor_out[4][22][10];
assign sum_out[1][22][10] = xor_out[5][22][10] + xor_out[6][22][10] + xor_out[7][22][10] + xor_out[8][22][10] + xor_out[9][22][10];
assign sum_out[2][22][10] = xor_out[10][22][10] + xor_out[11][22][10] + xor_out[12][22][10] + xor_out[13][22][10] + xor_out[14][22][10];
assign sum_out[3][22][10] = xor_out[15][22][10] + xor_out[16][22][10] + xor_out[17][22][10] + xor_out[18][22][10] + xor_out[19][22][10];
assign sum_out[4][22][10] = xor_out[20][22][10] + xor_out[21][22][10] + xor_out[22][22][10] + xor_out[23][22][10] + xor_out[24][22][10];
assign sum_out[5][22][10] = xor_out[25][22][10] + xor_out[26][22][10] + xor_out[27][22][10] + xor_out[28][22][10] + xor_out[29][22][10];
assign sum_out[6][22][10] = xor_out[30][22][10] + xor_out[31][22][10] + xor_out[32][22][10] + xor_out[33][22][10] + xor_out[34][22][10];
assign sum_out[7][22][10] = xor_out[35][22][10] + xor_out[36][22][10] + xor_out[37][22][10] + xor_out[38][22][10] + xor_out[39][22][10];
assign sum_out[8][22][10] = xor_out[40][22][10] + xor_out[41][22][10] + xor_out[42][22][10] + xor_out[43][22][10] + xor_out[44][22][10];
assign sum_out[9][22][10] = xor_out[45][22][10] + xor_out[46][22][10] + xor_out[47][22][10] + xor_out[48][22][10] + xor_out[49][22][10];
assign sum_out[10][22][10] = xor_out[50][22][10] + xor_out[51][22][10] + xor_out[52][22][10] + xor_out[53][22][10] + xor_out[54][22][10];
assign sum_out[11][22][10] = xor_out[55][22][10] + xor_out[56][22][10] + xor_out[57][22][10] + xor_out[58][22][10] + xor_out[59][22][10];
assign sum_out[12][22][10] = xor_out[60][22][10] + xor_out[61][22][10] + xor_out[62][22][10] + xor_out[63][22][10] + xor_out[64][22][10];
assign sum_out[13][22][10] = xor_out[65][22][10] + xor_out[66][22][10] + xor_out[67][22][10] + xor_out[68][22][10] + xor_out[69][22][10];
assign sum_out[14][22][10] = xor_out[70][22][10] + xor_out[71][22][10] + xor_out[72][22][10] + xor_out[73][22][10] + xor_out[74][22][10];
assign sum_out[15][22][10] = xor_out[75][22][10] + xor_out[76][22][10] + xor_out[77][22][10] + xor_out[78][22][10] + xor_out[79][22][10];
assign sum_out[16][22][10] = xor_out[80][22][10] + xor_out[81][22][10] + xor_out[82][22][10] + xor_out[83][22][10] + xor_out[84][22][10];
assign sum_out[17][22][10] = xor_out[85][22][10] + xor_out[86][22][10] + xor_out[87][22][10] + xor_out[88][22][10] + xor_out[89][22][10];
assign sum_out[18][22][10] = xor_out[90][22][10] + xor_out[91][22][10] + xor_out[92][22][10] + xor_out[93][22][10] + xor_out[94][22][10];
assign sum_out[19][22][10] = xor_out[95][22][10] + xor_out[96][22][10] + xor_out[97][22][10] + xor_out[98][22][10] + xor_out[99][22][10];

assign sum_out[0][22][11] = xor_out[0][22][11] + xor_out[1][22][11] + xor_out[2][22][11] + xor_out[3][22][11] + xor_out[4][22][11];
assign sum_out[1][22][11] = xor_out[5][22][11] + xor_out[6][22][11] + xor_out[7][22][11] + xor_out[8][22][11] + xor_out[9][22][11];
assign sum_out[2][22][11] = xor_out[10][22][11] + xor_out[11][22][11] + xor_out[12][22][11] + xor_out[13][22][11] + xor_out[14][22][11];
assign sum_out[3][22][11] = xor_out[15][22][11] + xor_out[16][22][11] + xor_out[17][22][11] + xor_out[18][22][11] + xor_out[19][22][11];
assign sum_out[4][22][11] = xor_out[20][22][11] + xor_out[21][22][11] + xor_out[22][22][11] + xor_out[23][22][11] + xor_out[24][22][11];
assign sum_out[5][22][11] = xor_out[25][22][11] + xor_out[26][22][11] + xor_out[27][22][11] + xor_out[28][22][11] + xor_out[29][22][11];
assign sum_out[6][22][11] = xor_out[30][22][11] + xor_out[31][22][11] + xor_out[32][22][11] + xor_out[33][22][11] + xor_out[34][22][11];
assign sum_out[7][22][11] = xor_out[35][22][11] + xor_out[36][22][11] + xor_out[37][22][11] + xor_out[38][22][11] + xor_out[39][22][11];
assign sum_out[8][22][11] = xor_out[40][22][11] + xor_out[41][22][11] + xor_out[42][22][11] + xor_out[43][22][11] + xor_out[44][22][11];
assign sum_out[9][22][11] = xor_out[45][22][11] + xor_out[46][22][11] + xor_out[47][22][11] + xor_out[48][22][11] + xor_out[49][22][11];
assign sum_out[10][22][11] = xor_out[50][22][11] + xor_out[51][22][11] + xor_out[52][22][11] + xor_out[53][22][11] + xor_out[54][22][11];
assign sum_out[11][22][11] = xor_out[55][22][11] + xor_out[56][22][11] + xor_out[57][22][11] + xor_out[58][22][11] + xor_out[59][22][11];
assign sum_out[12][22][11] = xor_out[60][22][11] + xor_out[61][22][11] + xor_out[62][22][11] + xor_out[63][22][11] + xor_out[64][22][11];
assign sum_out[13][22][11] = xor_out[65][22][11] + xor_out[66][22][11] + xor_out[67][22][11] + xor_out[68][22][11] + xor_out[69][22][11];
assign sum_out[14][22][11] = xor_out[70][22][11] + xor_out[71][22][11] + xor_out[72][22][11] + xor_out[73][22][11] + xor_out[74][22][11];
assign sum_out[15][22][11] = xor_out[75][22][11] + xor_out[76][22][11] + xor_out[77][22][11] + xor_out[78][22][11] + xor_out[79][22][11];
assign sum_out[16][22][11] = xor_out[80][22][11] + xor_out[81][22][11] + xor_out[82][22][11] + xor_out[83][22][11] + xor_out[84][22][11];
assign sum_out[17][22][11] = xor_out[85][22][11] + xor_out[86][22][11] + xor_out[87][22][11] + xor_out[88][22][11] + xor_out[89][22][11];
assign sum_out[18][22][11] = xor_out[90][22][11] + xor_out[91][22][11] + xor_out[92][22][11] + xor_out[93][22][11] + xor_out[94][22][11];
assign sum_out[19][22][11] = xor_out[95][22][11] + xor_out[96][22][11] + xor_out[97][22][11] + xor_out[98][22][11] + xor_out[99][22][11];

assign sum_out[0][22][12] = xor_out[0][22][12] + xor_out[1][22][12] + xor_out[2][22][12] + xor_out[3][22][12] + xor_out[4][22][12];
assign sum_out[1][22][12] = xor_out[5][22][12] + xor_out[6][22][12] + xor_out[7][22][12] + xor_out[8][22][12] + xor_out[9][22][12];
assign sum_out[2][22][12] = xor_out[10][22][12] + xor_out[11][22][12] + xor_out[12][22][12] + xor_out[13][22][12] + xor_out[14][22][12];
assign sum_out[3][22][12] = xor_out[15][22][12] + xor_out[16][22][12] + xor_out[17][22][12] + xor_out[18][22][12] + xor_out[19][22][12];
assign sum_out[4][22][12] = xor_out[20][22][12] + xor_out[21][22][12] + xor_out[22][22][12] + xor_out[23][22][12] + xor_out[24][22][12];
assign sum_out[5][22][12] = xor_out[25][22][12] + xor_out[26][22][12] + xor_out[27][22][12] + xor_out[28][22][12] + xor_out[29][22][12];
assign sum_out[6][22][12] = xor_out[30][22][12] + xor_out[31][22][12] + xor_out[32][22][12] + xor_out[33][22][12] + xor_out[34][22][12];
assign sum_out[7][22][12] = xor_out[35][22][12] + xor_out[36][22][12] + xor_out[37][22][12] + xor_out[38][22][12] + xor_out[39][22][12];
assign sum_out[8][22][12] = xor_out[40][22][12] + xor_out[41][22][12] + xor_out[42][22][12] + xor_out[43][22][12] + xor_out[44][22][12];
assign sum_out[9][22][12] = xor_out[45][22][12] + xor_out[46][22][12] + xor_out[47][22][12] + xor_out[48][22][12] + xor_out[49][22][12];
assign sum_out[10][22][12] = xor_out[50][22][12] + xor_out[51][22][12] + xor_out[52][22][12] + xor_out[53][22][12] + xor_out[54][22][12];
assign sum_out[11][22][12] = xor_out[55][22][12] + xor_out[56][22][12] + xor_out[57][22][12] + xor_out[58][22][12] + xor_out[59][22][12];
assign sum_out[12][22][12] = xor_out[60][22][12] + xor_out[61][22][12] + xor_out[62][22][12] + xor_out[63][22][12] + xor_out[64][22][12];
assign sum_out[13][22][12] = xor_out[65][22][12] + xor_out[66][22][12] + xor_out[67][22][12] + xor_out[68][22][12] + xor_out[69][22][12];
assign sum_out[14][22][12] = xor_out[70][22][12] + xor_out[71][22][12] + xor_out[72][22][12] + xor_out[73][22][12] + xor_out[74][22][12];
assign sum_out[15][22][12] = xor_out[75][22][12] + xor_out[76][22][12] + xor_out[77][22][12] + xor_out[78][22][12] + xor_out[79][22][12];
assign sum_out[16][22][12] = xor_out[80][22][12] + xor_out[81][22][12] + xor_out[82][22][12] + xor_out[83][22][12] + xor_out[84][22][12];
assign sum_out[17][22][12] = xor_out[85][22][12] + xor_out[86][22][12] + xor_out[87][22][12] + xor_out[88][22][12] + xor_out[89][22][12];
assign sum_out[18][22][12] = xor_out[90][22][12] + xor_out[91][22][12] + xor_out[92][22][12] + xor_out[93][22][12] + xor_out[94][22][12];
assign sum_out[19][22][12] = xor_out[95][22][12] + xor_out[96][22][12] + xor_out[97][22][12] + xor_out[98][22][12] + xor_out[99][22][12];

assign sum_out[0][22][13] = xor_out[0][22][13] + xor_out[1][22][13] + xor_out[2][22][13] + xor_out[3][22][13] + xor_out[4][22][13];
assign sum_out[1][22][13] = xor_out[5][22][13] + xor_out[6][22][13] + xor_out[7][22][13] + xor_out[8][22][13] + xor_out[9][22][13];
assign sum_out[2][22][13] = xor_out[10][22][13] + xor_out[11][22][13] + xor_out[12][22][13] + xor_out[13][22][13] + xor_out[14][22][13];
assign sum_out[3][22][13] = xor_out[15][22][13] + xor_out[16][22][13] + xor_out[17][22][13] + xor_out[18][22][13] + xor_out[19][22][13];
assign sum_out[4][22][13] = xor_out[20][22][13] + xor_out[21][22][13] + xor_out[22][22][13] + xor_out[23][22][13] + xor_out[24][22][13];
assign sum_out[5][22][13] = xor_out[25][22][13] + xor_out[26][22][13] + xor_out[27][22][13] + xor_out[28][22][13] + xor_out[29][22][13];
assign sum_out[6][22][13] = xor_out[30][22][13] + xor_out[31][22][13] + xor_out[32][22][13] + xor_out[33][22][13] + xor_out[34][22][13];
assign sum_out[7][22][13] = xor_out[35][22][13] + xor_out[36][22][13] + xor_out[37][22][13] + xor_out[38][22][13] + xor_out[39][22][13];
assign sum_out[8][22][13] = xor_out[40][22][13] + xor_out[41][22][13] + xor_out[42][22][13] + xor_out[43][22][13] + xor_out[44][22][13];
assign sum_out[9][22][13] = xor_out[45][22][13] + xor_out[46][22][13] + xor_out[47][22][13] + xor_out[48][22][13] + xor_out[49][22][13];
assign sum_out[10][22][13] = xor_out[50][22][13] + xor_out[51][22][13] + xor_out[52][22][13] + xor_out[53][22][13] + xor_out[54][22][13];
assign sum_out[11][22][13] = xor_out[55][22][13] + xor_out[56][22][13] + xor_out[57][22][13] + xor_out[58][22][13] + xor_out[59][22][13];
assign sum_out[12][22][13] = xor_out[60][22][13] + xor_out[61][22][13] + xor_out[62][22][13] + xor_out[63][22][13] + xor_out[64][22][13];
assign sum_out[13][22][13] = xor_out[65][22][13] + xor_out[66][22][13] + xor_out[67][22][13] + xor_out[68][22][13] + xor_out[69][22][13];
assign sum_out[14][22][13] = xor_out[70][22][13] + xor_out[71][22][13] + xor_out[72][22][13] + xor_out[73][22][13] + xor_out[74][22][13];
assign sum_out[15][22][13] = xor_out[75][22][13] + xor_out[76][22][13] + xor_out[77][22][13] + xor_out[78][22][13] + xor_out[79][22][13];
assign sum_out[16][22][13] = xor_out[80][22][13] + xor_out[81][22][13] + xor_out[82][22][13] + xor_out[83][22][13] + xor_out[84][22][13];
assign sum_out[17][22][13] = xor_out[85][22][13] + xor_out[86][22][13] + xor_out[87][22][13] + xor_out[88][22][13] + xor_out[89][22][13];
assign sum_out[18][22][13] = xor_out[90][22][13] + xor_out[91][22][13] + xor_out[92][22][13] + xor_out[93][22][13] + xor_out[94][22][13];
assign sum_out[19][22][13] = xor_out[95][22][13] + xor_out[96][22][13] + xor_out[97][22][13] + xor_out[98][22][13] + xor_out[99][22][13];

assign sum_out[0][22][14] = xor_out[0][22][14] + xor_out[1][22][14] + xor_out[2][22][14] + xor_out[3][22][14] + xor_out[4][22][14];
assign sum_out[1][22][14] = xor_out[5][22][14] + xor_out[6][22][14] + xor_out[7][22][14] + xor_out[8][22][14] + xor_out[9][22][14];
assign sum_out[2][22][14] = xor_out[10][22][14] + xor_out[11][22][14] + xor_out[12][22][14] + xor_out[13][22][14] + xor_out[14][22][14];
assign sum_out[3][22][14] = xor_out[15][22][14] + xor_out[16][22][14] + xor_out[17][22][14] + xor_out[18][22][14] + xor_out[19][22][14];
assign sum_out[4][22][14] = xor_out[20][22][14] + xor_out[21][22][14] + xor_out[22][22][14] + xor_out[23][22][14] + xor_out[24][22][14];
assign sum_out[5][22][14] = xor_out[25][22][14] + xor_out[26][22][14] + xor_out[27][22][14] + xor_out[28][22][14] + xor_out[29][22][14];
assign sum_out[6][22][14] = xor_out[30][22][14] + xor_out[31][22][14] + xor_out[32][22][14] + xor_out[33][22][14] + xor_out[34][22][14];
assign sum_out[7][22][14] = xor_out[35][22][14] + xor_out[36][22][14] + xor_out[37][22][14] + xor_out[38][22][14] + xor_out[39][22][14];
assign sum_out[8][22][14] = xor_out[40][22][14] + xor_out[41][22][14] + xor_out[42][22][14] + xor_out[43][22][14] + xor_out[44][22][14];
assign sum_out[9][22][14] = xor_out[45][22][14] + xor_out[46][22][14] + xor_out[47][22][14] + xor_out[48][22][14] + xor_out[49][22][14];
assign sum_out[10][22][14] = xor_out[50][22][14] + xor_out[51][22][14] + xor_out[52][22][14] + xor_out[53][22][14] + xor_out[54][22][14];
assign sum_out[11][22][14] = xor_out[55][22][14] + xor_out[56][22][14] + xor_out[57][22][14] + xor_out[58][22][14] + xor_out[59][22][14];
assign sum_out[12][22][14] = xor_out[60][22][14] + xor_out[61][22][14] + xor_out[62][22][14] + xor_out[63][22][14] + xor_out[64][22][14];
assign sum_out[13][22][14] = xor_out[65][22][14] + xor_out[66][22][14] + xor_out[67][22][14] + xor_out[68][22][14] + xor_out[69][22][14];
assign sum_out[14][22][14] = xor_out[70][22][14] + xor_out[71][22][14] + xor_out[72][22][14] + xor_out[73][22][14] + xor_out[74][22][14];
assign sum_out[15][22][14] = xor_out[75][22][14] + xor_out[76][22][14] + xor_out[77][22][14] + xor_out[78][22][14] + xor_out[79][22][14];
assign sum_out[16][22][14] = xor_out[80][22][14] + xor_out[81][22][14] + xor_out[82][22][14] + xor_out[83][22][14] + xor_out[84][22][14];
assign sum_out[17][22][14] = xor_out[85][22][14] + xor_out[86][22][14] + xor_out[87][22][14] + xor_out[88][22][14] + xor_out[89][22][14];
assign sum_out[18][22][14] = xor_out[90][22][14] + xor_out[91][22][14] + xor_out[92][22][14] + xor_out[93][22][14] + xor_out[94][22][14];
assign sum_out[19][22][14] = xor_out[95][22][14] + xor_out[96][22][14] + xor_out[97][22][14] + xor_out[98][22][14] + xor_out[99][22][14];

assign sum_out[0][22][15] = xor_out[0][22][15] + xor_out[1][22][15] + xor_out[2][22][15] + xor_out[3][22][15] + xor_out[4][22][15];
assign sum_out[1][22][15] = xor_out[5][22][15] + xor_out[6][22][15] + xor_out[7][22][15] + xor_out[8][22][15] + xor_out[9][22][15];
assign sum_out[2][22][15] = xor_out[10][22][15] + xor_out[11][22][15] + xor_out[12][22][15] + xor_out[13][22][15] + xor_out[14][22][15];
assign sum_out[3][22][15] = xor_out[15][22][15] + xor_out[16][22][15] + xor_out[17][22][15] + xor_out[18][22][15] + xor_out[19][22][15];
assign sum_out[4][22][15] = xor_out[20][22][15] + xor_out[21][22][15] + xor_out[22][22][15] + xor_out[23][22][15] + xor_out[24][22][15];
assign sum_out[5][22][15] = xor_out[25][22][15] + xor_out[26][22][15] + xor_out[27][22][15] + xor_out[28][22][15] + xor_out[29][22][15];
assign sum_out[6][22][15] = xor_out[30][22][15] + xor_out[31][22][15] + xor_out[32][22][15] + xor_out[33][22][15] + xor_out[34][22][15];
assign sum_out[7][22][15] = xor_out[35][22][15] + xor_out[36][22][15] + xor_out[37][22][15] + xor_out[38][22][15] + xor_out[39][22][15];
assign sum_out[8][22][15] = xor_out[40][22][15] + xor_out[41][22][15] + xor_out[42][22][15] + xor_out[43][22][15] + xor_out[44][22][15];
assign sum_out[9][22][15] = xor_out[45][22][15] + xor_out[46][22][15] + xor_out[47][22][15] + xor_out[48][22][15] + xor_out[49][22][15];
assign sum_out[10][22][15] = xor_out[50][22][15] + xor_out[51][22][15] + xor_out[52][22][15] + xor_out[53][22][15] + xor_out[54][22][15];
assign sum_out[11][22][15] = xor_out[55][22][15] + xor_out[56][22][15] + xor_out[57][22][15] + xor_out[58][22][15] + xor_out[59][22][15];
assign sum_out[12][22][15] = xor_out[60][22][15] + xor_out[61][22][15] + xor_out[62][22][15] + xor_out[63][22][15] + xor_out[64][22][15];
assign sum_out[13][22][15] = xor_out[65][22][15] + xor_out[66][22][15] + xor_out[67][22][15] + xor_out[68][22][15] + xor_out[69][22][15];
assign sum_out[14][22][15] = xor_out[70][22][15] + xor_out[71][22][15] + xor_out[72][22][15] + xor_out[73][22][15] + xor_out[74][22][15];
assign sum_out[15][22][15] = xor_out[75][22][15] + xor_out[76][22][15] + xor_out[77][22][15] + xor_out[78][22][15] + xor_out[79][22][15];
assign sum_out[16][22][15] = xor_out[80][22][15] + xor_out[81][22][15] + xor_out[82][22][15] + xor_out[83][22][15] + xor_out[84][22][15];
assign sum_out[17][22][15] = xor_out[85][22][15] + xor_out[86][22][15] + xor_out[87][22][15] + xor_out[88][22][15] + xor_out[89][22][15];
assign sum_out[18][22][15] = xor_out[90][22][15] + xor_out[91][22][15] + xor_out[92][22][15] + xor_out[93][22][15] + xor_out[94][22][15];
assign sum_out[19][22][15] = xor_out[95][22][15] + xor_out[96][22][15] + xor_out[97][22][15] + xor_out[98][22][15] + xor_out[99][22][15];

assign sum_out[0][22][16] = xor_out[0][22][16] + xor_out[1][22][16] + xor_out[2][22][16] + xor_out[3][22][16] + xor_out[4][22][16];
assign sum_out[1][22][16] = xor_out[5][22][16] + xor_out[6][22][16] + xor_out[7][22][16] + xor_out[8][22][16] + xor_out[9][22][16];
assign sum_out[2][22][16] = xor_out[10][22][16] + xor_out[11][22][16] + xor_out[12][22][16] + xor_out[13][22][16] + xor_out[14][22][16];
assign sum_out[3][22][16] = xor_out[15][22][16] + xor_out[16][22][16] + xor_out[17][22][16] + xor_out[18][22][16] + xor_out[19][22][16];
assign sum_out[4][22][16] = xor_out[20][22][16] + xor_out[21][22][16] + xor_out[22][22][16] + xor_out[23][22][16] + xor_out[24][22][16];
assign sum_out[5][22][16] = xor_out[25][22][16] + xor_out[26][22][16] + xor_out[27][22][16] + xor_out[28][22][16] + xor_out[29][22][16];
assign sum_out[6][22][16] = xor_out[30][22][16] + xor_out[31][22][16] + xor_out[32][22][16] + xor_out[33][22][16] + xor_out[34][22][16];
assign sum_out[7][22][16] = xor_out[35][22][16] + xor_out[36][22][16] + xor_out[37][22][16] + xor_out[38][22][16] + xor_out[39][22][16];
assign sum_out[8][22][16] = xor_out[40][22][16] + xor_out[41][22][16] + xor_out[42][22][16] + xor_out[43][22][16] + xor_out[44][22][16];
assign sum_out[9][22][16] = xor_out[45][22][16] + xor_out[46][22][16] + xor_out[47][22][16] + xor_out[48][22][16] + xor_out[49][22][16];
assign sum_out[10][22][16] = xor_out[50][22][16] + xor_out[51][22][16] + xor_out[52][22][16] + xor_out[53][22][16] + xor_out[54][22][16];
assign sum_out[11][22][16] = xor_out[55][22][16] + xor_out[56][22][16] + xor_out[57][22][16] + xor_out[58][22][16] + xor_out[59][22][16];
assign sum_out[12][22][16] = xor_out[60][22][16] + xor_out[61][22][16] + xor_out[62][22][16] + xor_out[63][22][16] + xor_out[64][22][16];
assign sum_out[13][22][16] = xor_out[65][22][16] + xor_out[66][22][16] + xor_out[67][22][16] + xor_out[68][22][16] + xor_out[69][22][16];
assign sum_out[14][22][16] = xor_out[70][22][16] + xor_out[71][22][16] + xor_out[72][22][16] + xor_out[73][22][16] + xor_out[74][22][16];
assign sum_out[15][22][16] = xor_out[75][22][16] + xor_out[76][22][16] + xor_out[77][22][16] + xor_out[78][22][16] + xor_out[79][22][16];
assign sum_out[16][22][16] = xor_out[80][22][16] + xor_out[81][22][16] + xor_out[82][22][16] + xor_out[83][22][16] + xor_out[84][22][16];
assign sum_out[17][22][16] = xor_out[85][22][16] + xor_out[86][22][16] + xor_out[87][22][16] + xor_out[88][22][16] + xor_out[89][22][16];
assign sum_out[18][22][16] = xor_out[90][22][16] + xor_out[91][22][16] + xor_out[92][22][16] + xor_out[93][22][16] + xor_out[94][22][16];
assign sum_out[19][22][16] = xor_out[95][22][16] + xor_out[96][22][16] + xor_out[97][22][16] + xor_out[98][22][16] + xor_out[99][22][16];

assign sum_out[0][22][17] = xor_out[0][22][17] + xor_out[1][22][17] + xor_out[2][22][17] + xor_out[3][22][17] + xor_out[4][22][17];
assign sum_out[1][22][17] = xor_out[5][22][17] + xor_out[6][22][17] + xor_out[7][22][17] + xor_out[8][22][17] + xor_out[9][22][17];
assign sum_out[2][22][17] = xor_out[10][22][17] + xor_out[11][22][17] + xor_out[12][22][17] + xor_out[13][22][17] + xor_out[14][22][17];
assign sum_out[3][22][17] = xor_out[15][22][17] + xor_out[16][22][17] + xor_out[17][22][17] + xor_out[18][22][17] + xor_out[19][22][17];
assign sum_out[4][22][17] = xor_out[20][22][17] + xor_out[21][22][17] + xor_out[22][22][17] + xor_out[23][22][17] + xor_out[24][22][17];
assign sum_out[5][22][17] = xor_out[25][22][17] + xor_out[26][22][17] + xor_out[27][22][17] + xor_out[28][22][17] + xor_out[29][22][17];
assign sum_out[6][22][17] = xor_out[30][22][17] + xor_out[31][22][17] + xor_out[32][22][17] + xor_out[33][22][17] + xor_out[34][22][17];
assign sum_out[7][22][17] = xor_out[35][22][17] + xor_out[36][22][17] + xor_out[37][22][17] + xor_out[38][22][17] + xor_out[39][22][17];
assign sum_out[8][22][17] = xor_out[40][22][17] + xor_out[41][22][17] + xor_out[42][22][17] + xor_out[43][22][17] + xor_out[44][22][17];
assign sum_out[9][22][17] = xor_out[45][22][17] + xor_out[46][22][17] + xor_out[47][22][17] + xor_out[48][22][17] + xor_out[49][22][17];
assign sum_out[10][22][17] = xor_out[50][22][17] + xor_out[51][22][17] + xor_out[52][22][17] + xor_out[53][22][17] + xor_out[54][22][17];
assign sum_out[11][22][17] = xor_out[55][22][17] + xor_out[56][22][17] + xor_out[57][22][17] + xor_out[58][22][17] + xor_out[59][22][17];
assign sum_out[12][22][17] = xor_out[60][22][17] + xor_out[61][22][17] + xor_out[62][22][17] + xor_out[63][22][17] + xor_out[64][22][17];
assign sum_out[13][22][17] = xor_out[65][22][17] + xor_out[66][22][17] + xor_out[67][22][17] + xor_out[68][22][17] + xor_out[69][22][17];
assign sum_out[14][22][17] = xor_out[70][22][17] + xor_out[71][22][17] + xor_out[72][22][17] + xor_out[73][22][17] + xor_out[74][22][17];
assign sum_out[15][22][17] = xor_out[75][22][17] + xor_out[76][22][17] + xor_out[77][22][17] + xor_out[78][22][17] + xor_out[79][22][17];
assign sum_out[16][22][17] = xor_out[80][22][17] + xor_out[81][22][17] + xor_out[82][22][17] + xor_out[83][22][17] + xor_out[84][22][17];
assign sum_out[17][22][17] = xor_out[85][22][17] + xor_out[86][22][17] + xor_out[87][22][17] + xor_out[88][22][17] + xor_out[89][22][17];
assign sum_out[18][22][17] = xor_out[90][22][17] + xor_out[91][22][17] + xor_out[92][22][17] + xor_out[93][22][17] + xor_out[94][22][17];
assign sum_out[19][22][17] = xor_out[95][22][17] + xor_out[96][22][17] + xor_out[97][22][17] + xor_out[98][22][17] + xor_out[99][22][17];

assign sum_out[0][22][18] = xor_out[0][22][18] + xor_out[1][22][18] + xor_out[2][22][18] + xor_out[3][22][18] + xor_out[4][22][18];
assign sum_out[1][22][18] = xor_out[5][22][18] + xor_out[6][22][18] + xor_out[7][22][18] + xor_out[8][22][18] + xor_out[9][22][18];
assign sum_out[2][22][18] = xor_out[10][22][18] + xor_out[11][22][18] + xor_out[12][22][18] + xor_out[13][22][18] + xor_out[14][22][18];
assign sum_out[3][22][18] = xor_out[15][22][18] + xor_out[16][22][18] + xor_out[17][22][18] + xor_out[18][22][18] + xor_out[19][22][18];
assign sum_out[4][22][18] = xor_out[20][22][18] + xor_out[21][22][18] + xor_out[22][22][18] + xor_out[23][22][18] + xor_out[24][22][18];
assign sum_out[5][22][18] = xor_out[25][22][18] + xor_out[26][22][18] + xor_out[27][22][18] + xor_out[28][22][18] + xor_out[29][22][18];
assign sum_out[6][22][18] = xor_out[30][22][18] + xor_out[31][22][18] + xor_out[32][22][18] + xor_out[33][22][18] + xor_out[34][22][18];
assign sum_out[7][22][18] = xor_out[35][22][18] + xor_out[36][22][18] + xor_out[37][22][18] + xor_out[38][22][18] + xor_out[39][22][18];
assign sum_out[8][22][18] = xor_out[40][22][18] + xor_out[41][22][18] + xor_out[42][22][18] + xor_out[43][22][18] + xor_out[44][22][18];
assign sum_out[9][22][18] = xor_out[45][22][18] + xor_out[46][22][18] + xor_out[47][22][18] + xor_out[48][22][18] + xor_out[49][22][18];
assign sum_out[10][22][18] = xor_out[50][22][18] + xor_out[51][22][18] + xor_out[52][22][18] + xor_out[53][22][18] + xor_out[54][22][18];
assign sum_out[11][22][18] = xor_out[55][22][18] + xor_out[56][22][18] + xor_out[57][22][18] + xor_out[58][22][18] + xor_out[59][22][18];
assign sum_out[12][22][18] = xor_out[60][22][18] + xor_out[61][22][18] + xor_out[62][22][18] + xor_out[63][22][18] + xor_out[64][22][18];
assign sum_out[13][22][18] = xor_out[65][22][18] + xor_out[66][22][18] + xor_out[67][22][18] + xor_out[68][22][18] + xor_out[69][22][18];
assign sum_out[14][22][18] = xor_out[70][22][18] + xor_out[71][22][18] + xor_out[72][22][18] + xor_out[73][22][18] + xor_out[74][22][18];
assign sum_out[15][22][18] = xor_out[75][22][18] + xor_out[76][22][18] + xor_out[77][22][18] + xor_out[78][22][18] + xor_out[79][22][18];
assign sum_out[16][22][18] = xor_out[80][22][18] + xor_out[81][22][18] + xor_out[82][22][18] + xor_out[83][22][18] + xor_out[84][22][18];
assign sum_out[17][22][18] = xor_out[85][22][18] + xor_out[86][22][18] + xor_out[87][22][18] + xor_out[88][22][18] + xor_out[89][22][18];
assign sum_out[18][22][18] = xor_out[90][22][18] + xor_out[91][22][18] + xor_out[92][22][18] + xor_out[93][22][18] + xor_out[94][22][18];
assign sum_out[19][22][18] = xor_out[95][22][18] + xor_out[96][22][18] + xor_out[97][22][18] + xor_out[98][22][18] + xor_out[99][22][18];

assign sum_out[0][22][19] = xor_out[0][22][19] + xor_out[1][22][19] + xor_out[2][22][19] + xor_out[3][22][19] + xor_out[4][22][19];
assign sum_out[1][22][19] = xor_out[5][22][19] + xor_out[6][22][19] + xor_out[7][22][19] + xor_out[8][22][19] + xor_out[9][22][19];
assign sum_out[2][22][19] = xor_out[10][22][19] + xor_out[11][22][19] + xor_out[12][22][19] + xor_out[13][22][19] + xor_out[14][22][19];
assign sum_out[3][22][19] = xor_out[15][22][19] + xor_out[16][22][19] + xor_out[17][22][19] + xor_out[18][22][19] + xor_out[19][22][19];
assign sum_out[4][22][19] = xor_out[20][22][19] + xor_out[21][22][19] + xor_out[22][22][19] + xor_out[23][22][19] + xor_out[24][22][19];
assign sum_out[5][22][19] = xor_out[25][22][19] + xor_out[26][22][19] + xor_out[27][22][19] + xor_out[28][22][19] + xor_out[29][22][19];
assign sum_out[6][22][19] = xor_out[30][22][19] + xor_out[31][22][19] + xor_out[32][22][19] + xor_out[33][22][19] + xor_out[34][22][19];
assign sum_out[7][22][19] = xor_out[35][22][19] + xor_out[36][22][19] + xor_out[37][22][19] + xor_out[38][22][19] + xor_out[39][22][19];
assign sum_out[8][22][19] = xor_out[40][22][19] + xor_out[41][22][19] + xor_out[42][22][19] + xor_out[43][22][19] + xor_out[44][22][19];
assign sum_out[9][22][19] = xor_out[45][22][19] + xor_out[46][22][19] + xor_out[47][22][19] + xor_out[48][22][19] + xor_out[49][22][19];
assign sum_out[10][22][19] = xor_out[50][22][19] + xor_out[51][22][19] + xor_out[52][22][19] + xor_out[53][22][19] + xor_out[54][22][19];
assign sum_out[11][22][19] = xor_out[55][22][19] + xor_out[56][22][19] + xor_out[57][22][19] + xor_out[58][22][19] + xor_out[59][22][19];
assign sum_out[12][22][19] = xor_out[60][22][19] + xor_out[61][22][19] + xor_out[62][22][19] + xor_out[63][22][19] + xor_out[64][22][19];
assign sum_out[13][22][19] = xor_out[65][22][19] + xor_out[66][22][19] + xor_out[67][22][19] + xor_out[68][22][19] + xor_out[69][22][19];
assign sum_out[14][22][19] = xor_out[70][22][19] + xor_out[71][22][19] + xor_out[72][22][19] + xor_out[73][22][19] + xor_out[74][22][19];
assign sum_out[15][22][19] = xor_out[75][22][19] + xor_out[76][22][19] + xor_out[77][22][19] + xor_out[78][22][19] + xor_out[79][22][19];
assign sum_out[16][22][19] = xor_out[80][22][19] + xor_out[81][22][19] + xor_out[82][22][19] + xor_out[83][22][19] + xor_out[84][22][19];
assign sum_out[17][22][19] = xor_out[85][22][19] + xor_out[86][22][19] + xor_out[87][22][19] + xor_out[88][22][19] + xor_out[89][22][19];
assign sum_out[18][22][19] = xor_out[90][22][19] + xor_out[91][22][19] + xor_out[92][22][19] + xor_out[93][22][19] + xor_out[94][22][19];
assign sum_out[19][22][19] = xor_out[95][22][19] + xor_out[96][22][19] + xor_out[97][22][19] + xor_out[98][22][19] + xor_out[99][22][19];

assign sum_out[0][22][20] = xor_out[0][22][20] + xor_out[1][22][20] + xor_out[2][22][20] + xor_out[3][22][20] + xor_out[4][22][20];
assign sum_out[1][22][20] = xor_out[5][22][20] + xor_out[6][22][20] + xor_out[7][22][20] + xor_out[8][22][20] + xor_out[9][22][20];
assign sum_out[2][22][20] = xor_out[10][22][20] + xor_out[11][22][20] + xor_out[12][22][20] + xor_out[13][22][20] + xor_out[14][22][20];
assign sum_out[3][22][20] = xor_out[15][22][20] + xor_out[16][22][20] + xor_out[17][22][20] + xor_out[18][22][20] + xor_out[19][22][20];
assign sum_out[4][22][20] = xor_out[20][22][20] + xor_out[21][22][20] + xor_out[22][22][20] + xor_out[23][22][20] + xor_out[24][22][20];
assign sum_out[5][22][20] = xor_out[25][22][20] + xor_out[26][22][20] + xor_out[27][22][20] + xor_out[28][22][20] + xor_out[29][22][20];
assign sum_out[6][22][20] = xor_out[30][22][20] + xor_out[31][22][20] + xor_out[32][22][20] + xor_out[33][22][20] + xor_out[34][22][20];
assign sum_out[7][22][20] = xor_out[35][22][20] + xor_out[36][22][20] + xor_out[37][22][20] + xor_out[38][22][20] + xor_out[39][22][20];
assign sum_out[8][22][20] = xor_out[40][22][20] + xor_out[41][22][20] + xor_out[42][22][20] + xor_out[43][22][20] + xor_out[44][22][20];
assign sum_out[9][22][20] = xor_out[45][22][20] + xor_out[46][22][20] + xor_out[47][22][20] + xor_out[48][22][20] + xor_out[49][22][20];
assign sum_out[10][22][20] = xor_out[50][22][20] + xor_out[51][22][20] + xor_out[52][22][20] + xor_out[53][22][20] + xor_out[54][22][20];
assign sum_out[11][22][20] = xor_out[55][22][20] + xor_out[56][22][20] + xor_out[57][22][20] + xor_out[58][22][20] + xor_out[59][22][20];
assign sum_out[12][22][20] = xor_out[60][22][20] + xor_out[61][22][20] + xor_out[62][22][20] + xor_out[63][22][20] + xor_out[64][22][20];
assign sum_out[13][22][20] = xor_out[65][22][20] + xor_out[66][22][20] + xor_out[67][22][20] + xor_out[68][22][20] + xor_out[69][22][20];
assign sum_out[14][22][20] = xor_out[70][22][20] + xor_out[71][22][20] + xor_out[72][22][20] + xor_out[73][22][20] + xor_out[74][22][20];
assign sum_out[15][22][20] = xor_out[75][22][20] + xor_out[76][22][20] + xor_out[77][22][20] + xor_out[78][22][20] + xor_out[79][22][20];
assign sum_out[16][22][20] = xor_out[80][22][20] + xor_out[81][22][20] + xor_out[82][22][20] + xor_out[83][22][20] + xor_out[84][22][20];
assign sum_out[17][22][20] = xor_out[85][22][20] + xor_out[86][22][20] + xor_out[87][22][20] + xor_out[88][22][20] + xor_out[89][22][20];
assign sum_out[18][22][20] = xor_out[90][22][20] + xor_out[91][22][20] + xor_out[92][22][20] + xor_out[93][22][20] + xor_out[94][22][20];
assign sum_out[19][22][20] = xor_out[95][22][20] + xor_out[96][22][20] + xor_out[97][22][20] + xor_out[98][22][20] + xor_out[99][22][20];

assign sum_out[0][22][21] = xor_out[0][22][21] + xor_out[1][22][21] + xor_out[2][22][21] + xor_out[3][22][21] + xor_out[4][22][21];
assign sum_out[1][22][21] = xor_out[5][22][21] + xor_out[6][22][21] + xor_out[7][22][21] + xor_out[8][22][21] + xor_out[9][22][21];
assign sum_out[2][22][21] = xor_out[10][22][21] + xor_out[11][22][21] + xor_out[12][22][21] + xor_out[13][22][21] + xor_out[14][22][21];
assign sum_out[3][22][21] = xor_out[15][22][21] + xor_out[16][22][21] + xor_out[17][22][21] + xor_out[18][22][21] + xor_out[19][22][21];
assign sum_out[4][22][21] = xor_out[20][22][21] + xor_out[21][22][21] + xor_out[22][22][21] + xor_out[23][22][21] + xor_out[24][22][21];
assign sum_out[5][22][21] = xor_out[25][22][21] + xor_out[26][22][21] + xor_out[27][22][21] + xor_out[28][22][21] + xor_out[29][22][21];
assign sum_out[6][22][21] = xor_out[30][22][21] + xor_out[31][22][21] + xor_out[32][22][21] + xor_out[33][22][21] + xor_out[34][22][21];
assign sum_out[7][22][21] = xor_out[35][22][21] + xor_out[36][22][21] + xor_out[37][22][21] + xor_out[38][22][21] + xor_out[39][22][21];
assign sum_out[8][22][21] = xor_out[40][22][21] + xor_out[41][22][21] + xor_out[42][22][21] + xor_out[43][22][21] + xor_out[44][22][21];
assign sum_out[9][22][21] = xor_out[45][22][21] + xor_out[46][22][21] + xor_out[47][22][21] + xor_out[48][22][21] + xor_out[49][22][21];
assign sum_out[10][22][21] = xor_out[50][22][21] + xor_out[51][22][21] + xor_out[52][22][21] + xor_out[53][22][21] + xor_out[54][22][21];
assign sum_out[11][22][21] = xor_out[55][22][21] + xor_out[56][22][21] + xor_out[57][22][21] + xor_out[58][22][21] + xor_out[59][22][21];
assign sum_out[12][22][21] = xor_out[60][22][21] + xor_out[61][22][21] + xor_out[62][22][21] + xor_out[63][22][21] + xor_out[64][22][21];
assign sum_out[13][22][21] = xor_out[65][22][21] + xor_out[66][22][21] + xor_out[67][22][21] + xor_out[68][22][21] + xor_out[69][22][21];
assign sum_out[14][22][21] = xor_out[70][22][21] + xor_out[71][22][21] + xor_out[72][22][21] + xor_out[73][22][21] + xor_out[74][22][21];
assign sum_out[15][22][21] = xor_out[75][22][21] + xor_out[76][22][21] + xor_out[77][22][21] + xor_out[78][22][21] + xor_out[79][22][21];
assign sum_out[16][22][21] = xor_out[80][22][21] + xor_out[81][22][21] + xor_out[82][22][21] + xor_out[83][22][21] + xor_out[84][22][21];
assign sum_out[17][22][21] = xor_out[85][22][21] + xor_out[86][22][21] + xor_out[87][22][21] + xor_out[88][22][21] + xor_out[89][22][21];
assign sum_out[18][22][21] = xor_out[90][22][21] + xor_out[91][22][21] + xor_out[92][22][21] + xor_out[93][22][21] + xor_out[94][22][21];
assign sum_out[19][22][21] = xor_out[95][22][21] + xor_out[96][22][21] + xor_out[97][22][21] + xor_out[98][22][21] + xor_out[99][22][21];

assign sum_out[0][22][22] = xor_out[0][22][22] + xor_out[1][22][22] + xor_out[2][22][22] + xor_out[3][22][22] + xor_out[4][22][22];
assign sum_out[1][22][22] = xor_out[5][22][22] + xor_out[6][22][22] + xor_out[7][22][22] + xor_out[8][22][22] + xor_out[9][22][22];
assign sum_out[2][22][22] = xor_out[10][22][22] + xor_out[11][22][22] + xor_out[12][22][22] + xor_out[13][22][22] + xor_out[14][22][22];
assign sum_out[3][22][22] = xor_out[15][22][22] + xor_out[16][22][22] + xor_out[17][22][22] + xor_out[18][22][22] + xor_out[19][22][22];
assign sum_out[4][22][22] = xor_out[20][22][22] + xor_out[21][22][22] + xor_out[22][22][22] + xor_out[23][22][22] + xor_out[24][22][22];
assign sum_out[5][22][22] = xor_out[25][22][22] + xor_out[26][22][22] + xor_out[27][22][22] + xor_out[28][22][22] + xor_out[29][22][22];
assign sum_out[6][22][22] = xor_out[30][22][22] + xor_out[31][22][22] + xor_out[32][22][22] + xor_out[33][22][22] + xor_out[34][22][22];
assign sum_out[7][22][22] = xor_out[35][22][22] + xor_out[36][22][22] + xor_out[37][22][22] + xor_out[38][22][22] + xor_out[39][22][22];
assign sum_out[8][22][22] = xor_out[40][22][22] + xor_out[41][22][22] + xor_out[42][22][22] + xor_out[43][22][22] + xor_out[44][22][22];
assign sum_out[9][22][22] = xor_out[45][22][22] + xor_out[46][22][22] + xor_out[47][22][22] + xor_out[48][22][22] + xor_out[49][22][22];
assign sum_out[10][22][22] = xor_out[50][22][22] + xor_out[51][22][22] + xor_out[52][22][22] + xor_out[53][22][22] + xor_out[54][22][22];
assign sum_out[11][22][22] = xor_out[55][22][22] + xor_out[56][22][22] + xor_out[57][22][22] + xor_out[58][22][22] + xor_out[59][22][22];
assign sum_out[12][22][22] = xor_out[60][22][22] + xor_out[61][22][22] + xor_out[62][22][22] + xor_out[63][22][22] + xor_out[64][22][22];
assign sum_out[13][22][22] = xor_out[65][22][22] + xor_out[66][22][22] + xor_out[67][22][22] + xor_out[68][22][22] + xor_out[69][22][22];
assign sum_out[14][22][22] = xor_out[70][22][22] + xor_out[71][22][22] + xor_out[72][22][22] + xor_out[73][22][22] + xor_out[74][22][22];
assign sum_out[15][22][22] = xor_out[75][22][22] + xor_out[76][22][22] + xor_out[77][22][22] + xor_out[78][22][22] + xor_out[79][22][22];
assign sum_out[16][22][22] = xor_out[80][22][22] + xor_out[81][22][22] + xor_out[82][22][22] + xor_out[83][22][22] + xor_out[84][22][22];
assign sum_out[17][22][22] = xor_out[85][22][22] + xor_out[86][22][22] + xor_out[87][22][22] + xor_out[88][22][22] + xor_out[89][22][22];
assign sum_out[18][22][22] = xor_out[90][22][22] + xor_out[91][22][22] + xor_out[92][22][22] + xor_out[93][22][22] + xor_out[94][22][22];
assign sum_out[19][22][22] = xor_out[95][22][22] + xor_out[96][22][22] + xor_out[97][22][22] + xor_out[98][22][22] + xor_out[99][22][22];

assign sum_out[0][22][23] = xor_out[0][22][23] + xor_out[1][22][23] + xor_out[2][22][23] + xor_out[3][22][23] + xor_out[4][22][23];
assign sum_out[1][22][23] = xor_out[5][22][23] + xor_out[6][22][23] + xor_out[7][22][23] + xor_out[8][22][23] + xor_out[9][22][23];
assign sum_out[2][22][23] = xor_out[10][22][23] + xor_out[11][22][23] + xor_out[12][22][23] + xor_out[13][22][23] + xor_out[14][22][23];
assign sum_out[3][22][23] = xor_out[15][22][23] + xor_out[16][22][23] + xor_out[17][22][23] + xor_out[18][22][23] + xor_out[19][22][23];
assign sum_out[4][22][23] = xor_out[20][22][23] + xor_out[21][22][23] + xor_out[22][22][23] + xor_out[23][22][23] + xor_out[24][22][23];
assign sum_out[5][22][23] = xor_out[25][22][23] + xor_out[26][22][23] + xor_out[27][22][23] + xor_out[28][22][23] + xor_out[29][22][23];
assign sum_out[6][22][23] = xor_out[30][22][23] + xor_out[31][22][23] + xor_out[32][22][23] + xor_out[33][22][23] + xor_out[34][22][23];
assign sum_out[7][22][23] = xor_out[35][22][23] + xor_out[36][22][23] + xor_out[37][22][23] + xor_out[38][22][23] + xor_out[39][22][23];
assign sum_out[8][22][23] = xor_out[40][22][23] + xor_out[41][22][23] + xor_out[42][22][23] + xor_out[43][22][23] + xor_out[44][22][23];
assign sum_out[9][22][23] = xor_out[45][22][23] + xor_out[46][22][23] + xor_out[47][22][23] + xor_out[48][22][23] + xor_out[49][22][23];
assign sum_out[10][22][23] = xor_out[50][22][23] + xor_out[51][22][23] + xor_out[52][22][23] + xor_out[53][22][23] + xor_out[54][22][23];
assign sum_out[11][22][23] = xor_out[55][22][23] + xor_out[56][22][23] + xor_out[57][22][23] + xor_out[58][22][23] + xor_out[59][22][23];
assign sum_out[12][22][23] = xor_out[60][22][23] + xor_out[61][22][23] + xor_out[62][22][23] + xor_out[63][22][23] + xor_out[64][22][23];
assign sum_out[13][22][23] = xor_out[65][22][23] + xor_out[66][22][23] + xor_out[67][22][23] + xor_out[68][22][23] + xor_out[69][22][23];
assign sum_out[14][22][23] = xor_out[70][22][23] + xor_out[71][22][23] + xor_out[72][22][23] + xor_out[73][22][23] + xor_out[74][22][23];
assign sum_out[15][22][23] = xor_out[75][22][23] + xor_out[76][22][23] + xor_out[77][22][23] + xor_out[78][22][23] + xor_out[79][22][23];
assign sum_out[16][22][23] = xor_out[80][22][23] + xor_out[81][22][23] + xor_out[82][22][23] + xor_out[83][22][23] + xor_out[84][22][23];
assign sum_out[17][22][23] = xor_out[85][22][23] + xor_out[86][22][23] + xor_out[87][22][23] + xor_out[88][22][23] + xor_out[89][22][23];
assign sum_out[18][22][23] = xor_out[90][22][23] + xor_out[91][22][23] + xor_out[92][22][23] + xor_out[93][22][23] + xor_out[94][22][23];
assign sum_out[19][22][23] = xor_out[95][22][23] + xor_out[96][22][23] + xor_out[97][22][23] + xor_out[98][22][23] + xor_out[99][22][23];

assign sum_out[0][23][0] = xor_out[0][23][0] + xor_out[1][23][0] + xor_out[2][23][0] + xor_out[3][23][0] + xor_out[4][23][0];
assign sum_out[1][23][0] = xor_out[5][23][0] + xor_out[6][23][0] + xor_out[7][23][0] + xor_out[8][23][0] + xor_out[9][23][0];
assign sum_out[2][23][0] = xor_out[10][23][0] + xor_out[11][23][0] + xor_out[12][23][0] + xor_out[13][23][0] + xor_out[14][23][0];
assign sum_out[3][23][0] = xor_out[15][23][0] + xor_out[16][23][0] + xor_out[17][23][0] + xor_out[18][23][0] + xor_out[19][23][0];
assign sum_out[4][23][0] = xor_out[20][23][0] + xor_out[21][23][0] + xor_out[22][23][0] + xor_out[23][23][0] + xor_out[24][23][0];
assign sum_out[5][23][0] = xor_out[25][23][0] + xor_out[26][23][0] + xor_out[27][23][0] + xor_out[28][23][0] + xor_out[29][23][0];
assign sum_out[6][23][0] = xor_out[30][23][0] + xor_out[31][23][0] + xor_out[32][23][0] + xor_out[33][23][0] + xor_out[34][23][0];
assign sum_out[7][23][0] = xor_out[35][23][0] + xor_out[36][23][0] + xor_out[37][23][0] + xor_out[38][23][0] + xor_out[39][23][0];
assign sum_out[8][23][0] = xor_out[40][23][0] + xor_out[41][23][0] + xor_out[42][23][0] + xor_out[43][23][0] + xor_out[44][23][0];
assign sum_out[9][23][0] = xor_out[45][23][0] + xor_out[46][23][0] + xor_out[47][23][0] + xor_out[48][23][0] + xor_out[49][23][0];
assign sum_out[10][23][0] = xor_out[50][23][0] + xor_out[51][23][0] + xor_out[52][23][0] + xor_out[53][23][0] + xor_out[54][23][0];
assign sum_out[11][23][0] = xor_out[55][23][0] + xor_out[56][23][0] + xor_out[57][23][0] + xor_out[58][23][0] + xor_out[59][23][0];
assign sum_out[12][23][0] = xor_out[60][23][0] + xor_out[61][23][0] + xor_out[62][23][0] + xor_out[63][23][0] + xor_out[64][23][0];
assign sum_out[13][23][0] = xor_out[65][23][0] + xor_out[66][23][0] + xor_out[67][23][0] + xor_out[68][23][0] + xor_out[69][23][0];
assign sum_out[14][23][0] = xor_out[70][23][0] + xor_out[71][23][0] + xor_out[72][23][0] + xor_out[73][23][0] + xor_out[74][23][0];
assign sum_out[15][23][0] = xor_out[75][23][0] + xor_out[76][23][0] + xor_out[77][23][0] + xor_out[78][23][0] + xor_out[79][23][0];
assign sum_out[16][23][0] = xor_out[80][23][0] + xor_out[81][23][0] + xor_out[82][23][0] + xor_out[83][23][0] + xor_out[84][23][0];
assign sum_out[17][23][0] = xor_out[85][23][0] + xor_out[86][23][0] + xor_out[87][23][0] + xor_out[88][23][0] + xor_out[89][23][0];
assign sum_out[18][23][0] = xor_out[90][23][0] + xor_out[91][23][0] + xor_out[92][23][0] + xor_out[93][23][0] + xor_out[94][23][0];
assign sum_out[19][23][0] = xor_out[95][23][0] + xor_out[96][23][0] + xor_out[97][23][0] + xor_out[98][23][0] + xor_out[99][23][0];

assign sum_out[0][23][1] = xor_out[0][23][1] + xor_out[1][23][1] + xor_out[2][23][1] + xor_out[3][23][1] + xor_out[4][23][1];
assign sum_out[1][23][1] = xor_out[5][23][1] + xor_out[6][23][1] + xor_out[7][23][1] + xor_out[8][23][1] + xor_out[9][23][1];
assign sum_out[2][23][1] = xor_out[10][23][1] + xor_out[11][23][1] + xor_out[12][23][1] + xor_out[13][23][1] + xor_out[14][23][1];
assign sum_out[3][23][1] = xor_out[15][23][1] + xor_out[16][23][1] + xor_out[17][23][1] + xor_out[18][23][1] + xor_out[19][23][1];
assign sum_out[4][23][1] = xor_out[20][23][1] + xor_out[21][23][1] + xor_out[22][23][1] + xor_out[23][23][1] + xor_out[24][23][1];
assign sum_out[5][23][1] = xor_out[25][23][1] + xor_out[26][23][1] + xor_out[27][23][1] + xor_out[28][23][1] + xor_out[29][23][1];
assign sum_out[6][23][1] = xor_out[30][23][1] + xor_out[31][23][1] + xor_out[32][23][1] + xor_out[33][23][1] + xor_out[34][23][1];
assign sum_out[7][23][1] = xor_out[35][23][1] + xor_out[36][23][1] + xor_out[37][23][1] + xor_out[38][23][1] + xor_out[39][23][1];
assign sum_out[8][23][1] = xor_out[40][23][1] + xor_out[41][23][1] + xor_out[42][23][1] + xor_out[43][23][1] + xor_out[44][23][1];
assign sum_out[9][23][1] = xor_out[45][23][1] + xor_out[46][23][1] + xor_out[47][23][1] + xor_out[48][23][1] + xor_out[49][23][1];
assign sum_out[10][23][1] = xor_out[50][23][1] + xor_out[51][23][1] + xor_out[52][23][1] + xor_out[53][23][1] + xor_out[54][23][1];
assign sum_out[11][23][1] = xor_out[55][23][1] + xor_out[56][23][1] + xor_out[57][23][1] + xor_out[58][23][1] + xor_out[59][23][1];
assign sum_out[12][23][1] = xor_out[60][23][1] + xor_out[61][23][1] + xor_out[62][23][1] + xor_out[63][23][1] + xor_out[64][23][1];
assign sum_out[13][23][1] = xor_out[65][23][1] + xor_out[66][23][1] + xor_out[67][23][1] + xor_out[68][23][1] + xor_out[69][23][1];
assign sum_out[14][23][1] = xor_out[70][23][1] + xor_out[71][23][1] + xor_out[72][23][1] + xor_out[73][23][1] + xor_out[74][23][1];
assign sum_out[15][23][1] = xor_out[75][23][1] + xor_out[76][23][1] + xor_out[77][23][1] + xor_out[78][23][1] + xor_out[79][23][1];
assign sum_out[16][23][1] = xor_out[80][23][1] + xor_out[81][23][1] + xor_out[82][23][1] + xor_out[83][23][1] + xor_out[84][23][1];
assign sum_out[17][23][1] = xor_out[85][23][1] + xor_out[86][23][1] + xor_out[87][23][1] + xor_out[88][23][1] + xor_out[89][23][1];
assign sum_out[18][23][1] = xor_out[90][23][1] + xor_out[91][23][1] + xor_out[92][23][1] + xor_out[93][23][1] + xor_out[94][23][1];
assign sum_out[19][23][1] = xor_out[95][23][1] + xor_out[96][23][1] + xor_out[97][23][1] + xor_out[98][23][1] + xor_out[99][23][1];

assign sum_out[0][23][2] = xor_out[0][23][2] + xor_out[1][23][2] + xor_out[2][23][2] + xor_out[3][23][2] + xor_out[4][23][2];
assign sum_out[1][23][2] = xor_out[5][23][2] + xor_out[6][23][2] + xor_out[7][23][2] + xor_out[8][23][2] + xor_out[9][23][2];
assign sum_out[2][23][2] = xor_out[10][23][2] + xor_out[11][23][2] + xor_out[12][23][2] + xor_out[13][23][2] + xor_out[14][23][2];
assign sum_out[3][23][2] = xor_out[15][23][2] + xor_out[16][23][2] + xor_out[17][23][2] + xor_out[18][23][2] + xor_out[19][23][2];
assign sum_out[4][23][2] = xor_out[20][23][2] + xor_out[21][23][2] + xor_out[22][23][2] + xor_out[23][23][2] + xor_out[24][23][2];
assign sum_out[5][23][2] = xor_out[25][23][2] + xor_out[26][23][2] + xor_out[27][23][2] + xor_out[28][23][2] + xor_out[29][23][2];
assign sum_out[6][23][2] = xor_out[30][23][2] + xor_out[31][23][2] + xor_out[32][23][2] + xor_out[33][23][2] + xor_out[34][23][2];
assign sum_out[7][23][2] = xor_out[35][23][2] + xor_out[36][23][2] + xor_out[37][23][2] + xor_out[38][23][2] + xor_out[39][23][2];
assign sum_out[8][23][2] = xor_out[40][23][2] + xor_out[41][23][2] + xor_out[42][23][2] + xor_out[43][23][2] + xor_out[44][23][2];
assign sum_out[9][23][2] = xor_out[45][23][2] + xor_out[46][23][2] + xor_out[47][23][2] + xor_out[48][23][2] + xor_out[49][23][2];
assign sum_out[10][23][2] = xor_out[50][23][2] + xor_out[51][23][2] + xor_out[52][23][2] + xor_out[53][23][2] + xor_out[54][23][2];
assign sum_out[11][23][2] = xor_out[55][23][2] + xor_out[56][23][2] + xor_out[57][23][2] + xor_out[58][23][2] + xor_out[59][23][2];
assign sum_out[12][23][2] = xor_out[60][23][2] + xor_out[61][23][2] + xor_out[62][23][2] + xor_out[63][23][2] + xor_out[64][23][2];
assign sum_out[13][23][2] = xor_out[65][23][2] + xor_out[66][23][2] + xor_out[67][23][2] + xor_out[68][23][2] + xor_out[69][23][2];
assign sum_out[14][23][2] = xor_out[70][23][2] + xor_out[71][23][2] + xor_out[72][23][2] + xor_out[73][23][2] + xor_out[74][23][2];
assign sum_out[15][23][2] = xor_out[75][23][2] + xor_out[76][23][2] + xor_out[77][23][2] + xor_out[78][23][2] + xor_out[79][23][2];
assign sum_out[16][23][2] = xor_out[80][23][2] + xor_out[81][23][2] + xor_out[82][23][2] + xor_out[83][23][2] + xor_out[84][23][2];
assign sum_out[17][23][2] = xor_out[85][23][2] + xor_out[86][23][2] + xor_out[87][23][2] + xor_out[88][23][2] + xor_out[89][23][2];
assign sum_out[18][23][2] = xor_out[90][23][2] + xor_out[91][23][2] + xor_out[92][23][2] + xor_out[93][23][2] + xor_out[94][23][2];
assign sum_out[19][23][2] = xor_out[95][23][2] + xor_out[96][23][2] + xor_out[97][23][2] + xor_out[98][23][2] + xor_out[99][23][2];

assign sum_out[0][23][3] = xor_out[0][23][3] + xor_out[1][23][3] + xor_out[2][23][3] + xor_out[3][23][3] + xor_out[4][23][3];
assign sum_out[1][23][3] = xor_out[5][23][3] + xor_out[6][23][3] + xor_out[7][23][3] + xor_out[8][23][3] + xor_out[9][23][3];
assign sum_out[2][23][3] = xor_out[10][23][3] + xor_out[11][23][3] + xor_out[12][23][3] + xor_out[13][23][3] + xor_out[14][23][3];
assign sum_out[3][23][3] = xor_out[15][23][3] + xor_out[16][23][3] + xor_out[17][23][3] + xor_out[18][23][3] + xor_out[19][23][3];
assign sum_out[4][23][3] = xor_out[20][23][3] + xor_out[21][23][3] + xor_out[22][23][3] + xor_out[23][23][3] + xor_out[24][23][3];
assign sum_out[5][23][3] = xor_out[25][23][3] + xor_out[26][23][3] + xor_out[27][23][3] + xor_out[28][23][3] + xor_out[29][23][3];
assign sum_out[6][23][3] = xor_out[30][23][3] + xor_out[31][23][3] + xor_out[32][23][3] + xor_out[33][23][3] + xor_out[34][23][3];
assign sum_out[7][23][3] = xor_out[35][23][3] + xor_out[36][23][3] + xor_out[37][23][3] + xor_out[38][23][3] + xor_out[39][23][3];
assign sum_out[8][23][3] = xor_out[40][23][3] + xor_out[41][23][3] + xor_out[42][23][3] + xor_out[43][23][3] + xor_out[44][23][3];
assign sum_out[9][23][3] = xor_out[45][23][3] + xor_out[46][23][3] + xor_out[47][23][3] + xor_out[48][23][3] + xor_out[49][23][3];
assign sum_out[10][23][3] = xor_out[50][23][3] + xor_out[51][23][3] + xor_out[52][23][3] + xor_out[53][23][3] + xor_out[54][23][3];
assign sum_out[11][23][3] = xor_out[55][23][3] + xor_out[56][23][3] + xor_out[57][23][3] + xor_out[58][23][3] + xor_out[59][23][3];
assign sum_out[12][23][3] = xor_out[60][23][3] + xor_out[61][23][3] + xor_out[62][23][3] + xor_out[63][23][3] + xor_out[64][23][3];
assign sum_out[13][23][3] = xor_out[65][23][3] + xor_out[66][23][3] + xor_out[67][23][3] + xor_out[68][23][3] + xor_out[69][23][3];
assign sum_out[14][23][3] = xor_out[70][23][3] + xor_out[71][23][3] + xor_out[72][23][3] + xor_out[73][23][3] + xor_out[74][23][3];
assign sum_out[15][23][3] = xor_out[75][23][3] + xor_out[76][23][3] + xor_out[77][23][3] + xor_out[78][23][3] + xor_out[79][23][3];
assign sum_out[16][23][3] = xor_out[80][23][3] + xor_out[81][23][3] + xor_out[82][23][3] + xor_out[83][23][3] + xor_out[84][23][3];
assign sum_out[17][23][3] = xor_out[85][23][3] + xor_out[86][23][3] + xor_out[87][23][3] + xor_out[88][23][3] + xor_out[89][23][3];
assign sum_out[18][23][3] = xor_out[90][23][3] + xor_out[91][23][3] + xor_out[92][23][3] + xor_out[93][23][3] + xor_out[94][23][3];
assign sum_out[19][23][3] = xor_out[95][23][3] + xor_out[96][23][3] + xor_out[97][23][3] + xor_out[98][23][3] + xor_out[99][23][3];

assign sum_out[0][23][4] = xor_out[0][23][4] + xor_out[1][23][4] + xor_out[2][23][4] + xor_out[3][23][4] + xor_out[4][23][4];
assign sum_out[1][23][4] = xor_out[5][23][4] + xor_out[6][23][4] + xor_out[7][23][4] + xor_out[8][23][4] + xor_out[9][23][4];
assign sum_out[2][23][4] = xor_out[10][23][4] + xor_out[11][23][4] + xor_out[12][23][4] + xor_out[13][23][4] + xor_out[14][23][4];
assign sum_out[3][23][4] = xor_out[15][23][4] + xor_out[16][23][4] + xor_out[17][23][4] + xor_out[18][23][4] + xor_out[19][23][4];
assign sum_out[4][23][4] = xor_out[20][23][4] + xor_out[21][23][4] + xor_out[22][23][4] + xor_out[23][23][4] + xor_out[24][23][4];
assign sum_out[5][23][4] = xor_out[25][23][4] + xor_out[26][23][4] + xor_out[27][23][4] + xor_out[28][23][4] + xor_out[29][23][4];
assign sum_out[6][23][4] = xor_out[30][23][4] + xor_out[31][23][4] + xor_out[32][23][4] + xor_out[33][23][4] + xor_out[34][23][4];
assign sum_out[7][23][4] = xor_out[35][23][4] + xor_out[36][23][4] + xor_out[37][23][4] + xor_out[38][23][4] + xor_out[39][23][4];
assign sum_out[8][23][4] = xor_out[40][23][4] + xor_out[41][23][4] + xor_out[42][23][4] + xor_out[43][23][4] + xor_out[44][23][4];
assign sum_out[9][23][4] = xor_out[45][23][4] + xor_out[46][23][4] + xor_out[47][23][4] + xor_out[48][23][4] + xor_out[49][23][4];
assign sum_out[10][23][4] = xor_out[50][23][4] + xor_out[51][23][4] + xor_out[52][23][4] + xor_out[53][23][4] + xor_out[54][23][4];
assign sum_out[11][23][4] = xor_out[55][23][4] + xor_out[56][23][4] + xor_out[57][23][4] + xor_out[58][23][4] + xor_out[59][23][4];
assign sum_out[12][23][4] = xor_out[60][23][4] + xor_out[61][23][4] + xor_out[62][23][4] + xor_out[63][23][4] + xor_out[64][23][4];
assign sum_out[13][23][4] = xor_out[65][23][4] + xor_out[66][23][4] + xor_out[67][23][4] + xor_out[68][23][4] + xor_out[69][23][4];
assign sum_out[14][23][4] = xor_out[70][23][4] + xor_out[71][23][4] + xor_out[72][23][4] + xor_out[73][23][4] + xor_out[74][23][4];
assign sum_out[15][23][4] = xor_out[75][23][4] + xor_out[76][23][4] + xor_out[77][23][4] + xor_out[78][23][4] + xor_out[79][23][4];
assign sum_out[16][23][4] = xor_out[80][23][4] + xor_out[81][23][4] + xor_out[82][23][4] + xor_out[83][23][4] + xor_out[84][23][4];
assign sum_out[17][23][4] = xor_out[85][23][4] + xor_out[86][23][4] + xor_out[87][23][4] + xor_out[88][23][4] + xor_out[89][23][4];
assign sum_out[18][23][4] = xor_out[90][23][4] + xor_out[91][23][4] + xor_out[92][23][4] + xor_out[93][23][4] + xor_out[94][23][4];
assign sum_out[19][23][4] = xor_out[95][23][4] + xor_out[96][23][4] + xor_out[97][23][4] + xor_out[98][23][4] + xor_out[99][23][4];

assign sum_out[0][23][5] = xor_out[0][23][5] + xor_out[1][23][5] + xor_out[2][23][5] + xor_out[3][23][5] + xor_out[4][23][5];
assign sum_out[1][23][5] = xor_out[5][23][5] + xor_out[6][23][5] + xor_out[7][23][5] + xor_out[8][23][5] + xor_out[9][23][5];
assign sum_out[2][23][5] = xor_out[10][23][5] + xor_out[11][23][5] + xor_out[12][23][5] + xor_out[13][23][5] + xor_out[14][23][5];
assign sum_out[3][23][5] = xor_out[15][23][5] + xor_out[16][23][5] + xor_out[17][23][5] + xor_out[18][23][5] + xor_out[19][23][5];
assign sum_out[4][23][5] = xor_out[20][23][5] + xor_out[21][23][5] + xor_out[22][23][5] + xor_out[23][23][5] + xor_out[24][23][5];
assign sum_out[5][23][5] = xor_out[25][23][5] + xor_out[26][23][5] + xor_out[27][23][5] + xor_out[28][23][5] + xor_out[29][23][5];
assign sum_out[6][23][5] = xor_out[30][23][5] + xor_out[31][23][5] + xor_out[32][23][5] + xor_out[33][23][5] + xor_out[34][23][5];
assign sum_out[7][23][5] = xor_out[35][23][5] + xor_out[36][23][5] + xor_out[37][23][5] + xor_out[38][23][5] + xor_out[39][23][5];
assign sum_out[8][23][5] = xor_out[40][23][5] + xor_out[41][23][5] + xor_out[42][23][5] + xor_out[43][23][5] + xor_out[44][23][5];
assign sum_out[9][23][5] = xor_out[45][23][5] + xor_out[46][23][5] + xor_out[47][23][5] + xor_out[48][23][5] + xor_out[49][23][5];
assign sum_out[10][23][5] = xor_out[50][23][5] + xor_out[51][23][5] + xor_out[52][23][5] + xor_out[53][23][5] + xor_out[54][23][5];
assign sum_out[11][23][5] = xor_out[55][23][5] + xor_out[56][23][5] + xor_out[57][23][5] + xor_out[58][23][5] + xor_out[59][23][5];
assign sum_out[12][23][5] = xor_out[60][23][5] + xor_out[61][23][5] + xor_out[62][23][5] + xor_out[63][23][5] + xor_out[64][23][5];
assign sum_out[13][23][5] = xor_out[65][23][5] + xor_out[66][23][5] + xor_out[67][23][5] + xor_out[68][23][5] + xor_out[69][23][5];
assign sum_out[14][23][5] = xor_out[70][23][5] + xor_out[71][23][5] + xor_out[72][23][5] + xor_out[73][23][5] + xor_out[74][23][5];
assign sum_out[15][23][5] = xor_out[75][23][5] + xor_out[76][23][5] + xor_out[77][23][5] + xor_out[78][23][5] + xor_out[79][23][5];
assign sum_out[16][23][5] = xor_out[80][23][5] + xor_out[81][23][5] + xor_out[82][23][5] + xor_out[83][23][5] + xor_out[84][23][5];
assign sum_out[17][23][5] = xor_out[85][23][5] + xor_out[86][23][5] + xor_out[87][23][5] + xor_out[88][23][5] + xor_out[89][23][5];
assign sum_out[18][23][5] = xor_out[90][23][5] + xor_out[91][23][5] + xor_out[92][23][5] + xor_out[93][23][5] + xor_out[94][23][5];
assign sum_out[19][23][5] = xor_out[95][23][5] + xor_out[96][23][5] + xor_out[97][23][5] + xor_out[98][23][5] + xor_out[99][23][5];

assign sum_out[0][23][6] = xor_out[0][23][6] + xor_out[1][23][6] + xor_out[2][23][6] + xor_out[3][23][6] + xor_out[4][23][6];
assign sum_out[1][23][6] = xor_out[5][23][6] + xor_out[6][23][6] + xor_out[7][23][6] + xor_out[8][23][6] + xor_out[9][23][6];
assign sum_out[2][23][6] = xor_out[10][23][6] + xor_out[11][23][6] + xor_out[12][23][6] + xor_out[13][23][6] + xor_out[14][23][6];
assign sum_out[3][23][6] = xor_out[15][23][6] + xor_out[16][23][6] + xor_out[17][23][6] + xor_out[18][23][6] + xor_out[19][23][6];
assign sum_out[4][23][6] = xor_out[20][23][6] + xor_out[21][23][6] + xor_out[22][23][6] + xor_out[23][23][6] + xor_out[24][23][6];
assign sum_out[5][23][6] = xor_out[25][23][6] + xor_out[26][23][6] + xor_out[27][23][6] + xor_out[28][23][6] + xor_out[29][23][6];
assign sum_out[6][23][6] = xor_out[30][23][6] + xor_out[31][23][6] + xor_out[32][23][6] + xor_out[33][23][6] + xor_out[34][23][6];
assign sum_out[7][23][6] = xor_out[35][23][6] + xor_out[36][23][6] + xor_out[37][23][6] + xor_out[38][23][6] + xor_out[39][23][6];
assign sum_out[8][23][6] = xor_out[40][23][6] + xor_out[41][23][6] + xor_out[42][23][6] + xor_out[43][23][6] + xor_out[44][23][6];
assign sum_out[9][23][6] = xor_out[45][23][6] + xor_out[46][23][6] + xor_out[47][23][6] + xor_out[48][23][6] + xor_out[49][23][6];
assign sum_out[10][23][6] = xor_out[50][23][6] + xor_out[51][23][6] + xor_out[52][23][6] + xor_out[53][23][6] + xor_out[54][23][6];
assign sum_out[11][23][6] = xor_out[55][23][6] + xor_out[56][23][6] + xor_out[57][23][6] + xor_out[58][23][6] + xor_out[59][23][6];
assign sum_out[12][23][6] = xor_out[60][23][6] + xor_out[61][23][6] + xor_out[62][23][6] + xor_out[63][23][6] + xor_out[64][23][6];
assign sum_out[13][23][6] = xor_out[65][23][6] + xor_out[66][23][6] + xor_out[67][23][6] + xor_out[68][23][6] + xor_out[69][23][6];
assign sum_out[14][23][6] = xor_out[70][23][6] + xor_out[71][23][6] + xor_out[72][23][6] + xor_out[73][23][6] + xor_out[74][23][6];
assign sum_out[15][23][6] = xor_out[75][23][6] + xor_out[76][23][6] + xor_out[77][23][6] + xor_out[78][23][6] + xor_out[79][23][6];
assign sum_out[16][23][6] = xor_out[80][23][6] + xor_out[81][23][6] + xor_out[82][23][6] + xor_out[83][23][6] + xor_out[84][23][6];
assign sum_out[17][23][6] = xor_out[85][23][6] + xor_out[86][23][6] + xor_out[87][23][6] + xor_out[88][23][6] + xor_out[89][23][6];
assign sum_out[18][23][6] = xor_out[90][23][6] + xor_out[91][23][6] + xor_out[92][23][6] + xor_out[93][23][6] + xor_out[94][23][6];
assign sum_out[19][23][6] = xor_out[95][23][6] + xor_out[96][23][6] + xor_out[97][23][6] + xor_out[98][23][6] + xor_out[99][23][6];

assign sum_out[0][23][7] = xor_out[0][23][7] + xor_out[1][23][7] + xor_out[2][23][7] + xor_out[3][23][7] + xor_out[4][23][7];
assign sum_out[1][23][7] = xor_out[5][23][7] + xor_out[6][23][7] + xor_out[7][23][7] + xor_out[8][23][7] + xor_out[9][23][7];
assign sum_out[2][23][7] = xor_out[10][23][7] + xor_out[11][23][7] + xor_out[12][23][7] + xor_out[13][23][7] + xor_out[14][23][7];
assign sum_out[3][23][7] = xor_out[15][23][7] + xor_out[16][23][7] + xor_out[17][23][7] + xor_out[18][23][7] + xor_out[19][23][7];
assign sum_out[4][23][7] = xor_out[20][23][7] + xor_out[21][23][7] + xor_out[22][23][7] + xor_out[23][23][7] + xor_out[24][23][7];
assign sum_out[5][23][7] = xor_out[25][23][7] + xor_out[26][23][7] + xor_out[27][23][7] + xor_out[28][23][7] + xor_out[29][23][7];
assign sum_out[6][23][7] = xor_out[30][23][7] + xor_out[31][23][7] + xor_out[32][23][7] + xor_out[33][23][7] + xor_out[34][23][7];
assign sum_out[7][23][7] = xor_out[35][23][7] + xor_out[36][23][7] + xor_out[37][23][7] + xor_out[38][23][7] + xor_out[39][23][7];
assign sum_out[8][23][7] = xor_out[40][23][7] + xor_out[41][23][7] + xor_out[42][23][7] + xor_out[43][23][7] + xor_out[44][23][7];
assign sum_out[9][23][7] = xor_out[45][23][7] + xor_out[46][23][7] + xor_out[47][23][7] + xor_out[48][23][7] + xor_out[49][23][7];
assign sum_out[10][23][7] = xor_out[50][23][7] + xor_out[51][23][7] + xor_out[52][23][7] + xor_out[53][23][7] + xor_out[54][23][7];
assign sum_out[11][23][7] = xor_out[55][23][7] + xor_out[56][23][7] + xor_out[57][23][7] + xor_out[58][23][7] + xor_out[59][23][7];
assign sum_out[12][23][7] = xor_out[60][23][7] + xor_out[61][23][7] + xor_out[62][23][7] + xor_out[63][23][7] + xor_out[64][23][7];
assign sum_out[13][23][7] = xor_out[65][23][7] + xor_out[66][23][7] + xor_out[67][23][7] + xor_out[68][23][7] + xor_out[69][23][7];
assign sum_out[14][23][7] = xor_out[70][23][7] + xor_out[71][23][7] + xor_out[72][23][7] + xor_out[73][23][7] + xor_out[74][23][7];
assign sum_out[15][23][7] = xor_out[75][23][7] + xor_out[76][23][7] + xor_out[77][23][7] + xor_out[78][23][7] + xor_out[79][23][7];
assign sum_out[16][23][7] = xor_out[80][23][7] + xor_out[81][23][7] + xor_out[82][23][7] + xor_out[83][23][7] + xor_out[84][23][7];
assign sum_out[17][23][7] = xor_out[85][23][7] + xor_out[86][23][7] + xor_out[87][23][7] + xor_out[88][23][7] + xor_out[89][23][7];
assign sum_out[18][23][7] = xor_out[90][23][7] + xor_out[91][23][7] + xor_out[92][23][7] + xor_out[93][23][7] + xor_out[94][23][7];
assign sum_out[19][23][7] = xor_out[95][23][7] + xor_out[96][23][7] + xor_out[97][23][7] + xor_out[98][23][7] + xor_out[99][23][7];

assign sum_out[0][23][8] = xor_out[0][23][8] + xor_out[1][23][8] + xor_out[2][23][8] + xor_out[3][23][8] + xor_out[4][23][8];
assign sum_out[1][23][8] = xor_out[5][23][8] + xor_out[6][23][8] + xor_out[7][23][8] + xor_out[8][23][8] + xor_out[9][23][8];
assign sum_out[2][23][8] = xor_out[10][23][8] + xor_out[11][23][8] + xor_out[12][23][8] + xor_out[13][23][8] + xor_out[14][23][8];
assign sum_out[3][23][8] = xor_out[15][23][8] + xor_out[16][23][8] + xor_out[17][23][8] + xor_out[18][23][8] + xor_out[19][23][8];
assign sum_out[4][23][8] = xor_out[20][23][8] + xor_out[21][23][8] + xor_out[22][23][8] + xor_out[23][23][8] + xor_out[24][23][8];
assign sum_out[5][23][8] = xor_out[25][23][8] + xor_out[26][23][8] + xor_out[27][23][8] + xor_out[28][23][8] + xor_out[29][23][8];
assign sum_out[6][23][8] = xor_out[30][23][8] + xor_out[31][23][8] + xor_out[32][23][8] + xor_out[33][23][8] + xor_out[34][23][8];
assign sum_out[7][23][8] = xor_out[35][23][8] + xor_out[36][23][8] + xor_out[37][23][8] + xor_out[38][23][8] + xor_out[39][23][8];
assign sum_out[8][23][8] = xor_out[40][23][8] + xor_out[41][23][8] + xor_out[42][23][8] + xor_out[43][23][8] + xor_out[44][23][8];
assign sum_out[9][23][8] = xor_out[45][23][8] + xor_out[46][23][8] + xor_out[47][23][8] + xor_out[48][23][8] + xor_out[49][23][8];
assign sum_out[10][23][8] = xor_out[50][23][8] + xor_out[51][23][8] + xor_out[52][23][8] + xor_out[53][23][8] + xor_out[54][23][8];
assign sum_out[11][23][8] = xor_out[55][23][8] + xor_out[56][23][8] + xor_out[57][23][8] + xor_out[58][23][8] + xor_out[59][23][8];
assign sum_out[12][23][8] = xor_out[60][23][8] + xor_out[61][23][8] + xor_out[62][23][8] + xor_out[63][23][8] + xor_out[64][23][8];
assign sum_out[13][23][8] = xor_out[65][23][8] + xor_out[66][23][8] + xor_out[67][23][8] + xor_out[68][23][8] + xor_out[69][23][8];
assign sum_out[14][23][8] = xor_out[70][23][8] + xor_out[71][23][8] + xor_out[72][23][8] + xor_out[73][23][8] + xor_out[74][23][8];
assign sum_out[15][23][8] = xor_out[75][23][8] + xor_out[76][23][8] + xor_out[77][23][8] + xor_out[78][23][8] + xor_out[79][23][8];
assign sum_out[16][23][8] = xor_out[80][23][8] + xor_out[81][23][8] + xor_out[82][23][8] + xor_out[83][23][8] + xor_out[84][23][8];
assign sum_out[17][23][8] = xor_out[85][23][8] + xor_out[86][23][8] + xor_out[87][23][8] + xor_out[88][23][8] + xor_out[89][23][8];
assign sum_out[18][23][8] = xor_out[90][23][8] + xor_out[91][23][8] + xor_out[92][23][8] + xor_out[93][23][8] + xor_out[94][23][8];
assign sum_out[19][23][8] = xor_out[95][23][8] + xor_out[96][23][8] + xor_out[97][23][8] + xor_out[98][23][8] + xor_out[99][23][8];

assign sum_out[0][23][9] = xor_out[0][23][9] + xor_out[1][23][9] + xor_out[2][23][9] + xor_out[3][23][9] + xor_out[4][23][9];
assign sum_out[1][23][9] = xor_out[5][23][9] + xor_out[6][23][9] + xor_out[7][23][9] + xor_out[8][23][9] + xor_out[9][23][9];
assign sum_out[2][23][9] = xor_out[10][23][9] + xor_out[11][23][9] + xor_out[12][23][9] + xor_out[13][23][9] + xor_out[14][23][9];
assign sum_out[3][23][9] = xor_out[15][23][9] + xor_out[16][23][9] + xor_out[17][23][9] + xor_out[18][23][9] + xor_out[19][23][9];
assign sum_out[4][23][9] = xor_out[20][23][9] + xor_out[21][23][9] + xor_out[22][23][9] + xor_out[23][23][9] + xor_out[24][23][9];
assign sum_out[5][23][9] = xor_out[25][23][9] + xor_out[26][23][9] + xor_out[27][23][9] + xor_out[28][23][9] + xor_out[29][23][9];
assign sum_out[6][23][9] = xor_out[30][23][9] + xor_out[31][23][9] + xor_out[32][23][9] + xor_out[33][23][9] + xor_out[34][23][9];
assign sum_out[7][23][9] = xor_out[35][23][9] + xor_out[36][23][9] + xor_out[37][23][9] + xor_out[38][23][9] + xor_out[39][23][9];
assign sum_out[8][23][9] = xor_out[40][23][9] + xor_out[41][23][9] + xor_out[42][23][9] + xor_out[43][23][9] + xor_out[44][23][9];
assign sum_out[9][23][9] = xor_out[45][23][9] + xor_out[46][23][9] + xor_out[47][23][9] + xor_out[48][23][9] + xor_out[49][23][9];
assign sum_out[10][23][9] = xor_out[50][23][9] + xor_out[51][23][9] + xor_out[52][23][9] + xor_out[53][23][9] + xor_out[54][23][9];
assign sum_out[11][23][9] = xor_out[55][23][9] + xor_out[56][23][9] + xor_out[57][23][9] + xor_out[58][23][9] + xor_out[59][23][9];
assign sum_out[12][23][9] = xor_out[60][23][9] + xor_out[61][23][9] + xor_out[62][23][9] + xor_out[63][23][9] + xor_out[64][23][9];
assign sum_out[13][23][9] = xor_out[65][23][9] + xor_out[66][23][9] + xor_out[67][23][9] + xor_out[68][23][9] + xor_out[69][23][9];
assign sum_out[14][23][9] = xor_out[70][23][9] + xor_out[71][23][9] + xor_out[72][23][9] + xor_out[73][23][9] + xor_out[74][23][9];
assign sum_out[15][23][9] = xor_out[75][23][9] + xor_out[76][23][9] + xor_out[77][23][9] + xor_out[78][23][9] + xor_out[79][23][9];
assign sum_out[16][23][9] = xor_out[80][23][9] + xor_out[81][23][9] + xor_out[82][23][9] + xor_out[83][23][9] + xor_out[84][23][9];
assign sum_out[17][23][9] = xor_out[85][23][9] + xor_out[86][23][9] + xor_out[87][23][9] + xor_out[88][23][9] + xor_out[89][23][9];
assign sum_out[18][23][9] = xor_out[90][23][9] + xor_out[91][23][9] + xor_out[92][23][9] + xor_out[93][23][9] + xor_out[94][23][9];
assign sum_out[19][23][9] = xor_out[95][23][9] + xor_out[96][23][9] + xor_out[97][23][9] + xor_out[98][23][9] + xor_out[99][23][9];

assign sum_out[0][23][10] = xor_out[0][23][10] + xor_out[1][23][10] + xor_out[2][23][10] + xor_out[3][23][10] + xor_out[4][23][10];
assign sum_out[1][23][10] = xor_out[5][23][10] + xor_out[6][23][10] + xor_out[7][23][10] + xor_out[8][23][10] + xor_out[9][23][10];
assign sum_out[2][23][10] = xor_out[10][23][10] + xor_out[11][23][10] + xor_out[12][23][10] + xor_out[13][23][10] + xor_out[14][23][10];
assign sum_out[3][23][10] = xor_out[15][23][10] + xor_out[16][23][10] + xor_out[17][23][10] + xor_out[18][23][10] + xor_out[19][23][10];
assign sum_out[4][23][10] = xor_out[20][23][10] + xor_out[21][23][10] + xor_out[22][23][10] + xor_out[23][23][10] + xor_out[24][23][10];
assign sum_out[5][23][10] = xor_out[25][23][10] + xor_out[26][23][10] + xor_out[27][23][10] + xor_out[28][23][10] + xor_out[29][23][10];
assign sum_out[6][23][10] = xor_out[30][23][10] + xor_out[31][23][10] + xor_out[32][23][10] + xor_out[33][23][10] + xor_out[34][23][10];
assign sum_out[7][23][10] = xor_out[35][23][10] + xor_out[36][23][10] + xor_out[37][23][10] + xor_out[38][23][10] + xor_out[39][23][10];
assign sum_out[8][23][10] = xor_out[40][23][10] + xor_out[41][23][10] + xor_out[42][23][10] + xor_out[43][23][10] + xor_out[44][23][10];
assign sum_out[9][23][10] = xor_out[45][23][10] + xor_out[46][23][10] + xor_out[47][23][10] + xor_out[48][23][10] + xor_out[49][23][10];
assign sum_out[10][23][10] = xor_out[50][23][10] + xor_out[51][23][10] + xor_out[52][23][10] + xor_out[53][23][10] + xor_out[54][23][10];
assign sum_out[11][23][10] = xor_out[55][23][10] + xor_out[56][23][10] + xor_out[57][23][10] + xor_out[58][23][10] + xor_out[59][23][10];
assign sum_out[12][23][10] = xor_out[60][23][10] + xor_out[61][23][10] + xor_out[62][23][10] + xor_out[63][23][10] + xor_out[64][23][10];
assign sum_out[13][23][10] = xor_out[65][23][10] + xor_out[66][23][10] + xor_out[67][23][10] + xor_out[68][23][10] + xor_out[69][23][10];
assign sum_out[14][23][10] = xor_out[70][23][10] + xor_out[71][23][10] + xor_out[72][23][10] + xor_out[73][23][10] + xor_out[74][23][10];
assign sum_out[15][23][10] = xor_out[75][23][10] + xor_out[76][23][10] + xor_out[77][23][10] + xor_out[78][23][10] + xor_out[79][23][10];
assign sum_out[16][23][10] = xor_out[80][23][10] + xor_out[81][23][10] + xor_out[82][23][10] + xor_out[83][23][10] + xor_out[84][23][10];
assign sum_out[17][23][10] = xor_out[85][23][10] + xor_out[86][23][10] + xor_out[87][23][10] + xor_out[88][23][10] + xor_out[89][23][10];
assign sum_out[18][23][10] = xor_out[90][23][10] + xor_out[91][23][10] + xor_out[92][23][10] + xor_out[93][23][10] + xor_out[94][23][10];
assign sum_out[19][23][10] = xor_out[95][23][10] + xor_out[96][23][10] + xor_out[97][23][10] + xor_out[98][23][10] + xor_out[99][23][10];

assign sum_out[0][23][11] = xor_out[0][23][11] + xor_out[1][23][11] + xor_out[2][23][11] + xor_out[3][23][11] + xor_out[4][23][11];
assign sum_out[1][23][11] = xor_out[5][23][11] + xor_out[6][23][11] + xor_out[7][23][11] + xor_out[8][23][11] + xor_out[9][23][11];
assign sum_out[2][23][11] = xor_out[10][23][11] + xor_out[11][23][11] + xor_out[12][23][11] + xor_out[13][23][11] + xor_out[14][23][11];
assign sum_out[3][23][11] = xor_out[15][23][11] + xor_out[16][23][11] + xor_out[17][23][11] + xor_out[18][23][11] + xor_out[19][23][11];
assign sum_out[4][23][11] = xor_out[20][23][11] + xor_out[21][23][11] + xor_out[22][23][11] + xor_out[23][23][11] + xor_out[24][23][11];
assign sum_out[5][23][11] = xor_out[25][23][11] + xor_out[26][23][11] + xor_out[27][23][11] + xor_out[28][23][11] + xor_out[29][23][11];
assign sum_out[6][23][11] = xor_out[30][23][11] + xor_out[31][23][11] + xor_out[32][23][11] + xor_out[33][23][11] + xor_out[34][23][11];
assign sum_out[7][23][11] = xor_out[35][23][11] + xor_out[36][23][11] + xor_out[37][23][11] + xor_out[38][23][11] + xor_out[39][23][11];
assign sum_out[8][23][11] = xor_out[40][23][11] + xor_out[41][23][11] + xor_out[42][23][11] + xor_out[43][23][11] + xor_out[44][23][11];
assign sum_out[9][23][11] = xor_out[45][23][11] + xor_out[46][23][11] + xor_out[47][23][11] + xor_out[48][23][11] + xor_out[49][23][11];
assign sum_out[10][23][11] = xor_out[50][23][11] + xor_out[51][23][11] + xor_out[52][23][11] + xor_out[53][23][11] + xor_out[54][23][11];
assign sum_out[11][23][11] = xor_out[55][23][11] + xor_out[56][23][11] + xor_out[57][23][11] + xor_out[58][23][11] + xor_out[59][23][11];
assign sum_out[12][23][11] = xor_out[60][23][11] + xor_out[61][23][11] + xor_out[62][23][11] + xor_out[63][23][11] + xor_out[64][23][11];
assign sum_out[13][23][11] = xor_out[65][23][11] + xor_out[66][23][11] + xor_out[67][23][11] + xor_out[68][23][11] + xor_out[69][23][11];
assign sum_out[14][23][11] = xor_out[70][23][11] + xor_out[71][23][11] + xor_out[72][23][11] + xor_out[73][23][11] + xor_out[74][23][11];
assign sum_out[15][23][11] = xor_out[75][23][11] + xor_out[76][23][11] + xor_out[77][23][11] + xor_out[78][23][11] + xor_out[79][23][11];
assign sum_out[16][23][11] = xor_out[80][23][11] + xor_out[81][23][11] + xor_out[82][23][11] + xor_out[83][23][11] + xor_out[84][23][11];
assign sum_out[17][23][11] = xor_out[85][23][11] + xor_out[86][23][11] + xor_out[87][23][11] + xor_out[88][23][11] + xor_out[89][23][11];
assign sum_out[18][23][11] = xor_out[90][23][11] + xor_out[91][23][11] + xor_out[92][23][11] + xor_out[93][23][11] + xor_out[94][23][11];
assign sum_out[19][23][11] = xor_out[95][23][11] + xor_out[96][23][11] + xor_out[97][23][11] + xor_out[98][23][11] + xor_out[99][23][11];

assign sum_out[0][23][12] = xor_out[0][23][12] + xor_out[1][23][12] + xor_out[2][23][12] + xor_out[3][23][12] + xor_out[4][23][12];
assign sum_out[1][23][12] = xor_out[5][23][12] + xor_out[6][23][12] + xor_out[7][23][12] + xor_out[8][23][12] + xor_out[9][23][12];
assign sum_out[2][23][12] = xor_out[10][23][12] + xor_out[11][23][12] + xor_out[12][23][12] + xor_out[13][23][12] + xor_out[14][23][12];
assign sum_out[3][23][12] = xor_out[15][23][12] + xor_out[16][23][12] + xor_out[17][23][12] + xor_out[18][23][12] + xor_out[19][23][12];
assign sum_out[4][23][12] = xor_out[20][23][12] + xor_out[21][23][12] + xor_out[22][23][12] + xor_out[23][23][12] + xor_out[24][23][12];
assign sum_out[5][23][12] = xor_out[25][23][12] + xor_out[26][23][12] + xor_out[27][23][12] + xor_out[28][23][12] + xor_out[29][23][12];
assign sum_out[6][23][12] = xor_out[30][23][12] + xor_out[31][23][12] + xor_out[32][23][12] + xor_out[33][23][12] + xor_out[34][23][12];
assign sum_out[7][23][12] = xor_out[35][23][12] + xor_out[36][23][12] + xor_out[37][23][12] + xor_out[38][23][12] + xor_out[39][23][12];
assign sum_out[8][23][12] = xor_out[40][23][12] + xor_out[41][23][12] + xor_out[42][23][12] + xor_out[43][23][12] + xor_out[44][23][12];
assign sum_out[9][23][12] = xor_out[45][23][12] + xor_out[46][23][12] + xor_out[47][23][12] + xor_out[48][23][12] + xor_out[49][23][12];
assign sum_out[10][23][12] = xor_out[50][23][12] + xor_out[51][23][12] + xor_out[52][23][12] + xor_out[53][23][12] + xor_out[54][23][12];
assign sum_out[11][23][12] = xor_out[55][23][12] + xor_out[56][23][12] + xor_out[57][23][12] + xor_out[58][23][12] + xor_out[59][23][12];
assign sum_out[12][23][12] = xor_out[60][23][12] + xor_out[61][23][12] + xor_out[62][23][12] + xor_out[63][23][12] + xor_out[64][23][12];
assign sum_out[13][23][12] = xor_out[65][23][12] + xor_out[66][23][12] + xor_out[67][23][12] + xor_out[68][23][12] + xor_out[69][23][12];
assign sum_out[14][23][12] = xor_out[70][23][12] + xor_out[71][23][12] + xor_out[72][23][12] + xor_out[73][23][12] + xor_out[74][23][12];
assign sum_out[15][23][12] = xor_out[75][23][12] + xor_out[76][23][12] + xor_out[77][23][12] + xor_out[78][23][12] + xor_out[79][23][12];
assign sum_out[16][23][12] = xor_out[80][23][12] + xor_out[81][23][12] + xor_out[82][23][12] + xor_out[83][23][12] + xor_out[84][23][12];
assign sum_out[17][23][12] = xor_out[85][23][12] + xor_out[86][23][12] + xor_out[87][23][12] + xor_out[88][23][12] + xor_out[89][23][12];
assign sum_out[18][23][12] = xor_out[90][23][12] + xor_out[91][23][12] + xor_out[92][23][12] + xor_out[93][23][12] + xor_out[94][23][12];
assign sum_out[19][23][12] = xor_out[95][23][12] + xor_out[96][23][12] + xor_out[97][23][12] + xor_out[98][23][12] + xor_out[99][23][12];

assign sum_out[0][23][13] = xor_out[0][23][13] + xor_out[1][23][13] + xor_out[2][23][13] + xor_out[3][23][13] + xor_out[4][23][13];
assign sum_out[1][23][13] = xor_out[5][23][13] + xor_out[6][23][13] + xor_out[7][23][13] + xor_out[8][23][13] + xor_out[9][23][13];
assign sum_out[2][23][13] = xor_out[10][23][13] + xor_out[11][23][13] + xor_out[12][23][13] + xor_out[13][23][13] + xor_out[14][23][13];
assign sum_out[3][23][13] = xor_out[15][23][13] + xor_out[16][23][13] + xor_out[17][23][13] + xor_out[18][23][13] + xor_out[19][23][13];
assign sum_out[4][23][13] = xor_out[20][23][13] + xor_out[21][23][13] + xor_out[22][23][13] + xor_out[23][23][13] + xor_out[24][23][13];
assign sum_out[5][23][13] = xor_out[25][23][13] + xor_out[26][23][13] + xor_out[27][23][13] + xor_out[28][23][13] + xor_out[29][23][13];
assign sum_out[6][23][13] = xor_out[30][23][13] + xor_out[31][23][13] + xor_out[32][23][13] + xor_out[33][23][13] + xor_out[34][23][13];
assign sum_out[7][23][13] = xor_out[35][23][13] + xor_out[36][23][13] + xor_out[37][23][13] + xor_out[38][23][13] + xor_out[39][23][13];
assign sum_out[8][23][13] = xor_out[40][23][13] + xor_out[41][23][13] + xor_out[42][23][13] + xor_out[43][23][13] + xor_out[44][23][13];
assign sum_out[9][23][13] = xor_out[45][23][13] + xor_out[46][23][13] + xor_out[47][23][13] + xor_out[48][23][13] + xor_out[49][23][13];
assign sum_out[10][23][13] = xor_out[50][23][13] + xor_out[51][23][13] + xor_out[52][23][13] + xor_out[53][23][13] + xor_out[54][23][13];
assign sum_out[11][23][13] = xor_out[55][23][13] + xor_out[56][23][13] + xor_out[57][23][13] + xor_out[58][23][13] + xor_out[59][23][13];
assign sum_out[12][23][13] = xor_out[60][23][13] + xor_out[61][23][13] + xor_out[62][23][13] + xor_out[63][23][13] + xor_out[64][23][13];
assign sum_out[13][23][13] = xor_out[65][23][13] + xor_out[66][23][13] + xor_out[67][23][13] + xor_out[68][23][13] + xor_out[69][23][13];
assign sum_out[14][23][13] = xor_out[70][23][13] + xor_out[71][23][13] + xor_out[72][23][13] + xor_out[73][23][13] + xor_out[74][23][13];
assign sum_out[15][23][13] = xor_out[75][23][13] + xor_out[76][23][13] + xor_out[77][23][13] + xor_out[78][23][13] + xor_out[79][23][13];
assign sum_out[16][23][13] = xor_out[80][23][13] + xor_out[81][23][13] + xor_out[82][23][13] + xor_out[83][23][13] + xor_out[84][23][13];
assign sum_out[17][23][13] = xor_out[85][23][13] + xor_out[86][23][13] + xor_out[87][23][13] + xor_out[88][23][13] + xor_out[89][23][13];
assign sum_out[18][23][13] = xor_out[90][23][13] + xor_out[91][23][13] + xor_out[92][23][13] + xor_out[93][23][13] + xor_out[94][23][13];
assign sum_out[19][23][13] = xor_out[95][23][13] + xor_out[96][23][13] + xor_out[97][23][13] + xor_out[98][23][13] + xor_out[99][23][13];

assign sum_out[0][23][14] = xor_out[0][23][14] + xor_out[1][23][14] + xor_out[2][23][14] + xor_out[3][23][14] + xor_out[4][23][14];
assign sum_out[1][23][14] = xor_out[5][23][14] + xor_out[6][23][14] + xor_out[7][23][14] + xor_out[8][23][14] + xor_out[9][23][14];
assign sum_out[2][23][14] = xor_out[10][23][14] + xor_out[11][23][14] + xor_out[12][23][14] + xor_out[13][23][14] + xor_out[14][23][14];
assign sum_out[3][23][14] = xor_out[15][23][14] + xor_out[16][23][14] + xor_out[17][23][14] + xor_out[18][23][14] + xor_out[19][23][14];
assign sum_out[4][23][14] = xor_out[20][23][14] + xor_out[21][23][14] + xor_out[22][23][14] + xor_out[23][23][14] + xor_out[24][23][14];
assign sum_out[5][23][14] = xor_out[25][23][14] + xor_out[26][23][14] + xor_out[27][23][14] + xor_out[28][23][14] + xor_out[29][23][14];
assign sum_out[6][23][14] = xor_out[30][23][14] + xor_out[31][23][14] + xor_out[32][23][14] + xor_out[33][23][14] + xor_out[34][23][14];
assign sum_out[7][23][14] = xor_out[35][23][14] + xor_out[36][23][14] + xor_out[37][23][14] + xor_out[38][23][14] + xor_out[39][23][14];
assign sum_out[8][23][14] = xor_out[40][23][14] + xor_out[41][23][14] + xor_out[42][23][14] + xor_out[43][23][14] + xor_out[44][23][14];
assign sum_out[9][23][14] = xor_out[45][23][14] + xor_out[46][23][14] + xor_out[47][23][14] + xor_out[48][23][14] + xor_out[49][23][14];
assign sum_out[10][23][14] = xor_out[50][23][14] + xor_out[51][23][14] + xor_out[52][23][14] + xor_out[53][23][14] + xor_out[54][23][14];
assign sum_out[11][23][14] = xor_out[55][23][14] + xor_out[56][23][14] + xor_out[57][23][14] + xor_out[58][23][14] + xor_out[59][23][14];
assign sum_out[12][23][14] = xor_out[60][23][14] + xor_out[61][23][14] + xor_out[62][23][14] + xor_out[63][23][14] + xor_out[64][23][14];
assign sum_out[13][23][14] = xor_out[65][23][14] + xor_out[66][23][14] + xor_out[67][23][14] + xor_out[68][23][14] + xor_out[69][23][14];
assign sum_out[14][23][14] = xor_out[70][23][14] + xor_out[71][23][14] + xor_out[72][23][14] + xor_out[73][23][14] + xor_out[74][23][14];
assign sum_out[15][23][14] = xor_out[75][23][14] + xor_out[76][23][14] + xor_out[77][23][14] + xor_out[78][23][14] + xor_out[79][23][14];
assign sum_out[16][23][14] = xor_out[80][23][14] + xor_out[81][23][14] + xor_out[82][23][14] + xor_out[83][23][14] + xor_out[84][23][14];
assign sum_out[17][23][14] = xor_out[85][23][14] + xor_out[86][23][14] + xor_out[87][23][14] + xor_out[88][23][14] + xor_out[89][23][14];
assign sum_out[18][23][14] = xor_out[90][23][14] + xor_out[91][23][14] + xor_out[92][23][14] + xor_out[93][23][14] + xor_out[94][23][14];
assign sum_out[19][23][14] = xor_out[95][23][14] + xor_out[96][23][14] + xor_out[97][23][14] + xor_out[98][23][14] + xor_out[99][23][14];

assign sum_out[0][23][15] = xor_out[0][23][15] + xor_out[1][23][15] + xor_out[2][23][15] + xor_out[3][23][15] + xor_out[4][23][15];
assign sum_out[1][23][15] = xor_out[5][23][15] + xor_out[6][23][15] + xor_out[7][23][15] + xor_out[8][23][15] + xor_out[9][23][15];
assign sum_out[2][23][15] = xor_out[10][23][15] + xor_out[11][23][15] + xor_out[12][23][15] + xor_out[13][23][15] + xor_out[14][23][15];
assign sum_out[3][23][15] = xor_out[15][23][15] + xor_out[16][23][15] + xor_out[17][23][15] + xor_out[18][23][15] + xor_out[19][23][15];
assign sum_out[4][23][15] = xor_out[20][23][15] + xor_out[21][23][15] + xor_out[22][23][15] + xor_out[23][23][15] + xor_out[24][23][15];
assign sum_out[5][23][15] = xor_out[25][23][15] + xor_out[26][23][15] + xor_out[27][23][15] + xor_out[28][23][15] + xor_out[29][23][15];
assign sum_out[6][23][15] = xor_out[30][23][15] + xor_out[31][23][15] + xor_out[32][23][15] + xor_out[33][23][15] + xor_out[34][23][15];
assign sum_out[7][23][15] = xor_out[35][23][15] + xor_out[36][23][15] + xor_out[37][23][15] + xor_out[38][23][15] + xor_out[39][23][15];
assign sum_out[8][23][15] = xor_out[40][23][15] + xor_out[41][23][15] + xor_out[42][23][15] + xor_out[43][23][15] + xor_out[44][23][15];
assign sum_out[9][23][15] = xor_out[45][23][15] + xor_out[46][23][15] + xor_out[47][23][15] + xor_out[48][23][15] + xor_out[49][23][15];
assign sum_out[10][23][15] = xor_out[50][23][15] + xor_out[51][23][15] + xor_out[52][23][15] + xor_out[53][23][15] + xor_out[54][23][15];
assign sum_out[11][23][15] = xor_out[55][23][15] + xor_out[56][23][15] + xor_out[57][23][15] + xor_out[58][23][15] + xor_out[59][23][15];
assign sum_out[12][23][15] = xor_out[60][23][15] + xor_out[61][23][15] + xor_out[62][23][15] + xor_out[63][23][15] + xor_out[64][23][15];
assign sum_out[13][23][15] = xor_out[65][23][15] + xor_out[66][23][15] + xor_out[67][23][15] + xor_out[68][23][15] + xor_out[69][23][15];
assign sum_out[14][23][15] = xor_out[70][23][15] + xor_out[71][23][15] + xor_out[72][23][15] + xor_out[73][23][15] + xor_out[74][23][15];
assign sum_out[15][23][15] = xor_out[75][23][15] + xor_out[76][23][15] + xor_out[77][23][15] + xor_out[78][23][15] + xor_out[79][23][15];
assign sum_out[16][23][15] = xor_out[80][23][15] + xor_out[81][23][15] + xor_out[82][23][15] + xor_out[83][23][15] + xor_out[84][23][15];
assign sum_out[17][23][15] = xor_out[85][23][15] + xor_out[86][23][15] + xor_out[87][23][15] + xor_out[88][23][15] + xor_out[89][23][15];
assign sum_out[18][23][15] = xor_out[90][23][15] + xor_out[91][23][15] + xor_out[92][23][15] + xor_out[93][23][15] + xor_out[94][23][15];
assign sum_out[19][23][15] = xor_out[95][23][15] + xor_out[96][23][15] + xor_out[97][23][15] + xor_out[98][23][15] + xor_out[99][23][15];

assign sum_out[0][23][16] = xor_out[0][23][16] + xor_out[1][23][16] + xor_out[2][23][16] + xor_out[3][23][16] + xor_out[4][23][16];
assign sum_out[1][23][16] = xor_out[5][23][16] + xor_out[6][23][16] + xor_out[7][23][16] + xor_out[8][23][16] + xor_out[9][23][16];
assign sum_out[2][23][16] = xor_out[10][23][16] + xor_out[11][23][16] + xor_out[12][23][16] + xor_out[13][23][16] + xor_out[14][23][16];
assign sum_out[3][23][16] = xor_out[15][23][16] + xor_out[16][23][16] + xor_out[17][23][16] + xor_out[18][23][16] + xor_out[19][23][16];
assign sum_out[4][23][16] = xor_out[20][23][16] + xor_out[21][23][16] + xor_out[22][23][16] + xor_out[23][23][16] + xor_out[24][23][16];
assign sum_out[5][23][16] = xor_out[25][23][16] + xor_out[26][23][16] + xor_out[27][23][16] + xor_out[28][23][16] + xor_out[29][23][16];
assign sum_out[6][23][16] = xor_out[30][23][16] + xor_out[31][23][16] + xor_out[32][23][16] + xor_out[33][23][16] + xor_out[34][23][16];
assign sum_out[7][23][16] = xor_out[35][23][16] + xor_out[36][23][16] + xor_out[37][23][16] + xor_out[38][23][16] + xor_out[39][23][16];
assign sum_out[8][23][16] = xor_out[40][23][16] + xor_out[41][23][16] + xor_out[42][23][16] + xor_out[43][23][16] + xor_out[44][23][16];
assign sum_out[9][23][16] = xor_out[45][23][16] + xor_out[46][23][16] + xor_out[47][23][16] + xor_out[48][23][16] + xor_out[49][23][16];
assign sum_out[10][23][16] = xor_out[50][23][16] + xor_out[51][23][16] + xor_out[52][23][16] + xor_out[53][23][16] + xor_out[54][23][16];
assign sum_out[11][23][16] = xor_out[55][23][16] + xor_out[56][23][16] + xor_out[57][23][16] + xor_out[58][23][16] + xor_out[59][23][16];
assign sum_out[12][23][16] = xor_out[60][23][16] + xor_out[61][23][16] + xor_out[62][23][16] + xor_out[63][23][16] + xor_out[64][23][16];
assign sum_out[13][23][16] = xor_out[65][23][16] + xor_out[66][23][16] + xor_out[67][23][16] + xor_out[68][23][16] + xor_out[69][23][16];
assign sum_out[14][23][16] = xor_out[70][23][16] + xor_out[71][23][16] + xor_out[72][23][16] + xor_out[73][23][16] + xor_out[74][23][16];
assign sum_out[15][23][16] = xor_out[75][23][16] + xor_out[76][23][16] + xor_out[77][23][16] + xor_out[78][23][16] + xor_out[79][23][16];
assign sum_out[16][23][16] = xor_out[80][23][16] + xor_out[81][23][16] + xor_out[82][23][16] + xor_out[83][23][16] + xor_out[84][23][16];
assign sum_out[17][23][16] = xor_out[85][23][16] + xor_out[86][23][16] + xor_out[87][23][16] + xor_out[88][23][16] + xor_out[89][23][16];
assign sum_out[18][23][16] = xor_out[90][23][16] + xor_out[91][23][16] + xor_out[92][23][16] + xor_out[93][23][16] + xor_out[94][23][16];
assign sum_out[19][23][16] = xor_out[95][23][16] + xor_out[96][23][16] + xor_out[97][23][16] + xor_out[98][23][16] + xor_out[99][23][16];

assign sum_out[0][23][17] = xor_out[0][23][17] + xor_out[1][23][17] + xor_out[2][23][17] + xor_out[3][23][17] + xor_out[4][23][17];
assign sum_out[1][23][17] = xor_out[5][23][17] + xor_out[6][23][17] + xor_out[7][23][17] + xor_out[8][23][17] + xor_out[9][23][17];
assign sum_out[2][23][17] = xor_out[10][23][17] + xor_out[11][23][17] + xor_out[12][23][17] + xor_out[13][23][17] + xor_out[14][23][17];
assign sum_out[3][23][17] = xor_out[15][23][17] + xor_out[16][23][17] + xor_out[17][23][17] + xor_out[18][23][17] + xor_out[19][23][17];
assign sum_out[4][23][17] = xor_out[20][23][17] + xor_out[21][23][17] + xor_out[22][23][17] + xor_out[23][23][17] + xor_out[24][23][17];
assign sum_out[5][23][17] = xor_out[25][23][17] + xor_out[26][23][17] + xor_out[27][23][17] + xor_out[28][23][17] + xor_out[29][23][17];
assign sum_out[6][23][17] = xor_out[30][23][17] + xor_out[31][23][17] + xor_out[32][23][17] + xor_out[33][23][17] + xor_out[34][23][17];
assign sum_out[7][23][17] = xor_out[35][23][17] + xor_out[36][23][17] + xor_out[37][23][17] + xor_out[38][23][17] + xor_out[39][23][17];
assign sum_out[8][23][17] = xor_out[40][23][17] + xor_out[41][23][17] + xor_out[42][23][17] + xor_out[43][23][17] + xor_out[44][23][17];
assign sum_out[9][23][17] = xor_out[45][23][17] + xor_out[46][23][17] + xor_out[47][23][17] + xor_out[48][23][17] + xor_out[49][23][17];
assign sum_out[10][23][17] = xor_out[50][23][17] + xor_out[51][23][17] + xor_out[52][23][17] + xor_out[53][23][17] + xor_out[54][23][17];
assign sum_out[11][23][17] = xor_out[55][23][17] + xor_out[56][23][17] + xor_out[57][23][17] + xor_out[58][23][17] + xor_out[59][23][17];
assign sum_out[12][23][17] = xor_out[60][23][17] + xor_out[61][23][17] + xor_out[62][23][17] + xor_out[63][23][17] + xor_out[64][23][17];
assign sum_out[13][23][17] = xor_out[65][23][17] + xor_out[66][23][17] + xor_out[67][23][17] + xor_out[68][23][17] + xor_out[69][23][17];
assign sum_out[14][23][17] = xor_out[70][23][17] + xor_out[71][23][17] + xor_out[72][23][17] + xor_out[73][23][17] + xor_out[74][23][17];
assign sum_out[15][23][17] = xor_out[75][23][17] + xor_out[76][23][17] + xor_out[77][23][17] + xor_out[78][23][17] + xor_out[79][23][17];
assign sum_out[16][23][17] = xor_out[80][23][17] + xor_out[81][23][17] + xor_out[82][23][17] + xor_out[83][23][17] + xor_out[84][23][17];
assign sum_out[17][23][17] = xor_out[85][23][17] + xor_out[86][23][17] + xor_out[87][23][17] + xor_out[88][23][17] + xor_out[89][23][17];
assign sum_out[18][23][17] = xor_out[90][23][17] + xor_out[91][23][17] + xor_out[92][23][17] + xor_out[93][23][17] + xor_out[94][23][17];
assign sum_out[19][23][17] = xor_out[95][23][17] + xor_out[96][23][17] + xor_out[97][23][17] + xor_out[98][23][17] + xor_out[99][23][17];

assign sum_out[0][23][18] = xor_out[0][23][18] + xor_out[1][23][18] + xor_out[2][23][18] + xor_out[3][23][18] + xor_out[4][23][18];
assign sum_out[1][23][18] = xor_out[5][23][18] + xor_out[6][23][18] + xor_out[7][23][18] + xor_out[8][23][18] + xor_out[9][23][18];
assign sum_out[2][23][18] = xor_out[10][23][18] + xor_out[11][23][18] + xor_out[12][23][18] + xor_out[13][23][18] + xor_out[14][23][18];
assign sum_out[3][23][18] = xor_out[15][23][18] + xor_out[16][23][18] + xor_out[17][23][18] + xor_out[18][23][18] + xor_out[19][23][18];
assign sum_out[4][23][18] = xor_out[20][23][18] + xor_out[21][23][18] + xor_out[22][23][18] + xor_out[23][23][18] + xor_out[24][23][18];
assign sum_out[5][23][18] = xor_out[25][23][18] + xor_out[26][23][18] + xor_out[27][23][18] + xor_out[28][23][18] + xor_out[29][23][18];
assign sum_out[6][23][18] = xor_out[30][23][18] + xor_out[31][23][18] + xor_out[32][23][18] + xor_out[33][23][18] + xor_out[34][23][18];
assign sum_out[7][23][18] = xor_out[35][23][18] + xor_out[36][23][18] + xor_out[37][23][18] + xor_out[38][23][18] + xor_out[39][23][18];
assign sum_out[8][23][18] = xor_out[40][23][18] + xor_out[41][23][18] + xor_out[42][23][18] + xor_out[43][23][18] + xor_out[44][23][18];
assign sum_out[9][23][18] = xor_out[45][23][18] + xor_out[46][23][18] + xor_out[47][23][18] + xor_out[48][23][18] + xor_out[49][23][18];
assign sum_out[10][23][18] = xor_out[50][23][18] + xor_out[51][23][18] + xor_out[52][23][18] + xor_out[53][23][18] + xor_out[54][23][18];
assign sum_out[11][23][18] = xor_out[55][23][18] + xor_out[56][23][18] + xor_out[57][23][18] + xor_out[58][23][18] + xor_out[59][23][18];
assign sum_out[12][23][18] = xor_out[60][23][18] + xor_out[61][23][18] + xor_out[62][23][18] + xor_out[63][23][18] + xor_out[64][23][18];
assign sum_out[13][23][18] = xor_out[65][23][18] + xor_out[66][23][18] + xor_out[67][23][18] + xor_out[68][23][18] + xor_out[69][23][18];
assign sum_out[14][23][18] = xor_out[70][23][18] + xor_out[71][23][18] + xor_out[72][23][18] + xor_out[73][23][18] + xor_out[74][23][18];
assign sum_out[15][23][18] = xor_out[75][23][18] + xor_out[76][23][18] + xor_out[77][23][18] + xor_out[78][23][18] + xor_out[79][23][18];
assign sum_out[16][23][18] = xor_out[80][23][18] + xor_out[81][23][18] + xor_out[82][23][18] + xor_out[83][23][18] + xor_out[84][23][18];
assign sum_out[17][23][18] = xor_out[85][23][18] + xor_out[86][23][18] + xor_out[87][23][18] + xor_out[88][23][18] + xor_out[89][23][18];
assign sum_out[18][23][18] = xor_out[90][23][18] + xor_out[91][23][18] + xor_out[92][23][18] + xor_out[93][23][18] + xor_out[94][23][18];
assign sum_out[19][23][18] = xor_out[95][23][18] + xor_out[96][23][18] + xor_out[97][23][18] + xor_out[98][23][18] + xor_out[99][23][18];

assign sum_out[0][23][19] = xor_out[0][23][19] + xor_out[1][23][19] + xor_out[2][23][19] + xor_out[3][23][19] + xor_out[4][23][19];
assign sum_out[1][23][19] = xor_out[5][23][19] + xor_out[6][23][19] + xor_out[7][23][19] + xor_out[8][23][19] + xor_out[9][23][19];
assign sum_out[2][23][19] = xor_out[10][23][19] + xor_out[11][23][19] + xor_out[12][23][19] + xor_out[13][23][19] + xor_out[14][23][19];
assign sum_out[3][23][19] = xor_out[15][23][19] + xor_out[16][23][19] + xor_out[17][23][19] + xor_out[18][23][19] + xor_out[19][23][19];
assign sum_out[4][23][19] = xor_out[20][23][19] + xor_out[21][23][19] + xor_out[22][23][19] + xor_out[23][23][19] + xor_out[24][23][19];
assign sum_out[5][23][19] = xor_out[25][23][19] + xor_out[26][23][19] + xor_out[27][23][19] + xor_out[28][23][19] + xor_out[29][23][19];
assign sum_out[6][23][19] = xor_out[30][23][19] + xor_out[31][23][19] + xor_out[32][23][19] + xor_out[33][23][19] + xor_out[34][23][19];
assign sum_out[7][23][19] = xor_out[35][23][19] + xor_out[36][23][19] + xor_out[37][23][19] + xor_out[38][23][19] + xor_out[39][23][19];
assign sum_out[8][23][19] = xor_out[40][23][19] + xor_out[41][23][19] + xor_out[42][23][19] + xor_out[43][23][19] + xor_out[44][23][19];
assign sum_out[9][23][19] = xor_out[45][23][19] + xor_out[46][23][19] + xor_out[47][23][19] + xor_out[48][23][19] + xor_out[49][23][19];
assign sum_out[10][23][19] = xor_out[50][23][19] + xor_out[51][23][19] + xor_out[52][23][19] + xor_out[53][23][19] + xor_out[54][23][19];
assign sum_out[11][23][19] = xor_out[55][23][19] + xor_out[56][23][19] + xor_out[57][23][19] + xor_out[58][23][19] + xor_out[59][23][19];
assign sum_out[12][23][19] = xor_out[60][23][19] + xor_out[61][23][19] + xor_out[62][23][19] + xor_out[63][23][19] + xor_out[64][23][19];
assign sum_out[13][23][19] = xor_out[65][23][19] + xor_out[66][23][19] + xor_out[67][23][19] + xor_out[68][23][19] + xor_out[69][23][19];
assign sum_out[14][23][19] = xor_out[70][23][19] + xor_out[71][23][19] + xor_out[72][23][19] + xor_out[73][23][19] + xor_out[74][23][19];
assign sum_out[15][23][19] = xor_out[75][23][19] + xor_out[76][23][19] + xor_out[77][23][19] + xor_out[78][23][19] + xor_out[79][23][19];
assign sum_out[16][23][19] = xor_out[80][23][19] + xor_out[81][23][19] + xor_out[82][23][19] + xor_out[83][23][19] + xor_out[84][23][19];
assign sum_out[17][23][19] = xor_out[85][23][19] + xor_out[86][23][19] + xor_out[87][23][19] + xor_out[88][23][19] + xor_out[89][23][19];
assign sum_out[18][23][19] = xor_out[90][23][19] + xor_out[91][23][19] + xor_out[92][23][19] + xor_out[93][23][19] + xor_out[94][23][19];
assign sum_out[19][23][19] = xor_out[95][23][19] + xor_out[96][23][19] + xor_out[97][23][19] + xor_out[98][23][19] + xor_out[99][23][19];

assign sum_out[0][23][20] = xor_out[0][23][20] + xor_out[1][23][20] + xor_out[2][23][20] + xor_out[3][23][20] + xor_out[4][23][20];
assign sum_out[1][23][20] = xor_out[5][23][20] + xor_out[6][23][20] + xor_out[7][23][20] + xor_out[8][23][20] + xor_out[9][23][20];
assign sum_out[2][23][20] = xor_out[10][23][20] + xor_out[11][23][20] + xor_out[12][23][20] + xor_out[13][23][20] + xor_out[14][23][20];
assign sum_out[3][23][20] = xor_out[15][23][20] + xor_out[16][23][20] + xor_out[17][23][20] + xor_out[18][23][20] + xor_out[19][23][20];
assign sum_out[4][23][20] = xor_out[20][23][20] + xor_out[21][23][20] + xor_out[22][23][20] + xor_out[23][23][20] + xor_out[24][23][20];
assign sum_out[5][23][20] = xor_out[25][23][20] + xor_out[26][23][20] + xor_out[27][23][20] + xor_out[28][23][20] + xor_out[29][23][20];
assign sum_out[6][23][20] = xor_out[30][23][20] + xor_out[31][23][20] + xor_out[32][23][20] + xor_out[33][23][20] + xor_out[34][23][20];
assign sum_out[7][23][20] = xor_out[35][23][20] + xor_out[36][23][20] + xor_out[37][23][20] + xor_out[38][23][20] + xor_out[39][23][20];
assign sum_out[8][23][20] = xor_out[40][23][20] + xor_out[41][23][20] + xor_out[42][23][20] + xor_out[43][23][20] + xor_out[44][23][20];
assign sum_out[9][23][20] = xor_out[45][23][20] + xor_out[46][23][20] + xor_out[47][23][20] + xor_out[48][23][20] + xor_out[49][23][20];
assign sum_out[10][23][20] = xor_out[50][23][20] + xor_out[51][23][20] + xor_out[52][23][20] + xor_out[53][23][20] + xor_out[54][23][20];
assign sum_out[11][23][20] = xor_out[55][23][20] + xor_out[56][23][20] + xor_out[57][23][20] + xor_out[58][23][20] + xor_out[59][23][20];
assign sum_out[12][23][20] = xor_out[60][23][20] + xor_out[61][23][20] + xor_out[62][23][20] + xor_out[63][23][20] + xor_out[64][23][20];
assign sum_out[13][23][20] = xor_out[65][23][20] + xor_out[66][23][20] + xor_out[67][23][20] + xor_out[68][23][20] + xor_out[69][23][20];
assign sum_out[14][23][20] = xor_out[70][23][20] + xor_out[71][23][20] + xor_out[72][23][20] + xor_out[73][23][20] + xor_out[74][23][20];
assign sum_out[15][23][20] = xor_out[75][23][20] + xor_out[76][23][20] + xor_out[77][23][20] + xor_out[78][23][20] + xor_out[79][23][20];
assign sum_out[16][23][20] = xor_out[80][23][20] + xor_out[81][23][20] + xor_out[82][23][20] + xor_out[83][23][20] + xor_out[84][23][20];
assign sum_out[17][23][20] = xor_out[85][23][20] + xor_out[86][23][20] + xor_out[87][23][20] + xor_out[88][23][20] + xor_out[89][23][20];
assign sum_out[18][23][20] = xor_out[90][23][20] + xor_out[91][23][20] + xor_out[92][23][20] + xor_out[93][23][20] + xor_out[94][23][20];
assign sum_out[19][23][20] = xor_out[95][23][20] + xor_out[96][23][20] + xor_out[97][23][20] + xor_out[98][23][20] + xor_out[99][23][20];

assign sum_out[0][23][21] = xor_out[0][23][21] + xor_out[1][23][21] + xor_out[2][23][21] + xor_out[3][23][21] + xor_out[4][23][21];
assign sum_out[1][23][21] = xor_out[5][23][21] + xor_out[6][23][21] + xor_out[7][23][21] + xor_out[8][23][21] + xor_out[9][23][21];
assign sum_out[2][23][21] = xor_out[10][23][21] + xor_out[11][23][21] + xor_out[12][23][21] + xor_out[13][23][21] + xor_out[14][23][21];
assign sum_out[3][23][21] = xor_out[15][23][21] + xor_out[16][23][21] + xor_out[17][23][21] + xor_out[18][23][21] + xor_out[19][23][21];
assign sum_out[4][23][21] = xor_out[20][23][21] + xor_out[21][23][21] + xor_out[22][23][21] + xor_out[23][23][21] + xor_out[24][23][21];
assign sum_out[5][23][21] = xor_out[25][23][21] + xor_out[26][23][21] + xor_out[27][23][21] + xor_out[28][23][21] + xor_out[29][23][21];
assign sum_out[6][23][21] = xor_out[30][23][21] + xor_out[31][23][21] + xor_out[32][23][21] + xor_out[33][23][21] + xor_out[34][23][21];
assign sum_out[7][23][21] = xor_out[35][23][21] + xor_out[36][23][21] + xor_out[37][23][21] + xor_out[38][23][21] + xor_out[39][23][21];
assign sum_out[8][23][21] = xor_out[40][23][21] + xor_out[41][23][21] + xor_out[42][23][21] + xor_out[43][23][21] + xor_out[44][23][21];
assign sum_out[9][23][21] = xor_out[45][23][21] + xor_out[46][23][21] + xor_out[47][23][21] + xor_out[48][23][21] + xor_out[49][23][21];
assign sum_out[10][23][21] = xor_out[50][23][21] + xor_out[51][23][21] + xor_out[52][23][21] + xor_out[53][23][21] + xor_out[54][23][21];
assign sum_out[11][23][21] = xor_out[55][23][21] + xor_out[56][23][21] + xor_out[57][23][21] + xor_out[58][23][21] + xor_out[59][23][21];
assign sum_out[12][23][21] = xor_out[60][23][21] + xor_out[61][23][21] + xor_out[62][23][21] + xor_out[63][23][21] + xor_out[64][23][21];
assign sum_out[13][23][21] = xor_out[65][23][21] + xor_out[66][23][21] + xor_out[67][23][21] + xor_out[68][23][21] + xor_out[69][23][21];
assign sum_out[14][23][21] = xor_out[70][23][21] + xor_out[71][23][21] + xor_out[72][23][21] + xor_out[73][23][21] + xor_out[74][23][21];
assign sum_out[15][23][21] = xor_out[75][23][21] + xor_out[76][23][21] + xor_out[77][23][21] + xor_out[78][23][21] + xor_out[79][23][21];
assign sum_out[16][23][21] = xor_out[80][23][21] + xor_out[81][23][21] + xor_out[82][23][21] + xor_out[83][23][21] + xor_out[84][23][21];
assign sum_out[17][23][21] = xor_out[85][23][21] + xor_out[86][23][21] + xor_out[87][23][21] + xor_out[88][23][21] + xor_out[89][23][21];
assign sum_out[18][23][21] = xor_out[90][23][21] + xor_out[91][23][21] + xor_out[92][23][21] + xor_out[93][23][21] + xor_out[94][23][21];
assign sum_out[19][23][21] = xor_out[95][23][21] + xor_out[96][23][21] + xor_out[97][23][21] + xor_out[98][23][21] + xor_out[99][23][21];

assign sum_out[0][23][22] = xor_out[0][23][22] + xor_out[1][23][22] + xor_out[2][23][22] + xor_out[3][23][22] + xor_out[4][23][22];
assign sum_out[1][23][22] = xor_out[5][23][22] + xor_out[6][23][22] + xor_out[7][23][22] + xor_out[8][23][22] + xor_out[9][23][22];
assign sum_out[2][23][22] = xor_out[10][23][22] + xor_out[11][23][22] + xor_out[12][23][22] + xor_out[13][23][22] + xor_out[14][23][22];
assign sum_out[3][23][22] = xor_out[15][23][22] + xor_out[16][23][22] + xor_out[17][23][22] + xor_out[18][23][22] + xor_out[19][23][22];
assign sum_out[4][23][22] = xor_out[20][23][22] + xor_out[21][23][22] + xor_out[22][23][22] + xor_out[23][23][22] + xor_out[24][23][22];
assign sum_out[5][23][22] = xor_out[25][23][22] + xor_out[26][23][22] + xor_out[27][23][22] + xor_out[28][23][22] + xor_out[29][23][22];
assign sum_out[6][23][22] = xor_out[30][23][22] + xor_out[31][23][22] + xor_out[32][23][22] + xor_out[33][23][22] + xor_out[34][23][22];
assign sum_out[7][23][22] = xor_out[35][23][22] + xor_out[36][23][22] + xor_out[37][23][22] + xor_out[38][23][22] + xor_out[39][23][22];
assign sum_out[8][23][22] = xor_out[40][23][22] + xor_out[41][23][22] + xor_out[42][23][22] + xor_out[43][23][22] + xor_out[44][23][22];
assign sum_out[9][23][22] = xor_out[45][23][22] + xor_out[46][23][22] + xor_out[47][23][22] + xor_out[48][23][22] + xor_out[49][23][22];
assign sum_out[10][23][22] = xor_out[50][23][22] + xor_out[51][23][22] + xor_out[52][23][22] + xor_out[53][23][22] + xor_out[54][23][22];
assign sum_out[11][23][22] = xor_out[55][23][22] + xor_out[56][23][22] + xor_out[57][23][22] + xor_out[58][23][22] + xor_out[59][23][22];
assign sum_out[12][23][22] = xor_out[60][23][22] + xor_out[61][23][22] + xor_out[62][23][22] + xor_out[63][23][22] + xor_out[64][23][22];
assign sum_out[13][23][22] = xor_out[65][23][22] + xor_out[66][23][22] + xor_out[67][23][22] + xor_out[68][23][22] + xor_out[69][23][22];
assign sum_out[14][23][22] = xor_out[70][23][22] + xor_out[71][23][22] + xor_out[72][23][22] + xor_out[73][23][22] + xor_out[74][23][22];
assign sum_out[15][23][22] = xor_out[75][23][22] + xor_out[76][23][22] + xor_out[77][23][22] + xor_out[78][23][22] + xor_out[79][23][22];
assign sum_out[16][23][22] = xor_out[80][23][22] + xor_out[81][23][22] + xor_out[82][23][22] + xor_out[83][23][22] + xor_out[84][23][22];
assign sum_out[17][23][22] = xor_out[85][23][22] + xor_out[86][23][22] + xor_out[87][23][22] + xor_out[88][23][22] + xor_out[89][23][22];
assign sum_out[18][23][22] = xor_out[90][23][22] + xor_out[91][23][22] + xor_out[92][23][22] + xor_out[93][23][22] + xor_out[94][23][22];
assign sum_out[19][23][22] = xor_out[95][23][22] + xor_out[96][23][22] + xor_out[97][23][22] + xor_out[98][23][22] + xor_out[99][23][22];

assign sum_out[0][23][23] = xor_out[0][23][23] + xor_out[1][23][23] + xor_out[2][23][23] + xor_out[3][23][23] + xor_out[4][23][23];
assign sum_out[1][23][23] = xor_out[5][23][23] + xor_out[6][23][23] + xor_out[7][23][23] + xor_out[8][23][23] + xor_out[9][23][23];
assign sum_out[2][23][23] = xor_out[10][23][23] + xor_out[11][23][23] + xor_out[12][23][23] + xor_out[13][23][23] + xor_out[14][23][23];
assign sum_out[3][23][23] = xor_out[15][23][23] + xor_out[16][23][23] + xor_out[17][23][23] + xor_out[18][23][23] + xor_out[19][23][23];
assign sum_out[4][23][23] = xor_out[20][23][23] + xor_out[21][23][23] + xor_out[22][23][23] + xor_out[23][23][23] + xor_out[24][23][23];
assign sum_out[5][23][23] = xor_out[25][23][23] + xor_out[26][23][23] + xor_out[27][23][23] + xor_out[28][23][23] + xor_out[29][23][23];
assign sum_out[6][23][23] = xor_out[30][23][23] + xor_out[31][23][23] + xor_out[32][23][23] + xor_out[33][23][23] + xor_out[34][23][23];
assign sum_out[7][23][23] = xor_out[35][23][23] + xor_out[36][23][23] + xor_out[37][23][23] + xor_out[38][23][23] + xor_out[39][23][23];
assign sum_out[8][23][23] = xor_out[40][23][23] + xor_out[41][23][23] + xor_out[42][23][23] + xor_out[43][23][23] + xor_out[44][23][23];
assign sum_out[9][23][23] = xor_out[45][23][23] + xor_out[46][23][23] + xor_out[47][23][23] + xor_out[48][23][23] + xor_out[49][23][23];
assign sum_out[10][23][23] = xor_out[50][23][23] + xor_out[51][23][23] + xor_out[52][23][23] + xor_out[53][23][23] + xor_out[54][23][23];
assign sum_out[11][23][23] = xor_out[55][23][23] + xor_out[56][23][23] + xor_out[57][23][23] + xor_out[58][23][23] + xor_out[59][23][23];
assign sum_out[12][23][23] = xor_out[60][23][23] + xor_out[61][23][23] + xor_out[62][23][23] + xor_out[63][23][23] + xor_out[64][23][23];
assign sum_out[13][23][23] = xor_out[65][23][23] + xor_out[66][23][23] + xor_out[67][23][23] + xor_out[68][23][23] + xor_out[69][23][23];
assign sum_out[14][23][23] = xor_out[70][23][23] + xor_out[71][23][23] + xor_out[72][23][23] + xor_out[73][23][23] + xor_out[74][23][23];
assign sum_out[15][23][23] = xor_out[75][23][23] + xor_out[76][23][23] + xor_out[77][23][23] + xor_out[78][23][23] + xor_out[79][23][23];
assign sum_out[16][23][23] = xor_out[80][23][23] + xor_out[81][23][23] + xor_out[82][23][23] + xor_out[83][23][23] + xor_out[84][23][23];
assign sum_out[17][23][23] = xor_out[85][23][23] + xor_out[86][23][23] + xor_out[87][23][23] + xor_out[88][23][23] + xor_out[89][23][23];
assign sum_out[18][23][23] = xor_out[90][23][23] + xor_out[91][23][23] + xor_out[92][23][23] + xor_out[93][23][23] + xor_out[94][23][23];
assign sum_out[19][23][23] = xor_out[95][23][23] + xor_out[96][23][23] + xor_out[97][23][23] + xor_out[98][23][23] + xor_out[99][23][23];


assign conv_one_out[0][0][0] = (sum_out[0][0][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][0][0] = (sum_out[1][0][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][0][0] = (sum_out[2][0][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][0][0] = (sum_out[3][0][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][0][0] = (sum_out[4][0][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][0][0] = (sum_out[5][0][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][0][0] = (sum_out[6][0][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][0][0] = (sum_out[7][0][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][0][0] = (sum_out[8][0][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][0][0] = (sum_out[9][0][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][0][0] = (sum_out[10][0][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][0][0] = (sum_out[11][0][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][0][0] = (sum_out[12][0][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][0][0] = (sum_out[13][0][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][0][0] = (sum_out[14][0][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][0][0] = (sum_out[15][0][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][0][0] = (sum_out[16][0][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][0][0] = (sum_out[17][0][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][0][0] = (sum_out[18][0][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][0][0] = (sum_out[19][0][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][0][1] = (sum_out[0][0][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][0][1] = (sum_out[1][0][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][0][1] = (sum_out[2][0][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][0][1] = (sum_out[3][0][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][0][1] = (sum_out[4][0][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][0][1] = (sum_out[5][0][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][0][1] = (sum_out[6][0][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][0][1] = (sum_out[7][0][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][0][1] = (sum_out[8][0][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][0][1] = (sum_out[9][0][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][0][1] = (sum_out[10][0][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][0][1] = (sum_out[11][0][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][0][1] = (sum_out[12][0][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][0][1] = (sum_out[13][0][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][0][1] = (sum_out[14][0][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][0][1] = (sum_out[15][0][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][0][1] = (sum_out[16][0][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][0][1] = (sum_out[17][0][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][0][1] = (sum_out[18][0][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][0][1] = (sum_out[19][0][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][0][2] = (sum_out[0][0][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][0][2] = (sum_out[1][0][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][0][2] = (sum_out[2][0][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][0][2] = (sum_out[3][0][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][0][2] = (sum_out[4][0][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][0][2] = (sum_out[5][0][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][0][2] = (sum_out[6][0][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][0][2] = (sum_out[7][0][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][0][2] = (sum_out[8][0][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][0][2] = (sum_out[9][0][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][0][2] = (sum_out[10][0][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][0][2] = (sum_out[11][0][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][0][2] = (sum_out[12][0][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][0][2] = (sum_out[13][0][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][0][2] = (sum_out[14][0][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][0][2] = (sum_out[15][0][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][0][2] = (sum_out[16][0][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][0][2] = (sum_out[17][0][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][0][2] = (sum_out[18][0][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][0][2] = (sum_out[19][0][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][0][3] = (sum_out[0][0][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][0][3] = (sum_out[1][0][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][0][3] = (sum_out[2][0][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][0][3] = (sum_out[3][0][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][0][3] = (sum_out[4][0][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][0][3] = (sum_out[5][0][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][0][3] = (sum_out[6][0][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][0][3] = (sum_out[7][0][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][0][3] = (sum_out[8][0][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][0][3] = (sum_out[9][0][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][0][3] = (sum_out[10][0][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][0][3] = (sum_out[11][0][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][0][3] = (sum_out[12][0][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][0][3] = (sum_out[13][0][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][0][3] = (sum_out[14][0][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][0][3] = (sum_out[15][0][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][0][3] = (sum_out[16][0][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][0][3] = (sum_out[17][0][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][0][3] = (sum_out[18][0][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][0][3] = (sum_out[19][0][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][0][4] = (sum_out[0][0][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][0][4] = (sum_out[1][0][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][0][4] = (sum_out[2][0][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][0][4] = (sum_out[3][0][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][0][4] = (sum_out[4][0][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][0][4] = (sum_out[5][0][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][0][4] = (sum_out[6][0][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][0][4] = (sum_out[7][0][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][0][4] = (sum_out[8][0][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][0][4] = (sum_out[9][0][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][0][4] = (sum_out[10][0][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][0][4] = (sum_out[11][0][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][0][4] = (sum_out[12][0][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][0][4] = (sum_out[13][0][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][0][4] = (sum_out[14][0][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][0][4] = (sum_out[15][0][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][0][4] = (sum_out[16][0][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][0][4] = (sum_out[17][0][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][0][4] = (sum_out[18][0][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][0][4] = (sum_out[19][0][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][0][5] = (sum_out[0][0][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][0][5] = (sum_out[1][0][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][0][5] = (sum_out[2][0][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][0][5] = (sum_out[3][0][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][0][5] = (sum_out[4][0][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][0][5] = (sum_out[5][0][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][0][5] = (sum_out[6][0][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][0][5] = (sum_out[7][0][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][0][5] = (sum_out[8][0][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][0][5] = (sum_out[9][0][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][0][5] = (sum_out[10][0][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][0][5] = (sum_out[11][0][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][0][5] = (sum_out[12][0][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][0][5] = (sum_out[13][0][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][0][5] = (sum_out[14][0][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][0][5] = (sum_out[15][0][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][0][5] = (sum_out[16][0][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][0][5] = (sum_out[17][0][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][0][5] = (sum_out[18][0][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][0][5] = (sum_out[19][0][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][0][6] = (sum_out[0][0][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][0][6] = (sum_out[1][0][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][0][6] = (sum_out[2][0][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][0][6] = (sum_out[3][0][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][0][6] = (sum_out[4][0][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][0][6] = (sum_out[5][0][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][0][6] = (sum_out[6][0][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][0][6] = (sum_out[7][0][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][0][6] = (sum_out[8][0][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][0][6] = (sum_out[9][0][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][0][6] = (sum_out[10][0][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][0][6] = (sum_out[11][0][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][0][6] = (sum_out[12][0][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][0][6] = (sum_out[13][0][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][0][6] = (sum_out[14][0][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][0][6] = (sum_out[15][0][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][0][6] = (sum_out[16][0][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][0][6] = (sum_out[17][0][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][0][6] = (sum_out[18][0][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][0][6] = (sum_out[19][0][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][0][7] = (sum_out[0][0][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][0][7] = (sum_out[1][0][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][0][7] = (sum_out[2][0][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][0][7] = (sum_out[3][0][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][0][7] = (sum_out[4][0][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][0][7] = (sum_out[5][0][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][0][7] = (sum_out[6][0][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][0][7] = (sum_out[7][0][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][0][7] = (sum_out[8][0][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][0][7] = (sum_out[9][0][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][0][7] = (sum_out[10][0][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][0][7] = (sum_out[11][0][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][0][7] = (sum_out[12][0][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][0][7] = (sum_out[13][0][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][0][7] = (sum_out[14][0][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][0][7] = (sum_out[15][0][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][0][7] = (sum_out[16][0][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][0][7] = (sum_out[17][0][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][0][7] = (sum_out[18][0][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][0][7] = (sum_out[19][0][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][0][8] = (sum_out[0][0][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][0][8] = (sum_out[1][0][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][0][8] = (sum_out[2][0][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][0][8] = (sum_out[3][0][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][0][8] = (sum_out[4][0][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][0][8] = (sum_out[5][0][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][0][8] = (sum_out[6][0][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][0][8] = (sum_out[7][0][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][0][8] = (sum_out[8][0][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][0][8] = (sum_out[9][0][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][0][8] = (sum_out[10][0][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][0][8] = (sum_out[11][0][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][0][8] = (sum_out[12][0][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][0][8] = (sum_out[13][0][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][0][8] = (sum_out[14][0][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][0][8] = (sum_out[15][0][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][0][8] = (sum_out[16][0][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][0][8] = (sum_out[17][0][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][0][8] = (sum_out[18][0][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][0][8] = (sum_out[19][0][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][0][9] = (sum_out[0][0][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][0][9] = (sum_out[1][0][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][0][9] = (sum_out[2][0][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][0][9] = (sum_out[3][0][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][0][9] = (sum_out[4][0][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][0][9] = (sum_out[5][0][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][0][9] = (sum_out[6][0][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][0][9] = (sum_out[7][0][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][0][9] = (sum_out[8][0][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][0][9] = (sum_out[9][0][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][0][9] = (sum_out[10][0][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][0][9] = (sum_out[11][0][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][0][9] = (sum_out[12][0][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][0][9] = (sum_out[13][0][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][0][9] = (sum_out[14][0][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][0][9] = (sum_out[15][0][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][0][9] = (sum_out[16][0][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][0][9] = (sum_out[17][0][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][0][9] = (sum_out[18][0][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][0][9] = (sum_out[19][0][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][0][10] = (sum_out[0][0][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][0][10] = (sum_out[1][0][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][0][10] = (sum_out[2][0][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][0][10] = (sum_out[3][0][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][0][10] = (sum_out[4][0][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][0][10] = (sum_out[5][0][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][0][10] = (sum_out[6][0][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][0][10] = (sum_out[7][0][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][0][10] = (sum_out[8][0][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][0][10] = (sum_out[9][0][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][0][10] = (sum_out[10][0][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][0][10] = (sum_out[11][0][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][0][10] = (sum_out[12][0][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][0][10] = (sum_out[13][0][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][0][10] = (sum_out[14][0][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][0][10] = (sum_out[15][0][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][0][10] = (sum_out[16][0][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][0][10] = (sum_out[17][0][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][0][10] = (sum_out[18][0][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][0][10] = (sum_out[19][0][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][0][11] = (sum_out[0][0][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][0][11] = (sum_out[1][0][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][0][11] = (sum_out[2][0][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][0][11] = (sum_out[3][0][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][0][11] = (sum_out[4][0][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][0][11] = (sum_out[5][0][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][0][11] = (sum_out[6][0][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][0][11] = (sum_out[7][0][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][0][11] = (sum_out[8][0][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][0][11] = (sum_out[9][0][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][0][11] = (sum_out[10][0][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][0][11] = (sum_out[11][0][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][0][11] = (sum_out[12][0][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][0][11] = (sum_out[13][0][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][0][11] = (sum_out[14][0][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][0][11] = (sum_out[15][0][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][0][11] = (sum_out[16][0][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][0][11] = (sum_out[17][0][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][0][11] = (sum_out[18][0][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][0][11] = (sum_out[19][0][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][0][12] = (sum_out[0][0][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][0][12] = (sum_out[1][0][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][0][12] = (sum_out[2][0][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][0][12] = (sum_out[3][0][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][0][12] = (sum_out[4][0][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][0][12] = (sum_out[5][0][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][0][12] = (sum_out[6][0][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][0][12] = (sum_out[7][0][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][0][12] = (sum_out[8][0][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][0][12] = (sum_out[9][0][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][0][12] = (sum_out[10][0][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][0][12] = (sum_out[11][0][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][0][12] = (sum_out[12][0][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][0][12] = (sum_out[13][0][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][0][12] = (sum_out[14][0][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][0][12] = (sum_out[15][0][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][0][12] = (sum_out[16][0][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][0][12] = (sum_out[17][0][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][0][12] = (sum_out[18][0][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][0][12] = (sum_out[19][0][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][0][13] = (sum_out[0][0][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][0][13] = (sum_out[1][0][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][0][13] = (sum_out[2][0][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][0][13] = (sum_out[3][0][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][0][13] = (sum_out[4][0][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][0][13] = (sum_out[5][0][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][0][13] = (sum_out[6][0][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][0][13] = (sum_out[7][0][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][0][13] = (sum_out[8][0][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][0][13] = (sum_out[9][0][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][0][13] = (sum_out[10][0][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][0][13] = (sum_out[11][0][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][0][13] = (sum_out[12][0][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][0][13] = (sum_out[13][0][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][0][13] = (sum_out[14][0][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][0][13] = (sum_out[15][0][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][0][13] = (sum_out[16][0][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][0][13] = (sum_out[17][0][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][0][13] = (sum_out[18][0][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][0][13] = (sum_out[19][0][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][0][14] = (sum_out[0][0][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][0][14] = (sum_out[1][0][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][0][14] = (sum_out[2][0][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][0][14] = (sum_out[3][0][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][0][14] = (sum_out[4][0][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][0][14] = (sum_out[5][0][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][0][14] = (sum_out[6][0][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][0][14] = (sum_out[7][0][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][0][14] = (sum_out[8][0][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][0][14] = (sum_out[9][0][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][0][14] = (sum_out[10][0][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][0][14] = (sum_out[11][0][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][0][14] = (sum_out[12][0][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][0][14] = (sum_out[13][0][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][0][14] = (sum_out[14][0][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][0][14] = (sum_out[15][0][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][0][14] = (sum_out[16][0][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][0][14] = (sum_out[17][0][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][0][14] = (sum_out[18][0][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][0][14] = (sum_out[19][0][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][0][15] = (sum_out[0][0][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][0][15] = (sum_out[1][0][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][0][15] = (sum_out[2][0][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][0][15] = (sum_out[3][0][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][0][15] = (sum_out[4][0][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][0][15] = (sum_out[5][0][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][0][15] = (sum_out[6][0][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][0][15] = (sum_out[7][0][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][0][15] = (sum_out[8][0][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][0][15] = (sum_out[9][0][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][0][15] = (sum_out[10][0][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][0][15] = (sum_out[11][0][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][0][15] = (sum_out[12][0][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][0][15] = (sum_out[13][0][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][0][15] = (sum_out[14][0][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][0][15] = (sum_out[15][0][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][0][15] = (sum_out[16][0][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][0][15] = (sum_out[17][0][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][0][15] = (sum_out[18][0][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][0][15] = (sum_out[19][0][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][0][16] = (sum_out[0][0][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][0][16] = (sum_out[1][0][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][0][16] = (sum_out[2][0][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][0][16] = (sum_out[3][0][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][0][16] = (sum_out[4][0][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][0][16] = (sum_out[5][0][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][0][16] = (sum_out[6][0][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][0][16] = (sum_out[7][0][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][0][16] = (sum_out[8][0][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][0][16] = (sum_out[9][0][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][0][16] = (sum_out[10][0][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][0][16] = (sum_out[11][0][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][0][16] = (sum_out[12][0][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][0][16] = (sum_out[13][0][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][0][16] = (sum_out[14][0][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][0][16] = (sum_out[15][0][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][0][16] = (sum_out[16][0][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][0][16] = (sum_out[17][0][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][0][16] = (sum_out[18][0][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][0][16] = (sum_out[19][0][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][0][17] = (sum_out[0][0][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][0][17] = (sum_out[1][0][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][0][17] = (sum_out[2][0][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][0][17] = (sum_out[3][0][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][0][17] = (sum_out[4][0][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][0][17] = (sum_out[5][0][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][0][17] = (sum_out[6][0][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][0][17] = (sum_out[7][0][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][0][17] = (sum_out[8][0][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][0][17] = (sum_out[9][0][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][0][17] = (sum_out[10][0][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][0][17] = (sum_out[11][0][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][0][17] = (sum_out[12][0][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][0][17] = (sum_out[13][0][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][0][17] = (sum_out[14][0][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][0][17] = (sum_out[15][0][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][0][17] = (sum_out[16][0][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][0][17] = (sum_out[17][0][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][0][17] = (sum_out[18][0][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][0][17] = (sum_out[19][0][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][0][18] = (sum_out[0][0][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][0][18] = (sum_out[1][0][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][0][18] = (sum_out[2][0][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][0][18] = (sum_out[3][0][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][0][18] = (sum_out[4][0][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][0][18] = (sum_out[5][0][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][0][18] = (sum_out[6][0][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][0][18] = (sum_out[7][0][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][0][18] = (sum_out[8][0][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][0][18] = (sum_out[9][0][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][0][18] = (sum_out[10][0][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][0][18] = (sum_out[11][0][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][0][18] = (sum_out[12][0][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][0][18] = (sum_out[13][0][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][0][18] = (sum_out[14][0][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][0][18] = (sum_out[15][0][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][0][18] = (sum_out[16][0][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][0][18] = (sum_out[17][0][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][0][18] = (sum_out[18][0][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][0][18] = (sum_out[19][0][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][0][19] = (sum_out[0][0][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][0][19] = (sum_out[1][0][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][0][19] = (sum_out[2][0][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][0][19] = (sum_out[3][0][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][0][19] = (sum_out[4][0][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][0][19] = (sum_out[5][0][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][0][19] = (sum_out[6][0][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][0][19] = (sum_out[7][0][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][0][19] = (sum_out[8][0][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][0][19] = (sum_out[9][0][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][0][19] = (sum_out[10][0][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][0][19] = (sum_out[11][0][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][0][19] = (sum_out[12][0][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][0][19] = (sum_out[13][0][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][0][19] = (sum_out[14][0][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][0][19] = (sum_out[15][0][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][0][19] = (sum_out[16][0][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][0][19] = (sum_out[17][0][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][0][19] = (sum_out[18][0][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][0][19] = (sum_out[19][0][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][0][20] = (sum_out[0][0][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][0][20] = (sum_out[1][0][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][0][20] = (sum_out[2][0][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][0][20] = (sum_out[3][0][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][0][20] = (sum_out[4][0][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][0][20] = (sum_out[5][0][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][0][20] = (sum_out[6][0][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][0][20] = (sum_out[7][0][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][0][20] = (sum_out[8][0][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][0][20] = (sum_out[9][0][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][0][20] = (sum_out[10][0][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][0][20] = (sum_out[11][0][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][0][20] = (sum_out[12][0][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][0][20] = (sum_out[13][0][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][0][20] = (sum_out[14][0][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][0][20] = (sum_out[15][0][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][0][20] = (sum_out[16][0][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][0][20] = (sum_out[17][0][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][0][20] = (sum_out[18][0][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][0][20] = (sum_out[19][0][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][0][21] = (sum_out[0][0][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][0][21] = (sum_out[1][0][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][0][21] = (sum_out[2][0][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][0][21] = (sum_out[3][0][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][0][21] = (sum_out[4][0][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][0][21] = (sum_out[5][0][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][0][21] = (sum_out[6][0][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][0][21] = (sum_out[7][0][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][0][21] = (sum_out[8][0][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][0][21] = (sum_out[9][0][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][0][21] = (sum_out[10][0][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][0][21] = (sum_out[11][0][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][0][21] = (sum_out[12][0][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][0][21] = (sum_out[13][0][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][0][21] = (sum_out[14][0][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][0][21] = (sum_out[15][0][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][0][21] = (sum_out[16][0][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][0][21] = (sum_out[17][0][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][0][21] = (sum_out[18][0][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][0][21] = (sum_out[19][0][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][0][22] = (sum_out[0][0][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][0][22] = (sum_out[1][0][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][0][22] = (sum_out[2][0][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][0][22] = (sum_out[3][0][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][0][22] = (sum_out[4][0][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][0][22] = (sum_out[5][0][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][0][22] = (sum_out[6][0][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][0][22] = (sum_out[7][0][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][0][22] = (sum_out[8][0][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][0][22] = (sum_out[9][0][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][0][22] = (sum_out[10][0][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][0][22] = (sum_out[11][0][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][0][22] = (sum_out[12][0][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][0][22] = (sum_out[13][0][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][0][22] = (sum_out[14][0][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][0][22] = (sum_out[15][0][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][0][22] = (sum_out[16][0][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][0][22] = (sum_out[17][0][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][0][22] = (sum_out[18][0][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][0][22] = (sum_out[19][0][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][0][23] = (sum_out[0][0][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][0][23] = (sum_out[1][0][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][0][23] = (sum_out[2][0][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][0][23] = (sum_out[3][0][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][0][23] = (sum_out[4][0][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][0][23] = (sum_out[5][0][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][0][23] = (sum_out[6][0][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][0][23] = (sum_out[7][0][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][0][23] = (sum_out[8][0][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][0][23] = (sum_out[9][0][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][0][23] = (sum_out[10][0][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][0][23] = (sum_out[11][0][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][0][23] = (sum_out[12][0][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][0][23] = (sum_out[13][0][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][0][23] = (sum_out[14][0][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][0][23] = (sum_out[15][0][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][0][23] = (sum_out[16][0][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][0][23] = (sum_out[17][0][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][0][23] = (sum_out[18][0][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][0][23] = (sum_out[19][0][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][1][0] = (sum_out[0][1][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][1][0] = (sum_out[1][1][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][1][0] = (sum_out[2][1][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][1][0] = (sum_out[3][1][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][1][0] = (sum_out[4][1][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][1][0] = (sum_out[5][1][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][1][0] = (sum_out[6][1][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][1][0] = (sum_out[7][1][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][1][0] = (sum_out[8][1][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][1][0] = (sum_out[9][1][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][1][0] = (sum_out[10][1][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][1][0] = (sum_out[11][1][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][1][0] = (sum_out[12][1][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][1][0] = (sum_out[13][1][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][1][0] = (sum_out[14][1][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][1][0] = (sum_out[15][1][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][1][0] = (sum_out[16][1][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][1][0] = (sum_out[17][1][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][1][0] = (sum_out[18][1][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][1][0] = (sum_out[19][1][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][1][1] = (sum_out[0][1][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][1][1] = (sum_out[1][1][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][1][1] = (sum_out[2][1][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][1][1] = (sum_out[3][1][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][1][1] = (sum_out[4][1][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][1][1] = (sum_out[5][1][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][1][1] = (sum_out[6][1][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][1][1] = (sum_out[7][1][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][1][1] = (sum_out[8][1][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][1][1] = (sum_out[9][1][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][1][1] = (sum_out[10][1][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][1][1] = (sum_out[11][1][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][1][1] = (sum_out[12][1][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][1][1] = (sum_out[13][1][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][1][1] = (sum_out[14][1][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][1][1] = (sum_out[15][1][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][1][1] = (sum_out[16][1][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][1][1] = (sum_out[17][1][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][1][1] = (sum_out[18][1][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][1][1] = (sum_out[19][1][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][1][2] = (sum_out[0][1][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][1][2] = (sum_out[1][1][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][1][2] = (sum_out[2][1][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][1][2] = (sum_out[3][1][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][1][2] = (sum_out[4][1][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][1][2] = (sum_out[5][1][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][1][2] = (sum_out[6][1][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][1][2] = (sum_out[7][1][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][1][2] = (sum_out[8][1][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][1][2] = (sum_out[9][1][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][1][2] = (sum_out[10][1][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][1][2] = (sum_out[11][1][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][1][2] = (sum_out[12][1][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][1][2] = (sum_out[13][1][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][1][2] = (sum_out[14][1][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][1][2] = (sum_out[15][1][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][1][2] = (sum_out[16][1][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][1][2] = (sum_out[17][1][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][1][2] = (sum_out[18][1][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][1][2] = (sum_out[19][1][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][1][3] = (sum_out[0][1][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][1][3] = (sum_out[1][1][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][1][3] = (sum_out[2][1][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][1][3] = (sum_out[3][1][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][1][3] = (sum_out[4][1][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][1][3] = (sum_out[5][1][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][1][3] = (sum_out[6][1][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][1][3] = (sum_out[7][1][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][1][3] = (sum_out[8][1][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][1][3] = (sum_out[9][1][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][1][3] = (sum_out[10][1][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][1][3] = (sum_out[11][1][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][1][3] = (sum_out[12][1][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][1][3] = (sum_out[13][1][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][1][3] = (sum_out[14][1][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][1][3] = (sum_out[15][1][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][1][3] = (sum_out[16][1][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][1][3] = (sum_out[17][1][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][1][3] = (sum_out[18][1][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][1][3] = (sum_out[19][1][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][1][4] = (sum_out[0][1][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][1][4] = (sum_out[1][1][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][1][4] = (sum_out[2][1][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][1][4] = (sum_out[3][1][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][1][4] = (sum_out[4][1][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][1][4] = (sum_out[5][1][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][1][4] = (sum_out[6][1][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][1][4] = (sum_out[7][1][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][1][4] = (sum_out[8][1][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][1][4] = (sum_out[9][1][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][1][4] = (sum_out[10][1][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][1][4] = (sum_out[11][1][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][1][4] = (sum_out[12][1][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][1][4] = (sum_out[13][1][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][1][4] = (sum_out[14][1][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][1][4] = (sum_out[15][1][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][1][4] = (sum_out[16][1][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][1][4] = (sum_out[17][1][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][1][4] = (sum_out[18][1][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][1][4] = (sum_out[19][1][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][1][5] = (sum_out[0][1][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][1][5] = (sum_out[1][1][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][1][5] = (sum_out[2][1][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][1][5] = (sum_out[3][1][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][1][5] = (sum_out[4][1][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][1][5] = (sum_out[5][1][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][1][5] = (sum_out[6][1][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][1][5] = (sum_out[7][1][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][1][5] = (sum_out[8][1][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][1][5] = (sum_out[9][1][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][1][5] = (sum_out[10][1][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][1][5] = (sum_out[11][1][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][1][5] = (sum_out[12][1][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][1][5] = (sum_out[13][1][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][1][5] = (sum_out[14][1][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][1][5] = (sum_out[15][1][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][1][5] = (sum_out[16][1][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][1][5] = (sum_out[17][1][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][1][5] = (sum_out[18][1][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][1][5] = (sum_out[19][1][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][1][6] = (sum_out[0][1][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][1][6] = (sum_out[1][1][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][1][6] = (sum_out[2][1][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][1][6] = (sum_out[3][1][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][1][6] = (sum_out[4][1][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][1][6] = (sum_out[5][1][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][1][6] = (sum_out[6][1][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][1][6] = (sum_out[7][1][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][1][6] = (sum_out[8][1][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][1][6] = (sum_out[9][1][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][1][6] = (sum_out[10][1][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][1][6] = (sum_out[11][1][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][1][6] = (sum_out[12][1][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][1][6] = (sum_out[13][1][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][1][6] = (sum_out[14][1][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][1][6] = (sum_out[15][1][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][1][6] = (sum_out[16][1][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][1][6] = (sum_out[17][1][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][1][6] = (sum_out[18][1][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][1][6] = (sum_out[19][1][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][1][7] = (sum_out[0][1][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][1][7] = (sum_out[1][1][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][1][7] = (sum_out[2][1][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][1][7] = (sum_out[3][1][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][1][7] = (sum_out[4][1][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][1][7] = (sum_out[5][1][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][1][7] = (sum_out[6][1][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][1][7] = (sum_out[7][1][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][1][7] = (sum_out[8][1][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][1][7] = (sum_out[9][1][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][1][7] = (sum_out[10][1][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][1][7] = (sum_out[11][1][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][1][7] = (sum_out[12][1][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][1][7] = (sum_out[13][1][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][1][7] = (sum_out[14][1][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][1][7] = (sum_out[15][1][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][1][7] = (sum_out[16][1][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][1][7] = (sum_out[17][1][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][1][7] = (sum_out[18][1][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][1][7] = (sum_out[19][1][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][1][8] = (sum_out[0][1][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][1][8] = (sum_out[1][1][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][1][8] = (sum_out[2][1][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][1][8] = (sum_out[3][1][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][1][8] = (sum_out[4][1][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][1][8] = (sum_out[5][1][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][1][8] = (sum_out[6][1][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][1][8] = (sum_out[7][1][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][1][8] = (sum_out[8][1][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][1][8] = (sum_out[9][1][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][1][8] = (sum_out[10][1][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][1][8] = (sum_out[11][1][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][1][8] = (sum_out[12][1][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][1][8] = (sum_out[13][1][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][1][8] = (sum_out[14][1][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][1][8] = (sum_out[15][1][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][1][8] = (sum_out[16][1][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][1][8] = (sum_out[17][1][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][1][8] = (sum_out[18][1][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][1][8] = (sum_out[19][1][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][1][9] = (sum_out[0][1][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][1][9] = (sum_out[1][1][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][1][9] = (sum_out[2][1][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][1][9] = (sum_out[3][1][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][1][9] = (sum_out[4][1][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][1][9] = (sum_out[5][1][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][1][9] = (sum_out[6][1][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][1][9] = (sum_out[7][1][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][1][9] = (sum_out[8][1][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][1][9] = (sum_out[9][1][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][1][9] = (sum_out[10][1][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][1][9] = (sum_out[11][1][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][1][9] = (sum_out[12][1][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][1][9] = (sum_out[13][1][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][1][9] = (sum_out[14][1][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][1][9] = (sum_out[15][1][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][1][9] = (sum_out[16][1][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][1][9] = (sum_out[17][1][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][1][9] = (sum_out[18][1][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][1][9] = (sum_out[19][1][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][1][10] = (sum_out[0][1][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][1][10] = (sum_out[1][1][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][1][10] = (sum_out[2][1][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][1][10] = (sum_out[3][1][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][1][10] = (sum_out[4][1][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][1][10] = (sum_out[5][1][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][1][10] = (sum_out[6][1][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][1][10] = (sum_out[7][1][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][1][10] = (sum_out[8][1][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][1][10] = (sum_out[9][1][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][1][10] = (sum_out[10][1][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][1][10] = (sum_out[11][1][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][1][10] = (sum_out[12][1][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][1][10] = (sum_out[13][1][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][1][10] = (sum_out[14][1][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][1][10] = (sum_out[15][1][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][1][10] = (sum_out[16][1][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][1][10] = (sum_out[17][1][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][1][10] = (sum_out[18][1][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][1][10] = (sum_out[19][1][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][1][11] = (sum_out[0][1][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][1][11] = (sum_out[1][1][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][1][11] = (sum_out[2][1][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][1][11] = (sum_out[3][1][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][1][11] = (sum_out[4][1][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][1][11] = (sum_out[5][1][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][1][11] = (sum_out[6][1][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][1][11] = (sum_out[7][1][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][1][11] = (sum_out[8][1][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][1][11] = (sum_out[9][1][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][1][11] = (sum_out[10][1][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][1][11] = (sum_out[11][1][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][1][11] = (sum_out[12][1][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][1][11] = (sum_out[13][1][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][1][11] = (sum_out[14][1][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][1][11] = (sum_out[15][1][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][1][11] = (sum_out[16][1][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][1][11] = (sum_out[17][1][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][1][11] = (sum_out[18][1][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][1][11] = (sum_out[19][1][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][1][12] = (sum_out[0][1][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][1][12] = (sum_out[1][1][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][1][12] = (sum_out[2][1][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][1][12] = (sum_out[3][1][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][1][12] = (sum_out[4][1][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][1][12] = (sum_out[5][1][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][1][12] = (sum_out[6][1][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][1][12] = (sum_out[7][1][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][1][12] = (sum_out[8][1][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][1][12] = (sum_out[9][1][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][1][12] = (sum_out[10][1][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][1][12] = (sum_out[11][1][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][1][12] = (sum_out[12][1][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][1][12] = (sum_out[13][1][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][1][12] = (sum_out[14][1][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][1][12] = (sum_out[15][1][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][1][12] = (sum_out[16][1][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][1][12] = (sum_out[17][1][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][1][12] = (sum_out[18][1][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][1][12] = (sum_out[19][1][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][1][13] = (sum_out[0][1][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][1][13] = (sum_out[1][1][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][1][13] = (sum_out[2][1][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][1][13] = (sum_out[3][1][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][1][13] = (sum_out[4][1][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][1][13] = (sum_out[5][1][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][1][13] = (sum_out[6][1][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][1][13] = (sum_out[7][1][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][1][13] = (sum_out[8][1][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][1][13] = (sum_out[9][1][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][1][13] = (sum_out[10][1][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][1][13] = (sum_out[11][1][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][1][13] = (sum_out[12][1][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][1][13] = (sum_out[13][1][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][1][13] = (sum_out[14][1][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][1][13] = (sum_out[15][1][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][1][13] = (sum_out[16][1][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][1][13] = (sum_out[17][1][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][1][13] = (sum_out[18][1][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][1][13] = (sum_out[19][1][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][1][14] = (sum_out[0][1][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][1][14] = (sum_out[1][1][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][1][14] = (sum_out[2][1][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][1][14] = (sum_out[3][1][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][1][14] = (sum_out[4][1][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][1][14] = (sum_out[5][1][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][1][14] = (sum_out[6][1][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][1][14] = (sum_out[7][1][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][1][14] = (sum_out[8][1][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][1][14] = (sum_out[9][1][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][1][14] = (sum_out[10][1][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][1][14] = (sum_out[11][1][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][1][14] = (sum_out[12][1][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][1][14] = (sum_out[13][1][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][1][14] = (sum_out[14][1][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][1][14] = (sum_out[15][1][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][1][14] = (sum_out[16][1][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][1][14] = (sum_out[17][1][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][1][14] = (sum_out[18][1][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][1][14] = (sum_out[19][1][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][1][15] = (sum_out[0][1][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][1][15] = (sum_out[1][1][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][1][15] = (sum_out[2][1][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][1][15] = (sum_out[3][1][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][1][15] = (sum_out[4][1][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][1][15] = (sum_out[5][1][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][1][15] = (sum_out[6][1][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][1][15] = (sum_out[7][1][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][1][15] = (sum_out[8][1][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][1][15] = (sum_out[9][1][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][1][15] = (sum_out[10][1][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][1][15] = (sum_out[11][1][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][1][15] = (sum_out[12][1][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][1][15] = (sum_out[13][1][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][1][15] = (sum_out[14][1][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][1][15] = (sum_out[15][1][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][1][15] = (sum_out[16][1][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][1][15] = (sum_out[17][1][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][1][15] = (sum_out[18][1][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][1][15] = (sum_out[19][1][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][1][16] = (sum_out[0][1][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][1][16] = (sum_out[1][1][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][1][16] = (sum_out[2][1][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][1][16] = (sum_out[3][1][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][1][16] = (sum_out[4][1][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][1][16] = (sum_out[5][1][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][1][16] = (sum_out[6][1][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][1][16] = (sum_out[7][1][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][1][16] = (sum_out[8][1][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][1][16] = (sum_out[9][1][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][1][16] = (sum_out[10][1][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][1][16] = (sum_out[11][1][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][1][16] = (sum_out[12][1][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][1][16] = (sum_out[13][1][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][1][16] = (sum_out[14][1][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][1][16] = (sum_out[15][1][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][1][16] = (sum_out[16][1][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][1][16] = (sum_out[17][1][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][1][16] = (sum_out[18][1][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][1][16] = (sum_out[19][1][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][1][17] = (sum_out[0][1][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][1][17] = (sum_out[1][1][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][1][17] = (sum_out[2][1][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][1][17] = (sum_out[3][1][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][1][17] = (sum_out[4][1][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][1][17] = (sum_out[5][1][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][1][17] = (sum_out[6][1][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][1][17] = (sum_out[7][1][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][1][17] = (sum_out[8][1][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][1][17] = (sum_out[9][1][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][1][17] = (sum_out[10][1][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][1][17] = (sum_out[11][1][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][1][17] = (sum_out[12][1][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][1][17] = (sum_out[13][1][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][1][17] = (sum_out[14][1][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][1][17] = (sum_out[15][1][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][1][17] = (sum_out[16][1][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][1][17] = (sum_out[17][1][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][1][17] = (sum_out[18][1][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][1][17] = (sum_out[19][1][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][1][18] = (sum_out[0][1][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][1][18] = (sum_out[1][1][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][1][18] = (sum_out[2][1][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][1][18] = (sum_out[3][1][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][1][18] = (sum_out[4][1][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][1][18] = (sum_out[5][1][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][1][18] = (sum_out[6][1][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][1][18] = (sum_out[7][1][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][1][18] = (sum_out[8][1][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][1][18] = (sum_out[9][1][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][1][18] = (sum_out[10][1][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][1][18] = (sum_out[11][1][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][1][18] = (sum_out[12][1][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][1][18] = (sum_out[13][1][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][1][18] = (sum_out[14][1][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][1][18] = (sum_out[15][1][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][1][18] = (sum_out[16][1][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][1][18] = (sum_out[17][1][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][1][18] = (sum_out[18][1][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][1][18] = (sum_out[19][1][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][1][19] = (sum_out[0][1][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][1][19] = (sum_out[1][1][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][1][19] = (sum_out[2][1][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][1][19] = (sum_out[3][1][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][1][19] = (sum_out[4][1][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][1][19] = (sum_out[5][1][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][1][19] = (sum_out[6][1][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][1][19] = (sum_out[7][1][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][1][19] = (sum_out[8][1][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][1][19] = (sum_out[9][1][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][1][19] = (sum_out[10][1][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][1][19] = (sum_out[11][1][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][1][19] = (sum_out[12][1][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][1][19] = (sum_out[13][1][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][1][19] = (sum_out[14][1][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][1][19] = (sum_out[15][1][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][1][19] = (sum_out[16][1][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][1][19] = (sum_out[17][1][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][1][19] = (sum_out[18][1][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][1][19] = (sum_out[19][1][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][1][20] = (sum_out[0][1][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][1][20] = (sum_out[1][1][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][1][20] = (sum_out[2][1][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][1][20] = (sum_out[3][1][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][1][20] = (sum_out[4][1][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][1][20] = (sum_out[5][1][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][1][20] = (sum_out[6][1][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][1][20] = (sum_out[7][1][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][1][20] = (sum_out[8][1][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][1][20] = (sum_out[9][1][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][1][20] = (sum_out[10][1][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][1][20] = (sum_out[11][1][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][1][20] = (sum_out[12][1][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][1][20] = (sum_out[13][1][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][1][20] = (sum_out[14][1][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][1][20] = (sum_out[15][1][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][1][20] = (sum_out[16][1][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][1][20] = (sum_out[17][1][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][1][20] = (sum_out[18][1][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][1][20] = (sum_out[19][1][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][1][21] = (sum_out[0][1][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][1][21] = (sum_out[1][1][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][1][21] = (sum_out[2][1][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][1][21] = (sum_out[3][1][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][1][21] = (sum_out[4][1][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][1][21] = (sum_out[5][1][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][1][21] = (sum_out[6][1][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][1][21] = (sum_out[7][1][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][1][21] = (sum_out[8][1][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][1][21] = (sum_out[9][1][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][1][21] = (sum_out[10][1][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][1][21] = (sum_out[11][1][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][1][21] = (sum_out[12][1][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][1][21] = (sum_out[13][1][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][1][21] = (sum_out[14][1][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][1][21] = (sum_out[15][1][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][1][21] = (sum_out[16][1][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][1][21] = (sum_out[17][1][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][1][21] = (sum_out[18][1][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][1][21] = (sum_out[19][1][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][1][22] = (sum_out[0][1][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][1][22] = (sum_out[1][1][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][1][22] = (sum_out[2][1][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][1][22] = (sum_out[3][1][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][1][22] = (sum_out[4][1][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][1][22] = (sum_out[5][1][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][1][22] = (sum_out[6][1][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][1][22] = (sum_out[7][1][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][1][22] = (sum_out[8][1][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][1][22] = (sum_out[9][1][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][1][22] = (sum_out[10][1][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][1][22] = (sum_out[11][1][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][1][22] = (sum_out[12][1][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][1][22] = (sum_out[13][1][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][1][22] = (sum_out[14][1][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][1][22] = (sum_out[15][1][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][1][22] = (sum_out[16][1][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][1][22] = (sum_out[17][1][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][1][22] = (sum_out[18][1][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][1][22] = (sum_out[19][1][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][1][23] = (sum_out[0][1][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][1][23] = (sum_out[1][1][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][1][23] = (sum_out[2][1][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][1][23] = (sum_out[3][1][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][1][23] = (sum_out[4][1][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][1][23] = (sum_out[5][1][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][1][23] = (sum_out[6][1][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][1][23] = (sum_out[7][1][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][1][23] = (sum_out[8][1][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][1][23] = (sum_out[9][1][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][1][23] = (sum_out[10][1][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][1][23] = (sum_out[11][1][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][1][23] = (sum_out[12][1][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][1][23] = (sum_out[13][1][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][1][23] = (sum_out[14][1][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][1][23] = (sum_out[15][1][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][1][23] = (sum_out[16][1][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][1][23] = (sum_out[17][1][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][1][23] = (sum_out[18][1][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][1][23] = (sum_out[19][1][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][2][0] = (sum_out[0][2][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][2][0] = (sum_out[1][2][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][2][0] = (sum_out[2][2][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][2][0] = (sum_out[3][2][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][2][0] = (sum_out[4][2][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][2][0] = (sum_out[5][2][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][2][0] = (sum_out[6][2][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][2][0] = (sum_out[7][2][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][2][0] = (sum_out[8][2][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][2][0] = (sum_out[9][2][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][2][0] = (sum_out[10][2][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][2][0] = (sum_out[11][2][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][2][0] = (sum_out[12][2][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][2][0] = (sum_out[13][2][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][2][0] = (sum_out[14][2][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][2][0] = (sum_out[15][2][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][2][0] = (sum_out[16][2][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][2][0] = (sum_out[17][2][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][2][0] = (sum_out[18][2][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][2][0] = (sum_out[19][2][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][2][1] = (sum_out[0][2][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][2][1] = (sum_out[1][2][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][2][1] = (sum_out[2][2][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][2][1] = (sum_out[3][2][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][2][1] = (sum_out[4][2][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][2][1] = (sum_out[5][2][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][2][1] = (sum_out[6][2][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][2][1] = (sum_out[7][2][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][2][1] = (sum_out[8][2][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][2][1] = (sum_out[9][2][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][2][1] = (sum_out[10][2][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][2][1] = (sum_out[11][2][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][2][1] = (sum_out[12][2][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][2][1] = (sum_out[13][2][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][2][1] = (sum_out[14][2][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][2][1] = (sum_out[15][2][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][2][1] = (sum_out[16][2][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][2][1] = (sum_out[17][2][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][2][1] = (sum_out[18][2][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][2][1] = (sum_out[19][2][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][2][2] = (sum_out[0][2][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][2][2] = (sum_out[1][2][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][2][2] = (sum_out[2][2][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][2][2] = (sum_out[3][2][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][2][2] = (sum_out[4][2][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][2][2] = (sum_out[5][2][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][2][2] = (sum_out[6][2][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][2][2] = (sum_out[7][2][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][2][2] = (sum_out[8][2][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][2][2] = (sum_out[9][2][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][2][2] = (sum_out[10][2][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][2][2] = (sum_out[11][2][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][2][2] = (sum_out[12][2][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][2][2] = (sum_out[13][2][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][2][2] = (sum_out[14][2][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][2][2] = (sum_out[15][2][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][2][2] = (sum_out[16][2][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][2][2] = (sum_out[17][2][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][2][2] = (sum_out[18][2][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][2][2] = (sum_out[19][2][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][2][3] = (sum_out[0][2][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][2][3] = (sum_out[1][2][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][2][3] = (sum_out[2][2][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][2][3] = (sum_out[3][2][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][2][3] = (sum_out[4][2][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][2][3] = (sum_out[5][2][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][2][3] = (sum_out[6][2][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][2][3] = (sum_out[7][2][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][2][3] = (sum_out[8][2][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][2][3] = (sum_out[9][2][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][2][3] = (sum_out[10][2][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][2][3] = (sum_out[11][2][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][2][3] = (sum_out[12][2][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][2][3] = (sum_out[13][2][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][2][3] = (sum_out[14][2][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][2][3] = (sum_out[15][2][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][2][3] = (sum_out[16][2][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][2][3] = (sum_out[17][2][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][2][3] = (sum_out[18][2][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][2][3] = (sum_out[19][2][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][2][4] = (sum_out[0][2][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][2][4] = (sum_out[1][2][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][2][4] = (sum_out[2][2][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][2][4] = (sum_out[3][2][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][2][4] = (sum_out[4][2][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][2][4] = (sum_out[5][2][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][2][4] = (sum_out[6][2][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][2][4] = (sum_out[7][2][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][2][4] = (sum_out[8][2][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][2][4] = (sum_out[9][2][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][2][4] = (sum_out[10][2][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][2][4] = (sum_out[11][2][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][2][4] = (sum_out[12][2][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][2][4] = (sum_out[13][2][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][2][4] = (sum_out[14][2][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][2][4] = (sum_out[15][2][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][2][4] = (sum_out[16][2][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][2][4] = (sum_out[17][2][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][2][4] = (sum_out[18][2][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][2][4] = (sum_out[19][2][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][2][5] = (sum_out[0][2][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][2][5] = (sum_out[1][2][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][2][5] = (sum_out[2][2][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][2][5] = (sum_out[3][2][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][2][5] = (sum_out[4][2][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][2][5] = (sum_out[5][2][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][2][5] = (sum_out[6][2][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][2][5] = (sum_out[7][2][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][2][5] = (sum_out[8][2][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][2][5] = (sum_out[9][2][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][2][5] = (sum_out[10][2][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][2][5] = (sum_out[11][2][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][2][5] = (sum_out[12][2][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][2][5] = (sum_out[13][2][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][2][5] = (sum_out[14][2][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][2][5] = (sum_out[15][2][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][2][5] = (sum_out[16][2][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][2][5] = (sum_out[17][2][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][2][5] = (sum_out[18][2][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][2][5] = (sum_out[19][2][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][2][6] = (sum_out[0][2][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][2][6] = (sum_out[1][2][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][2][6] = (sum_out[2][2][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][2][6] = (sum_out[3][2][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][2][6] = (sum_out[4][2][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][2][6] = (sum_out[5][2][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][2][6] = (sum_out[6][2][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][2][6] = (sum_out[7][2][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][2][6] = (sum_out[8][2][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][2][6] = (sum_out[9][2][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][2][6] = (sum_out[10][2][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][2][6] = (sum_out[11][2][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][2][6] = (sum_out[12][2][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][2][6] = (sum_out[13][2][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][2][6] = (sum_out[14][2][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][2][6] = (sum_out[15][2][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][2][6] = (sum_out[16][2][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][2][6] = (sum_out[17][2][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][2][6] = (sum_out[18][2][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][2][6] = (sum_out[19][2][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][2][7] = (sum_out[0][2][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][2][7] = (sum_out[1][2][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][2][7] = (sum_out[2][2][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][2][7] = (sum_out[3][2][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][2][7] = (sum_out[4][2][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][2][7] = (sum_out[5][2][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][2][7] = (sum_out[6][2][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][2][7] = (sum_out[7][2][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][2][7] = (sum_out[8][2][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][2][7] = (sum_out[9][2][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][2][7] = (sum_out[10][2][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][2][7] = (sum_out[11][2][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][2][7] = (sum_out[12][2][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][2][7] = (sum_out[13][2][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][2][7] = (sum_out[14][2][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][2][7] = (sum_out[15][2][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][2][7] = (sum_out[16][2][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][2][7] = (sum_out[17][2][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][2][7] = (sum_out[18][2][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][2][7] = (sum_out[19][2][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][2][8] = (sum_out[0][2][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][2][8] = (sum_out[1][2][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][2][8] = (sum_out[2][2][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][2][8] = (sum_out[3][2][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][2][8] = (sum_out[4][2][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][2][8] = (sum_out[5][2][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][2][8] = (sum_out[6][2][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][2][8] = (sum_out[7][2][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][2][8] = (sum_out[8][2][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][2][8] = (sum_out[9][2][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][2][8] = (sum_out[10][2][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][2][8] = (sum_out[11][2][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][2][8] = (sum_out[12][2][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][2][8] = (sum_out[13][2][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][2][8] = (sum_out[14][2][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][2][8] = (sum_out[15][2][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][2][8] = (sum_out[16][2][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][2][8] = (sum_out[17][2][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][2][8] = (sum_out[18][2][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][2][8] = (sum_out[19][2][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][2][9] = (sum_out[0][2][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][2][9] = (sum_out[1][2][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][2][9] = (sum_out[2][2][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][2][9] = (sum_out[3][2][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][2][9] = (sum_out[4][2][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][2][9] = (sum_out[5][2][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][2][9] = (sum_out[6][2][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][2][9] = (sum_out[7][2][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][2][9] = (sum_out[8][2][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][2][9] = (sum_out[9][2][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][2][9] = (sum_out[10][2][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][2][9] = (sum_out[11][2][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][2][9] = (sum_out[12][2][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][2][9] = (sum_out[13][2][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][2][9] = (sum_out[14][2][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][2][9] = (sum_out[15][2][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][2][9] = (sum_out[16][2][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][2][9] = (sum_out[17][2][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][2][9] = (sum_out[18][2][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][2][9] = (sum_out[19][2][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][2][10] = (sum_out[0][2][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][2][10] = (sum_out[1][2][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][2][10] = (sum_out[2][2][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][2][10] = (sum_out[3][2][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][2][10] = (sum_out[4][2][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][2][10] = (sum_out[5][2][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][2][10] = (sum_out[6][2][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][2][10] = (sum_out[7][2][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][2][10] = (sum_out[8][2][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][2][10] = (sum_out[9][2][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][2][10] = (sum_out[10][2][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][2][10] = (sum_out[11][2][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][2][10] = (sum_out[12][2][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][2][10] = (sum_out[13][2][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][2][10] = (sum_out[14][2][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][2][10] = (sum_out[15][2][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][2][10] = (sum_out[16][2][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][2][10] = (sum_out[17][2][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][2][10] = (sum_out[18][2][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][2][10] = (sum_out[19][2][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][2][11] = (sum_out[0][2][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][2][11] = (sum_out[1][2][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][2][11] = (sum_out[2][2][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][2][11] = (sum_out[3][2][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][2][11] = (sum_out[4][2][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][2][11] = (sum_out[5][2][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][2][11] = (sum_out[6][2][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][2][11] = (sum_out[7][2][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][2][11] = (sum_out[8][2][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][2][11] = (sum_out[9][2][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][2][11] = (sum_out[10][2][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][2][11] = (sum_out[11][2][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][2][11] = (sum_out[12][2][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][2][11] = (sum_out[13][2][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][2][11] = (sum_out[14][2][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][2][11] = (sum_out[15][2][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][2][11] = (sum_out[16][2][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][2][11] = (sum_out[17][2][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][2][11] = (sum_out[18][2][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][2][11] = (sum_out[19][2][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][2][12] = (sum_out[0][2][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][2][12] = (sum_out[1][2][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][2][12] = (sum_out[2][2][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][2][12] = (sum_out[3][2][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][2][12] = (sum_out[4][2][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][2][12] = (sum_out[5][2][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][2][12] = (sum_out[6][2][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][2][12] = (sum_out[7][2][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][2][12] = (sum_out[8][2][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][2][12] = (sum_out[9][2][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][2][12] = (sum_out[10][2][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][2][12] = (sum_out[11][2][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][2][12] = (sum_out[12][2][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][2][12] = (sum_out[13][2][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][2][12] = (sum_out[14][2][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][2][12] = (sum_out[15][2][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][2][12] = (sum_out[16][2][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][2][12] = (sum_out[17][2][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][2][12] = (sum_out[18][2][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][2][12] = (sum_out[19][2][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][2][13] = (sum_out[0][2][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][2][13] = (sum_out[1][2][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][2][13] = (sum_out[2][2][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][2][13] = (sum_out[3][2][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][2][13] = (sum_out[4][2][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][2][13] = (sum_out[5][2][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][2][13] = (sum_out[6][2][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][2][13] = (sum_out[7][2][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][2][13] = (sum_out[8][2][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][2][13] = (sum_out[9][2][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][2][13] = (sum_out[10][2][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][2][13] = (sum_out[11][2][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][2][13] = (sum_out[12][2][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][2][13] = (sum_out[13][2][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][2][13] = (sum_out[14][2][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][2][13] = (sum_out[15][2][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][2][13] = (sum_out[16][2][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][2][13] = (sum_out[17][2][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][2][13] = (sum_out[18][2][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][2][13] = (sum_out[19][2][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][2][14] = (sum_out[0][2][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][2][14] = (sum_out[1][2][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][2][14] = (sum_out[2][2][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][2][14] = (sum_out[3][2][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][2][14] = (sum_out[4][2][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][2][14] = (sum_out[5][2][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][2][14] = (sum_out[6][2][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][2][14] = (sum_out[7][2][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][2][14] = (sum_out[8][2][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][2][14] = (sum_out[9][2][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][2][14] = (sum_out[10][2][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][2][14] = (sum_out[11][2][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][2][14] = (sum_out[12][2][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][2][14] = (sum_out[13][2][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][2][14] = (sum_out[14][2][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][2][14] = (sum_out[15][2][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][2][14] = (sum_out[16][2][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][2][14] = (sum_out[17][2][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][2][14] = (sum_out[18][2][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][2][14] = (sum_out[19][2][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][2][15] = (sum_out[0][2][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][2][15] = (sum_out[1][2][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][2][15] = (sum_out[2][2][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][2][15] = (sum_out[3][2][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][2][15] = (sum_out[4][2][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][2][15] = (sum_out[5][2][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][2][15] = (sum_out[6][2][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][2][15] = (sum_out[7][2][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][2][15] = (sum_out[8][2][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][2][15] = (sum_out[9][2][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][2][15] = (sum_out[10][2][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][2][15] = (sum_out[11][2][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][2][15] = (sum_out[12][2][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][2][15] = (sum_out[13][2][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][2][15] = (sum_out[14][2][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][2][15] = (sum_out[15][2][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][2][15] = (sum_out[16][2][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][2][15] = (sum_out[17][2][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][2][15] = (sum_out[18][2][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][2][15] = (sum_out[19][2][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][2][16] = (sum_out[0][2][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][2][16] = (sum_out[1][2][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][2][16] = (sum_out[2][2][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][2][16] = (sum_out[3][2][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][2][16] = (sum_out[4][2][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][2][16] = (sum_out[5][2][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][2][16] = (sum_out[6][2][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][2][16] = (sum_out[7][2][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][2][16] = (sum_out[8][2][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][2][16] = (sum_out[9][2][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][2][16] = (sum_out[10][2][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][2][16] = (sum_out[11][2][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][2][16] = (sum_out[12][2][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][2][16] = (sum_out[13][2][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][2][16] = (sum_out[14][2][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][2][16] = (sum_out[15][2][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][2][16] = (sum_out[16][2][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][2][16] = (sum_out[17][2][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][2][16] = (sum_out[18][2][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][2][16] = (sum_out[19][2][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][2][17] = (sum_out[0][2][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][2][17] = (sum_out[1][2][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][2][17] = (sum_out[2][2][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][2][17] = (sum_out[3][2][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][2][17] = (sum_out[4][2][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][2][17] = (sum_out[5][2][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][2][17] = (sum_out[6][2][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][2][17] = (sum_out[7][2][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][2][17] = (sum_out[8][2][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][2][17] = (sum_out[9][2][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][2][17] = (sum_out[10][2][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][2][17] = (sum_out[11][2][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][2][17] = (sum_out[12][2][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][2][17] = (sum_out[13][2][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][2][17] = (sum_out[14][2][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][2][17] = (sum_out[15][2][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][2][17] = (sum_out[16][2][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][2][17] = (sum_out[17][2][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][2][17] = (sum_out[18][2][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][2][17] = (sum_out[19][2][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][2][18] = (sum_out[0][2][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][2][18] = (sum_out[1][2][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][2][18] = (sum_out[2][2][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][2][18] = (sum_out[3][2][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][2][18] = (sum_out[4][2][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][2][18] = (sum_out[5][2][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][2][18] = (sum_out[6][2][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][2][18] = (sum_out[7][2][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][2][18] = (sum_out[8][2][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][2][18] = (sum_out[9][2][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][2][18] = (sum_out[10][2][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][2][18] = (sum_out[11][2][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][2][18] = (sum_out[12][2][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][2][18] = (sum_out[13][2][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][2][18] = (sum_out[14][2][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][2][18] = (sum_out[15][2][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][2][18] = (sum_out[16][2][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][2][18] = (sum_out[17][2][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][2][18] = (sum_out[18][2][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][2][18] = (sum_out[19][2][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][2][19] = (sum_out[0][2][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][2][19] = (sum_out[1][2][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][2][19] = (sum_out[2][2][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][2][19] = (sum_out[3][2][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][2][19] = (sum_out[4][2][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][2][19] = (sum_out[5][2][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][2][19] = (sum_out[6][2][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][2][19] = (sum_out[7][2][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][2][19] = (sum_out[8][2][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][2][19] = (sum_out[9][2][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][2][19] = (sum_out[10][2][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][2][19] = (sum_out[11][2][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][2][19] = (sum_out[12][2][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][2][19] = (sum_out[13][2][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][2][19] = (sum_out[14][2][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][2][19] = (sum_out[15][2][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][2][19] = (sum_out[16][2][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][2][19] = (sum_out[17][2][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][2][19] = (sum_out[18][2][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][2][19] = (sum_out[19][2][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][2][20] = (sum_out[0][2][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][2][20] = (sum_out[1][2][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][2][20] = (sum_out[2][2][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][2][20] = (sum_out[3][2][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][2][20] = (sum_out[4][2][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][2][20] = (sum_out[5][2][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][2][20] = (sum_out[6][2][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][2][20] = (sum_out[7][2][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][2][20] = (sum_out[8][2][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][2][20] = (sum_out[9][2][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][2][20] = (sum_out[10][2][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][2][20] = (sum_out[11][2][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][2][20] = (sum_out[12][2][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][2][20] = (sum_out[13][2][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][2][20] = (sum_out[14][2][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][2][20] = (sum_out[15][2][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][2][20] = (sum_out[16][2][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][2][20] = (sum_out[17][2][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][2][20] = (sum_out[18][2][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][2][20] = (sum_out[19][2][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][2][21] = (sum_out[0][2][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][2][21] = (sum_out[1][2][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][2][21] = (sum_out[2][2][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][2][21] = (sum_out[3][2][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][2][21] = (sum_out[4][2][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][2][21] = (sum_out[5][2][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][2][21] = (sum_out[6][2][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][2][21] = (sum_out[7][2][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][2][21] = (sum_out[8][2][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][2][21] = (sum_out[9][2][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][2][21] = (sum_out[10][2][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][2][21] = (sum_out[11][2][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][2][21] = (sum_out[12][2][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][2][21] = (sum_out[13][2][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][2][21] = (sum_out[14][2][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][2][21] = (sum_out[15][2][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][2][21] = (sum_out[16][2][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][2][21] = (sum_out[17][2][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][2][21] = (sum_out[18][2][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][2][21] = (sum_out[19][2][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][2][22] = (sum_out[0][2][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][2][22] = (sum_out[1][2][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][2][22] = (sum_out[2][2][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][2][22] = (sum_out[3][2][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][2][22] = (sum_out[4][2][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][2][22] = (sum_out[5][2][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][2][22] = (sum_out[6][2][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][2][22] = (sum_out[7][2][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][2][22] = (sum_out[8][2][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][2][22] = (sum_out[9][2][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][2][22] = (sum_out[10][2][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][2][22] = (sum_out[11][2][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][2][22] = (sum_out[12][2][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][2][22] = (sum_out[13][2][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][2][22] = (sum_out[14][2][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][2][22] = (sum_out[15][2][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][2][22] = (sum_out[16][2][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][2][22] = (sum_out[17][2][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][2][22] = (sum_out[18][2][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][2][22] = (sum_out[19][2][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][2][23] = (sum_out[0][2][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][2][23] = (sum_out[1][2][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][2][23] = (sum_out[2][2][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][2][23] = (sum_out[3][2][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][2][23] = (sum_out[4][2][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][2][23] = (sum_out[5][2][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][2][23] = (sum_out[6][2][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][2][23] = (sum_out[7][2][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][2][23] = (sum_out[8][2][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][2][23] = (sum_out[9][2][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][2][23] = (sum_out[10][2][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][2][23] = (sum_out[11][2][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][2][23] = (sum_out[12][2][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][2][23] = (sum_out[13][2][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][2][23] = (sum_out[14][2][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][2][23] = (sum_out[15][2][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][2][23] = (sum_out[16][2][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][2][23] = (sum_out[17][2][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][2][23] = (sum_out[18][2][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][2][23] = (sum_out[19][2][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][3][0] = (sum_out[0][3][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][3][0] = (sum_out[1][3][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][3][0] = (sum_out[2][3][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][3][0] = (sum_out[3][3][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][3][0] = (sum_out[4][3][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][3][0] = (sum_out[5][3][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][3][0] = (sum_out[6][3][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][3][0] = (sum_out[7][3][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][3][0] = (sum_out[8][3][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][3][0] = (sum_out[9][3][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][3][0] = (sum_out[10][3][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][3][0] = (sum_out[11][3][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][3][0] = (sum_out[12][3][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][3][0] = (sum_out[13][3][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][3][0] = (sum_out[14][3][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][3][0] = (sum_out[15][3][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][3][0] = (sum_out[16][3][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][3][0] = (sum_out[17][3][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][3][0] = (sum_out[18][3][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][3][0] = (sum_out[19][3][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][3][1] = (sum_out[0][3][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][3][1] = (sum_out[1][3][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][3][1] = (sum_out[2][3][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][3][1] = (sum_out[3][3][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][3][1] = (sum_out[4][3][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][3][1] = (sum_out[5][3][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][3][1] = (sum_out[6][3][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][3][1] = (sum_out[7][3][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][3][1] = (sum_out[8][3][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][3][1] = (sum_out[9][3][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][3][1] = (sum_out[10][3][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][3][1] = (sum_out[11][3][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][3][1] = (sum_out[12][3][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][3][1] = (sum_out[13][3][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][3][1] = (sum_out[14][3][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][3][1] = (sum_out[15][3][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][3][1] = (sum_out[16][3][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][3][1] = (sum_out[17][3][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][3][1] = (sum_out[18][3][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][3][1] = (sum_out[19][3][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][3][2] = (sum_out[0][3][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][3][2] = (sum_out[1][3][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][3][2] = (sum_out[2][3][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][3][2] = (sum_out[3][3][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][3][2] = (sum_out[4][3][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][3][2] = (sum_out[5][3][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][3][2] = (sum_out[6][3][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][3][2] = (sum_out[7][3][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][3][2] = (sum_out[8][3][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][3][2] = (sum_out[9][3][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][3][2] = (sum_out[10][3][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][3][2] = (sum_out[11][3][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][3][2] = (sum_out[12][3][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][3][2] = (sum_out[13][3][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][3][2] = (sum_out[14][3][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][3][2] = (sum_out[15][3][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][3][2] = (sum_out[16][3][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][3][2] = (sum_out[17][3][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][3][2] = (sum_out[18][3][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][3][2] = (sum_out[19][3][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][3][3] = (sum_out[0][3][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][3][3] = (sum_out[1][3][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][3][3] = (sum_out[2][3][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][3][3] = (sum_out[3][3][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][3][3] = (sum_out[4][3][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][3][3] = (sum_out[5][3][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][3][3] = (sum_out[6][3][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][3][3] = (sum_out[7][3][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][3][3] = (sum_out[8][3][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][3][3] = (sum_out[9][3][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][3][3] = (sum_out[10][3][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][3][3] = (sum_out[11][3][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][3][3] = (sum_out[12][3][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][3][3] = (sum_out[13][3][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][3][3] = (sum_out[14][3][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][3][3] = (sum_out[15][3][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][3][3] = (sum_out[16][3][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][3][3] = (sum_out[17][3][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][3][3] = (sum_out[18][3][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][3][3] = (sum_out[19][3][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][3][4] = (sum_out[0][3][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][3][4] = (sum_out[1][3][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][3][4] = (sum_out[2][3][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][3][4] = (sum_out[3][3][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][3][4] = (sum_out[4][3][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][3][4] = (sum_out[5][3][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][3][4] = (sum_out[6][3][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][3][4] = (sum_out[7][3][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][3][4] = (sum_out[8][3][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][3][4] = (sum_out[9][3][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][3][4] = (sum_out[10][3][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][3][4] = (sum_out[11][3][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][3][4] = (sum_out[12][3][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][3][4] = (sum_out[13][3][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][3][4] = (sum_out[14][3][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][3][4] = (sum_out[15][3][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][3][4] = (sum_out[16][3][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][3][4] = (sum_out[17][3][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][3][4] = (sum_out[18][3][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][3][4] = (sum_out[19][3][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][3][5] = (sum_out[0][3][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][3][5] = (sum_out[1][3][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][3][5] = (sum_out[2][3][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][3][5] = (sum_out[3][3][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][3][5] = (sum_out[4][3][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][3][5] = (sum_out[5][3][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][3][5] = (sum_out[6][3][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][3][5] = (sum_out[7][3][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][3][5] = (sum_out[8][3][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][3][5] = (sum_out[9][3][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][3][5] = (sum_out[10][3][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][3][5] = (sum_out[11][3][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][3][5] = (sum_out[12][3][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][3][5] = (sum_out[13][3][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][3][5] = (sum_out[14][3][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][3][5] = (sum_out[15][3][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][3][5] = (sum_out[16][3][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][3][5] = (sum_out[17][3][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][3][5] = (sum_out[18][3][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][3][5] = (sum_out[19][3][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][3][6] = (sum_out[0][3][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][3][6] = (sum_out[1][3][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][3][6] = (sum_out[2][3][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][3][6] = (sum_out[3][3][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][3][6] = (sum_out[4][3][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][3][6] = (sum_out[5][3][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][3][6] = (sum_out[6][3][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][3][6] = (sum_out[7][3][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][3][6] = (sum_out[8][3][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][3][6] = (sum_out[9][3][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][3][6] = (sum_out[10][3][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][3][6] = (sum_out[11][3][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][3][6] = (sum_out[12][3][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][3][6] = (sum_out[13][3][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][3][6] = (sum_out[14][3][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][3][6] = (sum_out[15][3][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][3][6] = (sum_out[16][3][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][3][6] = (sum_out[17][3][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][3][6] = (sum_out[18][3][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][3][6] = (sum_out[19][3][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][3][7] = (sum_out[0][3][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][3][7] = (sum_out[1][3][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][3][7] = (sum_out[2][3][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][3][7] = (sum_out[3][3][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][3][7] = (sum_out[4][3][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][3][7] = (sum_out[5][3][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][3][7] = (sum_out[6][3][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][3][7] = (sum_out[7][3][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][3][7] = (sum_out[8][3][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][3][7] = (sum_out[9][3][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][3][7] = (sum_out[10][3][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][3][7] = (sum_out[11][3][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][3][7] = (sum_out[12][3][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][3][7] = (sum_out[13][3][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][3][7] = (sum_out[14][3][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][3][7] = (sum_out[15][3][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][3][7] = (sum_out[16][3][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][3][7] = (sum_out[17][3][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][3][7] = (sum_out[18][3][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][3][7] = (sum_out[19][3][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][3][8] = (sum_out[0][3][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][3][8] = (sum_out[1][3][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][3][8] = (sum_out[2][3][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][3][8] = (sum_out[3][3][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][3][8] = (sum_out[4][3][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][3][8] = (sum_out[5][3][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][3][8] = (sum_out[6][3][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][3][8] = (sum_out[7][3][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][3][8] = (sum_out[8][3][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][3][8] = (sum_out[9][3][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][3][8] = (sum_out[10][3][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][3][8] = (sum_out[11][3][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][3][8] = (sum_out[12][3][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][3][8] = (sum_out[13][3][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][3][8] = (sum_out[14][3][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][3][8] = (sum_out[15][3][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][3][8] = (sum_out[16][3][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][3][8] = (sum_out[17][3][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][3][8] = (sum_out[18][3][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][3][8] = (sum_out[19][3][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][3][9] = (sum_out[0][3][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][3][9] = (sum_out[1][3][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][3][9] = (sum_out[2][3][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][3][9] = (sum_out[3][3][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][3][9] = (sum_out[4][3][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][3][9] = (sum_out[5][3][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][3][9] = (sum_out[6][3][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][3][9] = (sum_out[7][3][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][3][9] = (sum_out[8][3][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][3][9] = (sum_out[9][3][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][3][9] = (sum_out[10][3][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][3][9] = (sum_out[11][3][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][3][9] = (sum_out[12][3][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][3][9] = (sum_out[13][3][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][3][9] = (sum_out[14][3][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][3][9] = (sum_out[15][3][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][3][9] = (sum_out[16][3][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][3][9] = (sum_out[17][3][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][3][9] = (sum_out[18][3][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][3][9] = (sum_out[19][3][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][3][10] = (sum_out[0][3][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][3][10] = (sum_out[1][3][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][3][10] = (sum_out[2][3][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][3][10] = (sum_out[3][3][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][3][10] = (sum_out[4][3][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][3][10] = (sum_out[5][3][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][3][10] = (sum_out[6][3][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][3][10] = (sum_out[7][3][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][3][10] = (sum_out[8][3][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][3][10] = (sum_out[9][3][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][3][10] = (sum_out[10][3][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][3][10] = (sum_out[11][3][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][3][10] = (sum_out[12][3][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][3][10] = (sum_out[13][3][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][3][10] = (sum_out[14][3][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][3][10] = (sum_out[15][3][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][3][10] = (sum_out[16][3][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][3][10] = (sum_out[17][3][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][3][10] = (sum_out[18][3][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][3][10] = (sum_out[19][3][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][3][11] = (sum_out[0][3][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][3][11] = (sum_out[1][3][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][3][11] = (sum_out[2][3][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][3][11] = (sum_out[3][3][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][3][11] = (sum_out[4][3][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][3][11] = (sum_out[5][3][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][3][11] = (sum_out[6][3][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][3][11] = (sum_out[7][3][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][3][11] = (sum_out[8][3][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][3][11] = (sum_out[9][3][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][3][11] = (sum_out[10][3][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][3][11] = (sum_out[11][3][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][3][11] = (sum_out[12][3][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][3][11] = (sum_out[13][3][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][3][11] = (sum_out[14][3][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][3][11] = (sum_out[15][3][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][3][11] = (sum_out[16][3][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][3][11] = (sum_out[17][3][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][3][11] = (sum_out[18][3][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][3][11] = (sum_out[19][3][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][3][12] = (sum_out[0][3][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][3][12] = (sum_out[1][3][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][3][12] = (sum_out[2][3][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][3][12] = (sum_out[3][3][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][3][12] = (sum_out[4][3][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][3][12] = (sum_out[5][3][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][3][12] = (sum_out[6][3][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][3][12] = (sum_out[7][3][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][3][12] = (sum_out[8][3][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][3][12] = (sum_out[9][3][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][3][12] = (sum_out[10][3][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][3][12] = (sum_out[11][3][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][3][12] = (sum_out[12][3][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][3][12] = (sum_out[13][3][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][3][12] = (sum_out[14][3][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][3][12] = (sum_out[15][3][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][3][12] = (sum_out[16][3][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][3][12] = (sum_out[17][3][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][3][12] = (sum_out[18][3][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][3][12] = (sum_out[19][3][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][3][13] = (sum_out[0][3][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][3][13] = (sum_out[1][3][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][3][13] = (sum_out[2][3][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][3][13] = (sum_out[3][3][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][3][13] = (sum_out[4][3][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][3][13] = (sum_out[5][3][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][3][13] = (sum_out[6][3][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][3][13] = (sum_out[7][3][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][3][13] = (sum_out[8][3][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][3][13] = (sum_out[9][3][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][3][13] = (sum_out[10][3][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][3][13] = (sum_out[11][3][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][3][13] = (sum_out[12][3][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][3][13] = (sum_out[13][3][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][3][13] = (sum_out[14][3][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][3][13] = (sum_out[15][3][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][3][13] = (sum_out[16][3][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][3][13] = (sum_out[17][3][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][3][13] = (sum_out[18][3][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][3][13] = (sum_out[19][3][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][3][14] = (sum_out[0][3][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][3][14] = (sum_out[1][3][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][3][14] = (sum_out[2][3][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][3][14] = (sum_out[3][3][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][3][14] = (sum_out[4][3][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][3][14] = (sum_out[5][3][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][3][14] = (sum_out[6][3][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][3][14] = (sum_out[7][3][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][3][14] = (sum_out[8][3][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][3][14] = (sum_out[9][3][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][3][14] = (sum_out[10][3][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][3][14] = (sum_out[11][3][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][3][14] = (sum_out[12][3][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][3][14] = (sum_out[13][3][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][3][14] = (sum_out[14][3][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][3][14] = (sum_out[15][3][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][3][14] = (sum_out[16][3][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][3][14] = (sum_out[17][3][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][3][14] = (sum_out[18][3][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][3][14] = (sum_out[19][3][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][3][15] = (sum_out[0][3][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][3][15] = (sum_out[1][3][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][3][15] = (sum_out[2][3][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][3][15] = (sum_out[3][3][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][3][15] = (sum_out[4][3][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][3][15] = (sum_out[5][3][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][3][15] = (sum_out[6][3][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][3][15] = (sum_out[7][3][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][3][15] = (sum_out[8][3][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][3][15] = (sum_out[9][3][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][3][15] = (sum_out[10][3][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][3][15] = (sum_out[11][3][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][3][15] = (sum_out[12][3][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][3][15] = (sum_out[13][3][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][3][15] = (sum_out[14][3][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][3][15] = (sum_out[15][3][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][3][15] = (sum_out[16][3][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][3][15] = (sum_out[17][3][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][3][15] = (sum_out[18][3][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][3][15] = (sum_out[19][3][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][3][16] = (sum_out[0][3][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][3][16] = (sum_out[1][3][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][3][16] = (sum_out[2][3][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][3][16] = (sum_out[3][3][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][3][16] = (sum_out[4][3][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][3][16] = (sum_out[5][3][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][3][16] = (sum_out[6][3][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][3][16] = (sum_out[7][3][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][3][16] = (sum_out[8][3][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][3][16] = (sum_out[9][3][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][3][16] = (sum_out[10][3][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][3][16] = (sum_out[11][3][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][3][16] = (sum_out[12][3][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][3][16] = (sum_out[13][3][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][3][16] = (sum_out[14][3][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][3][16] = (sum_out[15][3][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][3][16] = (sum_out[16][3][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][3][16] = (sum_out[17][3][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][3][16] = (sum_out[18][3][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][3][16] = (sum_out[19][3][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][3][17] = (sum_out[0][3][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][3][17] = (sum_out[1][3][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][3][17] = (sum_out[2][3][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][3][17] = (sum_out[3][3][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][3][17] = (sum_out[4][3][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][3][17] = (sum_out[5][3][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][3][17] = (sum_out[6][3][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][3][17] = (sum_out[7][3][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][3][17] = (sum_out[8][3][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][3][17] = (sum_out[9][3][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][3][17] = (sum_out[10][3][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][3][17] = (sum_out[11][3][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][3][17] = (sum_out[12][3][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][3][17] = (sum_out[13][3][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][3][17] = (sum_out[14][3][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][3][17] = (sum_out[15][3][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][3][17] = (sum_out[16][3][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][3][17] = (sum_out[17][3][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][3][17] = (sum_out[18][3][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][3][17] = (sum_out[19][3][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][3][18] = (sum_out[0][3][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][3][18] = (sum_out[1][3][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][3][18] = (sum_out[2][3][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][3][18] = (sum_out[3][3][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][3][18] = (sum_out[4][3][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][3][18] = (sum_out[5][3][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][3][18] = (sum_out[6][3][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][3][18] = (sum_out[7][3][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][3][18] = (sum_out[8][3][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][3][18] = (sum_out[9][3][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][3][18] = (sum_out[10][3][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][3][18] = (sum_out[11][3][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][3][18] = (sum_out[12][3][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][3][18] = (sum_out[13][3][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][3][18] = (sum_out[14][3][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][3][18] = (sum_out[15][3][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][3][18] = (sum_out[16][3][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][3][18] = (sum_out[17][3][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][3][18] = (sum_out[18][3][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][3][18] = (sum_out[19][3][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][3][19] = (sum_out[0][3][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][3][19] = (sum_out[1][3][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][3][19] = (sum_out[2][3][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][3][19] = (sum_out[3][3][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][3][19] = (sum_out[4][3][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][3][19] = (sum_out[5][3][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][3][19] = (sum_out[6][3][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][3][19] = (sum_out[7][3][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][3][19] = (sum_out[8][3][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][3][19] = (sum_out[9][3][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][3][19] = (sum_out[10][3][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][3][19] = (sum_out[11][3][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][3][19] = (sum_out[12][3][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][3][19] = (sum_out[13][3][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][3][19] = (sum_out[14][3][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][3][19] = (sum_out[15][3][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][3][19] = (sum_out[16][3][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][3][19] = (sum_out[17][3][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][3][19] = (sum_out[18][3][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][3][19] = (sum_out[19][3][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][3][20] = (sum_out[0][3][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][3][20] = (sum_out[1][3][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][3][20] = (sum_out[2][3][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][3][20] = (sum_out[3][3][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][3][20] = (sum_out[4][3][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][3][20] = (sum_out[5][3][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][3][20] = (sum_out[6][3][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][3][20] = (sum_out[7][3][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][3][20] = (sum_out[8][3][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][3][20] = (sum_out[9][3][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][3][20] = (sum_out[10][3][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][3][20] = (sum_out[11][3][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][3][20] = (sum_out[12][3][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][3][20] = (sum_out[13][3][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][3][20] = (sum_out[14][3][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][3][20] = (sum_out[15][3][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][3][20] = (sum_out[16][3][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][3][20] = (sum_out[17][3][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][3][20] = (sum_out[18][3][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][3][20] = (sum_out[19][3][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][3][21] = (sum_out[0][3][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][3][21] = (sum_out[1][3][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][3][21] = (sum_out[2][3][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][3][21] = (sum_out[3][3][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][3][21] = (sum_out[4][3][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][3][21] = (sum_out[5][3][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][3][21] = (sum_out[6][3][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][3][21] = (sum_out[7][3][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][3][21] = (sum_out[8][3][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][3][21] = (sum_out[9][3][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][3][21] = (sum_out[10][3][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][3][21] = (sum_out[11][3][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][3][21] = (sum_out[12][3][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][3][21] = (sum_out[13][3][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][3][21] = (sum_out[14][3][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][3][21] = (sum_out[15][3][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][3][21] = (sum_out[16][3][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][3][21] = (sum_out[17][3][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][3][21] = (sum_out[18][3][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][3][21] = (sum_out[19][3][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][3][22] = (sum_out[0][3][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][3][22] = (sum_out[1][3][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][3][22] = (sum_out[2][3][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][3][22] = (sum_out[3][3][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][3][22] = (sum_out[4][3][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][3][22] = (sum_out[5][3][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][3][22] = (sum_out[6][3][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][3][22] = (sum_out[7][3][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][3][22] = (sum_out[8][3][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][3][22] = (sum_out[9][3][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][3][22] = (sum_out[10][3][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][3][22] = (sum_out[11][3][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][3][22] = (sum_out[12][3][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][3][22] = (sum_out[13][3][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][3][22] = (sum_out[14][3][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][3][22] = (sum_out[15][3][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][3][22] = (sum_out[16][3][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][3][22] = (sum_out[17][3][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][3][22] = (sum_out[18][3][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][3][22] = (sum_out[19][3][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][3][23] = (sum_out[0][3][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][3][23] = (sum_out[1][3][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][3][23] = (sum_out[2][3][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][3][23] = (sum_out[3][3][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][3][23] = (sum_out[4][3][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][3][23] = (sum_out[5][3][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][3][23] = (sum_out[6][3][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][3][23] = (sum_out[7][3][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][3][23] = (sum_out[8][3][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][3][23] = (sum_out[9][3][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][3][23] = (sum_out[10][3][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][3][23] = (sum_out[11][3][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][3][23] = (sum_out[12][3][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][3][23] = (sum_out[13][3][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][3][23] = (sum_out[14][3][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][3][23] = (sum_out[15][3][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][3][23] = (sum_out[16][3][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][3][23] = (sum_out[17][3][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][3][23] = (sum_out[18][3][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][3][23] = (sum_out[19][3][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][4][0] = (sum_out[0][4][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][4][0] = (sum_out[1][4][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][4][0] = (sum_out[2][4][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][4][0] = (sum_out[3][4][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][4][0] = (sum_out[4][4][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][4][0] = (sum_out[5][4][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][4][0] = (sum_out[6][4][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][4][0] = (sum_out[7][4][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][4][0] = (sum_out[8][4][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][4][0] = (sum_out[9][4][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][4][0] = (sum_out[10][4][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][4][0] = (sum_out[11][4][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][4][0] = (sum_out[12][4][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][4][0] = (sum_out[13][4][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][4][0] = (sum_out[14][4][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][4][0] = (sum_out[15][4][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][4][0] = (sum_out[16][4][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][4][0] = (sum_out[17][4][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][4][0] = (sum_out[18][4][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][4][0] = (sum_out[19][4][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][4][1] = (sum_out[0][4][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][4][1] = (sum_out[1][4][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][4][1] = (sum_out[2][4][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][4][1] = (sum_out[3][4][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][4][1] = (sum_out[4][4][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][4][1] = (sum_out[5][4][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][4][1] = (sum_out[6][4][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][4][1] = (sum_out[7][4][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][4][1] = (sum_out[8][4][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][4][1] = (sum_out[9][4][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][4][1] = (sum_out[10][4][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][4][1] = (sum_out[11][4][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][4][1] = (sum_out[12][4][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][4][1] = (sum_out[13][4][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][4][1] = (sum_out[14][4][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][4][1] = (sum_out[15][4][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][4][1] = (sum_out[16][4][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][4][1] = (sum_out[17][4][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][4][1] = (sum_out[18][4][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][4][1] = (sum_out[19][4][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][4][2] = (sum_out[0][4][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][4][2] = (sum_out[1][4][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][4][2] = (sum_out[2][4][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][4][2] = (sum_out[3][4][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][4][2] = (sum_out[4][4][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][4][2] = (sum_out[5][4][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][4][2] = (sum_out[6][4][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][4][2] = (sum_out[7][4][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][4][2] = (sum_out[8][4][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][4][2] = (sum_out[9][4][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][4][2] = (sum_out[10][4][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][4][2] = (sum_out[11][4][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][4][2] = (sum_out[12][4][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][4][2] = (sum_out[13][4][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][4][2] = (sum_out[14][4][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][4][2] = (sum_out[15][4][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][4][2] = (sum_out[16][4][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][4][2] = (sum_out[17][4][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][4][2] = (sum_out[18][4][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][4][2] = (sum_out[19][4][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][4][3] = (sum_out[0][4][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][4][3] = (sum_out[1][4][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][4][3] = (sum_out[2][4][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][4][3] = (sum_out[3][4][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][4][3] = (sum_out[4][4][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][4][3] = (sum_out[5][4][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][4][3] = (sum_out[6][4][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][4][3] = (sum_out[7][4][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][4][3] = (sum_out[8][4][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][4][3] = (sum_out[9][4][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][4][3] = (sum_out[10][4][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][4][3] = (sum_out[11][4][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][4][3] = (sum_out[12][4][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][4][3] = (sum_out[13][4][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][4][3] = (sum_out[14][4][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][4][3] = (sum_out[15][4][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][4][3] = (sum_out[16][4][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][4][3] = (sum_out[17][4][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][4][3] = (sum_out[18][4][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][4][3] = (sum_out[19][4][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][4][4] = (sum_out[0][4][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][4][4] = (sum_out[1][4][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][4][4] = (sum_out[2][4][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][4][4] = (sum_out[3][4][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][4][4] = (sum_out[4][4][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][4][4] = (sum_out[5][4][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][4][4] = (sum_out[6][4][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][4][4] = (sum_out[7][4][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][4][4] = (sum_out[8][4][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][4][4] = (sum_out[9][4][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][4][4] = (sum_out[10][4][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][4][4] = (sum_out[11][4][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][4][4] = (sum_out[12][4][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][4][4] = (sum_out[13][4][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][4][4] = (sum_out[14][4][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][4][4] = (sum_out[15][4][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][4][4] = (sum_out[16][4][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][4][4] = (sum_out[17][4][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][4][4] = (sum_out[18][4][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][4][4] = (sum_out[19][4][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][4][5] = (sum_out[0][4][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][4][5] = (sum_out[1][4][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][4][5] = (sum_out[2][4][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][4][5] = (sum_out[3][4][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][4][5] = (sum_out[4][4][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][4][5] = (sum_out[5][4][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][4][5] = (sum_out[6][4][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][4][5] = (sum_out[7][4][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][4][5] = (sum_out[8][4][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][4][5] = (sum_out[9][4][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][4][5] = (sum_out[10][4][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][4][5] = (sum_out[11][4][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][4][5] = (sum_out[12][4][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][4][5] = (sum_out[13][4][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][4][5] = (sum_out[14][4][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][4][5] = (sum_out[15][4][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][4][5] = (sum_out[16][4][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][4][5] = (sum_out[17][4][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][4][5] = (sum_out[18][4][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][4][5] = (sum_out[19][4][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][4][6] = (sum_out[0][4][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][4][6] = (sum_out[1][4][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][4][6] = (sum_out[2][4][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][4][6] = (sum_out[3][4][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][4][6] = (sum_out[4][4][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][4][6] = (sum_out[5][4][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][4][6] = (sum_out[6][4][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][4][6] = (sum_out[7][4][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][4][6] = (sum_out[8][4][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][4][6] = (sum_out[9][4][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][4][6] = (sum_out[10][4][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][4][6] = (sum_out[11][4][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][4][6] = (sum_out[12][4][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][4][6] = (sum_out[13][4][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][4][6] = (sum_out[14][4][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][4][6] = (sum_out[15][4][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][4][6] = (sum_out[16][4][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][4][6] = (sum_out[17][4][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][4][6] = (sum_out[18][4][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][4][6] = (sum_out[19][4][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][4][7] = (sum_out[0][4][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][4][7] = (sum_out[1][4][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][4][7] = (sum_out[2][4][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][4][7] = (sum_out[3][4][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][4][7] = (sum_out[4][4][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][4][7] = (sum_out[5][4][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][4][7] = (sum_out[6][4][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][4][7] = (sum_out[7][4][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][4][7] = (sum_out[8][4][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][4][7] = (sum_out[9][4][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][4][7] = (sum_out[10][4][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][4][7] = (sum_out[11][4][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][4][7] = (sum_out[12][4][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][4][7] = (sum_out[13][4][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][4][7] = (sum_out[14][4][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][4][7] = (sum_out[15][4][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][4][7] = (sum_out[16][4][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][4][7] = (sum_out[17][4][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][4][7] = (sum_out[18][4][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][4][7] = (sum_out[19][4][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][4][8] = (sum_out[0][4][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][4][8] = (sum_out[1][4][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][4][8] = (sum_out[2][4][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][4][8] = (sum_out[3][4][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][4][8] = (sum_out[4][4][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][4][8] = (sum_out[5][4][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][4][8] = (sum_out[6][4][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][4][8] = (sum_out[7][4][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][4][8] = (sum_out[8][4][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][4][8] = (sum_out[9][4][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][4][8] = (sum_out[10][4][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][4][8] = (sum_out[11][4][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][4][8] = (sum_out[12][4][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][4][8] = (sum_out[13][4][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][4][8] = (sum_out[14][4][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][4][8] = (sum_out[15][4][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][4][8] = (sum_out[16][4][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][4][8] = (sum_out[17][4][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][4][8] = (sum_out[18][4][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][4][8] = (sum_out[19][4][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][4][9] = (sum_out[0][4][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][4][9] = (sum_out[1][4][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][4][9] = (sum_out[2][4][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][4][9] = (sum_out[3][4][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][4][9] = (sum_out[4][4][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][4][9] = (sum_out[5][4][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][4][9] = (sum_out[6][4][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][4][9] = (sum_out[7][4][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][4][9] = (sum_out[8][4][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][4][9] = (sum_out[9][4][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][4][9] = (sum_out[10][4][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][4][9] = (sum_out[11][4][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][4][9] = (sum_out[12][4][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][4][9] = (sum_out[13][4][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][4][9] = (sum_out[14][4][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][4][9] = (sum_out[15][4][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][4][9] = (sum_out[16][4][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][4][9] = (sum_out[17][4][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][4][9] = (sum_out[18][4][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][4][9] = (sum_out[19][4][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][4][10] = (sum_out[0][4][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][4][10] = (sum_out[1][4][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][4][10] = (sum_out[2][4][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][4][10] = (sum_out[3][4][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][4][10] = (sum_out[4][4][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][4][10] = (sum_out[5][4][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][4][10] = (sum_out[6][4][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][4][10] = (sum_out[7][4][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][4][10] = (sum_out[8][4][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][4][10] = (sum_out[9][4][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][4][10] = (sum_out[10][4][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][4][10] = (sum_out[11][4][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][4][10] = (sum_out[12][4][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][4][10] = (sum_out[13][4][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][4][10] = (sum_out[14][4][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][4][10] = (sum_out[15][4][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][4][10] = (sum_out[16][4][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][4][10] = (sum_out[17][4][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][4][10] = (sum_out[18][4][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][4][10] = (sum_out[19][4][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][4][11] = (sum_out[0][4][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][4][11] = (sum_out[1][4][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][4][11] = (sum_out[2][4][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][4][11] = (sum_out[3][4][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][4][11] = (sum_out[4][4][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][4][11] = (sum_out[5][4][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][4][11] = (sum_out[6][4][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][4][11] = (sum_out[7][4][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][4][11] = (sum_out[8][4][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][4][11] = (sum_out[9][4][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][4][11] = (sum_out[10][4][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][4][11] = (sum_out[11][4][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][4][11] = (sum_out[12][4][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][4][11] = (sum_out[13][4][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][4][11] = (sum_out[14][4][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][4][11] = (sum_out[15][4][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][4][11] = (sum_out[16][4][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][4][11] = (sum_out[17][4][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][4][11] = (sum_out[18][4][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][4][11] = (sum_out[19][4][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][4][12] = (sum_out[0][4][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][4][12] = (sum_out[1][4][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][4][12] = (sum_out[2][4][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][4][12] = (sum_out[3][4][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][4][12] = (sum_out[4][4][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][4][12] = (sum_out[5][4][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][4][12] = (sum_out[6][4][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][4][12] = (sum_out[7][4][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][4][12] = (sum_out[8][4][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][4][12] = (sum_out[9][4][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][4][12] = (sum_out[10][4][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][4][12] = (sum_out[11][4][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][4][12] = (sum_out[12][4][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][4][12] = (sum_out[13][4][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][4][12] = (sum_out[14][4][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][4][12] = (sum_out[15][4][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][4][12] = (sum_out[16][4][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][4][12] = (sum_out[17][4][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][4][12] = (sum_out[18][4][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][4][12] = (sum_out[19][4][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][4][13] = (sum_out[0][4][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][4][13] = (sum_out[1][4][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][4][13] = (sum_out[2][4][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][4][13] = (sum_out[3][4][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][4][13] = (sum_out[4][4][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][4][13] = (sum_out[5][4][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][4][13] = (sum_out[6][4][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][4][13] = (sum_out[7][4][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][4][13] = (sum_out[8][4][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][4][13] = (sum_out[9][4][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][4][13] = (sum_out[10][4][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][4][13] = (sum_out[11][4][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][4][13] = (sum_out[12][4][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][4][13] = (sum_out[13][4][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][4][13] = (sum_out[14][4][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][4][13] = (sum_out[15][4][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][4][13] = (sum_out[16][4][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][4][13] = (sum_out[17][4][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][4][13] = (sum_out[18][4][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][4][13] = (sum_out[19][4][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][4][14] = (sum_out[0][4][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][4][14] = (sum_out[1][4][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][4][14] = (sum_out[2][4][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][4][14] = (sum_out[3][4][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][4][14] = (sum_out[4][4][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][4][14] = (sum_out[5][4][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][4][14] = (sum_out[6][4][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][4][14] = (sum_out[7][4][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][4][14] = (sum_out[8][4][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][4][14] = (sum_out[9][4][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][4][14] = (sum_out[10][4][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][4][14] = (sum_out[11][4][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][4][14] = (sum_out[12][4][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][4][14] = (sum_out[13][4][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][4][14] = (sum_out[14][4][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][4][14] = (sum_out[15][4][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][4][14] = (sum_out[16][4][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][4][14] = (sum_out[17][4][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][4][14] = (sum_out[18][4][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][4][14] = (sum_out[19][4][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][4][15] = (sum_out[0][4][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][4][15] = (sum_out[1][4][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][4][15] = (sum_out[2][4][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][4][15] = (sum_out[3][4][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][4][15] = (sum_out[4][4][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][4][15] = (sum_out[5][4][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][4][15] = (sum_out[6][4][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][4][15] = (sum_out[7][4][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][4][15] = (sum_out[8][4][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][4][15] = (sum_out[9][4][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][4][15] = (sum_out[10][4][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][4][15] = (sum_out[11][4][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][4][15] = (sum_out[12][4][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][4][15] = (sum_out[13][4][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][4][15] = (sum_out[14][4][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][4][15] = (sum_out[15][4][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][4][15] = (sum_out[16][4][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][4][15] = (sum_out[17][4][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][4][15] = (sum_out[18][4][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][4][15] = (sum_out[19][4][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][4][16] = (sum_out[0][4][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][4][16] = (sum_out[1][4][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][4][16] = (sum_out[2][4][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][4][16] = (sum_out[3][4][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][4][16] = (sum_out[4][4][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][4][16] = (sum_out[5][4][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][4][16] = (sum_out[6][4][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][4][16] = (sum_out[7][4][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][4][16] = (sum_out[8][4][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][4][16] = (sum_out[9][4][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][4][16] = (sum_out[10][4][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][4][16] = (sum_out[11][4][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][4][16] = (sum_out[12][4][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][4][16] = (sum_out[13][4][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][4][16] = (sum_out[14][4][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][4][16] = (sum_out[15][4][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][4][16] = (sum_out[16][4][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][4][16] = (sum_out[17][4][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][4][16] = (sum_out[18][4][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][4][16] = (sum_out[19][4][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][4][17] = (sum_out[0][4][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][4][17] = (sum_out[1][4][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][4][17] = (sum_out[2][4][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][4][17] = (sum_out[3][4][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][4][17] = (sum_out[4][4][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][4][17] = (sum_out[5][4][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][4][17] = (sum_out[6][4][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][4][17] = (sum_out[7][4][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][4][17] = (sum_out[8][4][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][4][17] = (sum_out[9][4][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][4][17] = (sum_out[10][4][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][4][17] = (sum_out[11][4][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][4][17] = (sum_out[12][4][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][4][17] = (sum_out[13][4][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][4][17] = (sum_out[14][4][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][4][17] = (sum_out[15][4][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][4][17] = (sum_out[16][4][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][4][17] = (sum_out[17][4][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][4][17] = (sum_out[18][4][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][4][17] = (sum_out[19][4][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][4][18] = (sum_out[0][4][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][4][18] = (sum_out[1][4][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][4][18] = (sum_out[2][4][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][4][18] = (sum_out[3][4][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][4][18] = (sum_out[4][4][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][4][18] = (sum_out[5][4][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][4][18] = (sum_out[6][4][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][4][18] = (sum_out[7][4][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][4][18] = (sum_out[8][4][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][4][18] = (sum_out[9][4][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][4][18] = (sum_out[10][4][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][4][18] = (sum_out[11][4][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][4][18] = (sum_out[12][4][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][4][18] = (sum_out[13][4][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][4][18] = (sum_out[14][4][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][4][18] = (sum_out[15][4][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][4][18] = (sum_out[16][4][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][4][18] = (sum_out[17][4][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][4][18] = (sum_out[18][4][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][4][18] = (sum_out[19][4][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][4][19] = (sum_out[0][4][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][4][19] = (sum_out[1][4][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][4][19] = (sum_out[2][4][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][4][19] = (sum_out[3][4][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][4][19] = (sum_out[4][4][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][4][19] = (sum_out[5][4][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][4][19] = (sum_out[6][4][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][4][19] = (sum_out[7][4][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][4][19] = (sum_out[8][4][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][4][19] = (sum_out[9][4][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][4][19] = (sum_out[10][4][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][4][19] = (sum_out[11][4][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][4][19] = (sum_out[12][4][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][4][19] = (sum_out[13][4][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][4][19] = (sum_out[14][4][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][4][19] = (sum_out[15][4][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][4][19] = (sum_out[16][4][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][4][19] = (sum_out[17][4][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][4][19] = (sum_out[18][4][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][4][19] = (sum_out[19][4][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][4][20] = (sum_out[0][4][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][4][20] = (sum_out[1][4][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][4][20] = (sum_out[2][4][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][4][20] = (sum_out[3][4][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][4][20] = (sum_out[4][4][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][4][20] = (sum_out[5][4][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][4][20] = (sum_out[6][4][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][4][20] = (sum_out[7][4][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][4][20] = (sum_out[8][4][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][4][20] = (sum_out[9][4][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][4][20] = (sum_out[10][4][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][4][20] = (sum_out[11][4][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][4][20] = (sum_out[12][4][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][4][20] = (sum_out[13][4][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][4][20] = (sum_out[14][4][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][4][20] = (sum_out[15][4][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][4][20] = (sum_out[16][4][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][4][20] = (sum_out[17][4][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][4][20] = (sum_out[18][4][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][4][20] = (sum_out[19][4][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][4][21] = (sum_out[0][4][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][4][21] = (sum_out[1][4][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][4][21] = (sum_out[2][4][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][4][21] = (sum_out[3][4][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][4][21] = (sum_out[4][4][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][4][21] = (sum_out[5][4][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][4][21] = (sum_out[6][4][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][4][21] = (sum_out[7][4][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][4][21] = (sum_out[8][4][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][4][21] = (sum_out[9][4][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][4][21] = (sum_out[10][4][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][4][21] = (sum_out[11][4][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][4][21] = (sum_out[12][4][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][4][21] = (sum_out[13][4][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][4][21] = (sum_out[14][4][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][4][21] = (sum_out[15][4][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][4][21] = (sum_out[16][4][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][4][21] = (sum_out[17][4][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][4][21] = (sum_out[18][4][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][4][21] = (sum_out[19][4][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][4][22] = (sum_out[0][4][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][4][22] = (sum_out[1][4][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][4][22] = (sum_out[2][4][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][4][22] = (sum_out[3][4][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][4][22] = (sum_out[4][4][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][4][22] = (sum_out[5][4][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][4][22] = (sum_out[6][4][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][4][22] = (sum_out[7][4][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][4][22] = (sum_out[8][4][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][4][22] = (sum_out[9][4][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][4][22] = (sum_out[10][4][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][4][22] = (sum_out[11][4][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][4][22] = (sum_out[12][4][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][4][22] = (sum_out[13][4][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][4][22] = (sum_out[14][4][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][4][22] = (sum_out[15][4][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][4][22] = (sum_out[16][4][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][4][22] = (sum_out[17][4][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][4][22] = (sum_out[18][4][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][4][22] = (sum_out[19][4][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][4][23] = (sum_out[0][4][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][4][23] = (sum_out[1][4][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][4][23] = (sum_out[2][4][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][4][23] = (sum_out[3][4][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][4][23] = (sum_out[4][4][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][4][23] = (sum_out[5][4][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][4][23] = (sum_out[6][4][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][4][23] = (sum_out[7][4][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][4][23] = (sum_out[8][4][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][4][23] = (sum_out[9][4][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][4][23] = (sum_out[10][4][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][4][23] = (sum_out[11][4][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][4][23] = (sum_out[12][4][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][4][23] = (sum_out[13][4][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][4][23] = (sum_out[14][4][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][4][23] = (sum_out[15][4][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][4][23] = (sum_out[16][4][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][4][23] = (sum_out[17][4][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][4][23] = (sum_out[18][4][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][4][23] = (sum_out[19][4][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][5][0] = (sum_out[0][5][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][5][0] = (sum_out[1][5][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][5][0] = (sum_out[2][5][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][5][0] = (sum_out[3][5][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][5][0] = (sum_out[4][5][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][5][0] = (sum_out[5][5][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][5][0] = (sum_out[6][5][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][5][0] = (sum_out[7][5][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][5][0] = (sum_out[8][5][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][5][0] = (sum_out[9][5][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][5][0] = (sum_out[10][5][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][5][0] = (sum_out[11][5][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][5][0] = (sum_out[12][5][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][5][0] = (sum_out[13][5][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][5][0] = (sum_out[14][5][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][5][0] = (sum_out[15][5][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][5][0] = (sum_out[16][5][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][5][0] = (sum_out[17][5][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][5][0] = (sum_out[18][5][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][5][0] = (sum_out[19][5][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][5][1] = (sum_out[0][5][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][5][1] = (sum_out[1][5][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][5][1] = (sum_out[2][5][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][5][1] = (sum_out[3][5][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][5][1] = (sum_out[4][5][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][5][1] = (sum_out[5][5][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][5][1] = (sum_out[6][5][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][5][1] = (sum_out[7][5][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][5][1] = (sum_out[8][5][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][5][1] = (sum_out[9][5][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][5][1] = (sum_out[10][5][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][5][1] = (sum_out[11][5][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][5][1] = (sum_out[12][5][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][5][1] = (sum_out[13][5][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][5][1] = (sum_out[14][5][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][5][1] = (sum_out[15][5][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][5][1] = (sum_out[16][5][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][5][1] = (sum_out[17][5][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][5][1] = (sum_out[18][5][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][5][1] = (sum_out[19][5][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][5][2] = (sum_out[0][5][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][5][2] = (sum_out[1][5][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][5][2] = (sum_out[2][5][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][5][2] = (sum_out[3][5][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][5][2] = (sum_out[4][5][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][5][2] = (sum_out[5][5][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][5][2] = (sum_out[6][5][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][5][2] = (sum_out[7][5][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][5][2] = (sum_out[8][5][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][5][2] = (sum_out[9][5][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][5][2] = (sum_out[10][5][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][5][2] = (sum_out[11][5][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][5][2] = (sum_out[12][5][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][5][2] = (sum_out[13][5][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][5][2] = (sum_out[14][5][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][5][2] = (sum_out[15][5][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][5][2] = (sum_out[16][5][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][5][2] = (sum_out[17][5][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][5][2] = (sum_out[18][5][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][5][2] = (sum_out[19][5][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][5][3] = (sum_out[0][5][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][5][3] = (sum_out[1][5][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][5][3] = (sum_out[2][5][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][5][3] = (sum_out[3][5][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][5][3] = (sum_out[4][5][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][5][3] = (sum_out[5][5][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][5][3] = (sum_out[6][5][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][5][3] = (sum_out[7][5][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][5][3] = (sum_out[8][5][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][5][3] = (sum_out[9][5][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][5][3] = (sum_out[10][5][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][5][3] = (sum_out[11][5][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][5][3] = (sum_out[12][5][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][5][3] = (sum_out[13][5][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][5][3] = (sum_out[14][5][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][5][3] = (sum_out[15][5][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][5][3] = (sum_out[16][5][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][5][3] = (sum_out[17][5][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][5][3] = (sum_out[18][5][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][5][3] = (sum_out[19][5][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][5][4] = (sum_out[0][5][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][5][4] = (sum_out[1][5][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][5][4] = (sum_out[2][5][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][5][4] = (sum_out[3][5][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][5][4] = (sum_out[4][5][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][5][4] = (sum_out[5][5][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][5][4] = (sum_out[6][5][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][5][4] = (sum_out[7][5][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][5][4] = (sum_out[8][5][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][5][4] = (sum_out[9][5][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][5][4] = (sum_out[10][5][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][5][4] = (sum_out[11][5][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][5][4] = (sum_out[12][5][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][5][4] = (sum_out[13][5][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][5][4] = (sum_out[14][5][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][5][4] = (sum_out[15][5][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][5][4] = (sum_out[16][5][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][5][4] = (sum_out[17][5][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][5][4] = (sum_out[18][5][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][5][4] = (sum_out[19][5][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][5][5] = (sum_out[0][5][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][5][5] = (sum_out[1][5][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][5][5] = (sum_out[2][5][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][5][5] = (sum_out[3][5][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][5][5] = (sum_out[4][5][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][5][5] = (sum_out[5][5][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][5][5] = (sum_out[6][5][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][5][5] = (sum_out[7][5][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][5][5] = (sum_out[8][5][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][5][5] = (sum_out[9][5][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][5][5] = (sum_out[10][5][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][5][5] = (sum_out[11][5][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][5][5] = (sum_out[12][5][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][5][5] = (sum_out[13][5][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][5][5] = (sum_out[14][5][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][5][5] = (sum_out[15][5][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][5][5] = (sum_out[16][5][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][5][5] = (sum_out[17][5][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][5][5] = (sum_out[18][5][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][5][5] = (sum_out[19][5][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][5][6] = (sum_out[0][5][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][5][6] = (sum_out[1][5][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][5][6] = (sum_out[2][5][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][5][6] = (sum_out[3][5][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][5][6] = (sum_out[4][5][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][5][6] = (sum_out[5][5][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][5][6] = (sum_out[6][5][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][5][6] = (sum_out[7][5][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][5][6] = (sum_out[8][5][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][5][6] = (sum_out[9][5][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][5][6] = (sum_out[10][5][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][5][6] = (sum_out[11][5][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][5][6] = (sum_out[12][5][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][5][6] = (sum_out[13][5][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][5][6] = (sum_out[14][5][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][5][6] = (sum_out[15][5][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][5][6] = (sum_out[16][5][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][5][6] = (sum_out[17][5][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][5][6] = (sum_out[18][5][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][5][6] = (sum_out[19][5][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][5][7] = (sum_out[0][5][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][5][7] = (sum_out[1][5][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][5][7] = (sum_out[2][5][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][5][7] = (sum_out[3][5][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][5][7] = (sum_out[4][5][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][5][7] = (sum_out[5][5][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][5][7] = (sum_out[6][5][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][5][7] = (sum_out[7][5][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][5][7] = (sum_out[8][5][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][5][7] = (sum_out[9][5][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][5][7] = (sum_out[10][5][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][5][7] = (sum_out[11][5][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][5][7] = (sum_out[12][5][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][5][7] = (sum_out[13][5][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][5][7] = (sum_out[14][5][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][5][7] = (sum_out[15][5][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][5][7] = (sum_out[16][5][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][5][7] = (sum_out[17][5][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][5][7] = (sum_out[18][5][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][5][7] = (sum_out[19][5][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][5][8] = (sum_out[0][5][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][5][8] = (sum_out[1][5][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][5][8] = (sum_out[2][5][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][5][8] = (sum_out[3][5][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][5][8] = (sum_out[4][5][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][5][8] = (sum_out[5][5][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][5][8] = (sum_out[6][5][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][5][8] = (sum_out[7][5][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][5][8] = (sum_out[8][5][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][5][8] = (sum_out[9][5][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][5][8] = (sum_out[10][5][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][5][8] = (sum_out[11][5][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][5][8] = (sum_out[12][5][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][5][8] = (sum_out[13][5][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][5][8] = (sum_out[14][5][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][5][8] = (sum_out[15][5][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][5][8] = (sum_out[16][5][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][5][8] = (sum_out[17][5][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][5][8] = (sum_out[18][5][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][5][8] = (sum_out[19][5][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][5][9] = (sum_out[0][5][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][5][9] = (sum_out[1][5][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][5][9] = (sum_out[2][5][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][5][9] = (sum_out[3][5][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][5][9] = (sum_out[4][5][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][5][9] = (sum_out[5][5][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][5][9] = (sum_out[6][5][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][5][9] = (sum_out[7][5][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][5][9] = (sum_out[8][5][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][5][9] = (sum_out[9][5][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][5][9] = (sum_out[10][5][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][5][9] = (sum_out[11][5][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][5][9] = (sum_out[12][5][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][5][9] = (sum_out[13][5][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][5][9] = (sum_out[14][5][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][5][9] = (sum_out[15][5][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][5][9] = (sum_out[16][5][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][5][9] = (sum_out[17][5][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][5][9] = (sum_out[18][5][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][5][9] = (sum_out[19][5][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][5][10] = (sum_out[0][5][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][5][10] = (sum_out[1][5][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][5][10] = (sum_out[2][5][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][5][10] = (sum_out[3][5][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][5][10] = (sum_out[4][5][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][5][10] = (sum_out[5][5][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][5][10] = (sum_out[6][5][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][5][10] = (sum_out[7][5][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][5][10] = (sum_out[8][5][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][5][10] = (sum_out[9][5][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][5][10] = (sum_out[10][5][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][5][10] = (sum_out[11][5][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][5][10] = (sum_out[12][5][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][5][10] = (sum_out[13][5][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][5][10] = (sum_out[14][5][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][5][10] = (sum_out[15][5][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][5][10] = (sum_out[16][5][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][5][10] = (sum_out[17][5][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][5][10] = (sum_out[18][5][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][5][10] = (sum_out[19][5][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][5][11] = (sum_out[0][5][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][5][11] = (sum_out[1][5][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][5][11] = (sum_out[2][5][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][5][11] = (sum_out[3][5][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][5][11] = (sum_out[4][5][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][5][11] = (sum_out[5][5][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][5][11] = (sum_out[6][5][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][5][11] = (sum_out[7][5][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][5][11] = (sum_out[8][5][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][5][11] = (sum_out[9][5][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][5][11] = (sum_out[10][5][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][5][11] = (sum_out[11][5][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][5][11] = (sum_out[12][5][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][5][11] = (sum_out[13][5][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][5][11] = (sum_out[14][5][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][5][11] = (sum_out[15][5][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][5][11] = (sum_out[16][5][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][5][11] = (sum_out[17][5][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][5][11] = (sum_out[18][5][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][5][11] = (sum_out[19][5][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][5][12] = (sum_out[0][5][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][5][12] = (sum_out[1][5][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][5][12] = (sum_out[2][5][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][5][12] = (sum_out[3][5][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][5][12] = (sum_out[4][5][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][5][12] = (sum_out[5][5][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][5][12] = (sum_out[6][5][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][5][12] = (sum_out[7][5][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][5][12] = (sum_out[8][5][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][5][12] = (sum_out[9][5][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][5][12] = (sum_out[10][5][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][5][12] = (sum_out[11][5][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][5][12] = (sum_out[12][5][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][5][12] = (sum_out[13][5][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][5][12] = (sum_out[14][5][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][5][12] = (sum_out[15][5][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][5][12] = (sum_out[16][5][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][5][12] = (sum_out[17][5][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][5][12] = (sum_out[18][5][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][5][12] = (sum_out[19][5][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][5][13] = (sum_out[0][5][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][5][13] = (sum_out[1][5][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][5][13] = (sum_out[2][5][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][5][13] = (sum_out[3][5][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][5][13] = (sum_out[4][5][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][5][13] = (sum_out[5][5][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][5][13] = (sum_out[6][5][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][5][13] = (sum_out[7][5][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][5][13] = (sum_out[8][5][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][5][13] = (sum_out[9][5][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][5][13] = (sum_out[10][5][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][5][13] = (sum_out[11][5][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][5][13] = (sum_out[12][5][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][5][13] = (sum_out[13][5][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][5][13] = (sum_out[14][5][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][5][13] = (sum_out[15][5][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][5][13] = (sum_out[16][5][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][5][13] = (sum_out[17][5][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][5][13] = (sum_out[18][5][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][5][13] = (sum_out[19][5][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][5][14] = (sum_out[0][5][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][5][14] = (sum_out[1][5][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][5][14] = (sum_out[2][5][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][5][14] = (sum_out[3][5][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][5][14] = (sum_out[4][5][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][5][14] = (sum_out[5][5][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][5][14] = (sum_out[6][5][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][5][14] = (sum_out[7][5][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][5][14] = (sum_out[8][5][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][5][14] = (sum_out[9][5][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][5][14] = (sum_out[10][5][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][5][14] = (sum_out[11][5][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][5][14] = (sum_out[12][5][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][5][14] = (sum_out[13][5][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][5][14] = (sum_out[14][5][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][5][14] = (sum_out[15][5][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][5][14] = (sum_out[16][5][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][5][14] = (sum_out[17][5][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][5][14] = (sum_out[18][5][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][5][14] = (sum_out[19][5][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][5][15] = (sum_out[0][5][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][5][15] = (sum_out[1][5][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][5][15] = (sum_out[2][5][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][5][15] = (sum_out[3][5][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][5][15] = (sum_out[4][5][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][5][15] = (sum_out[5][5][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][5][15] = (sum_out[6][5][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][5][15] = (sum_out[7][5][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][5][15] = (sum_out[8][5][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][5][15] = (sum_out[9][5][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][5][15] = (sum_out[10][5][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][5][15] = (sum_out[11][5][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][5][15] = (sum_out[12][5][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][5][15] = (sum_out[13][5][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][5][15] = (sum_out[14][5][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][5][15] = (sum_out[15][5][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][5][15] = (sum_out[16][5][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][5][15] = (sum_out[17][5][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][5][15] = (sum_out[18][5][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][5][15] = (sum_out[19][5][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][5][16] = (sum_out[0][5][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][5][16] = (sum_out[1][5][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][5][16] = (sum_out[2][5][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][5][16] = (sum_out[3][5][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][5][16] = (sum_out[4][5][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][5][16] = (sum_out[5][5][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][5][16] = (sum_out[6][5][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][5][16] = (sum_out[7][5][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][5][16] = (sum_out[8][5][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][5][16] = (sum_out[9][5][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][5][16] = (sum_out[10][5][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][5][16] = (sum_out[11][5][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][5][16] = (sum_out[12][5][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][5][16] = (sum_out[13][5][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][5][16] = (sum_out[14][5][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][5][16] = (sum_out[15][5][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][5][16] = (sum_out[16][5][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][5][16] = (sum_out[17][5][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][5][16] = (sum_out[18][5][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][5][16] = (sum_out[19][5][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][5][17] = (sum_out[0][5][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][5][17] = (sum_out[1][5][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][5][17] = (sum_out[2][5][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][5][17] = (sum_out[3][5][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][5][17] = (sum_out[4][5][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][5][17] = (sum_out[5][5][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][5][17] = (sum_out[6][5][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][5][17] = (sum_out[7][5][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][5][17] = (sum_out[8][5][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][5][17] = (sum_out[9][5][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][5][17] = (sum_out[10][5][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][5][17] = (sum_out[11][5][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][5][17] = (sum_out[12][5][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][5][17] = (sum_out[13][5][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][5][17] = (sum_out[14][5][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][5][17] = (sum_out[15][5][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][5][17] = (sum_out[16][5][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][5][17] = (sum_out[17][5][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][5][17] = (sum_out[18][5][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][5][17] = (sum_out[19][5][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][5][18] = (sum_out[0][5][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][5][18] = (sum_out[1][5][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][5][18] = (sum_out[2][5][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][5][18] = (sum_out[3][5][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][5][18] = (sum_out[4][5][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][5][18] = (sum_out[5][5][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][5][18] = (sum_out[6][5][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][5][18] = (sum_out[7][5][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][5][18] = (sum_out[8][5][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][5][18] = (sum_out[9][5][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][5][18] = (sum_out[10][5][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][5][18] = (sum_out[11][5][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][5][18] = (sum_out[12][5][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][5][18] = (sum_out[13][5][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][5][18] = (sum_out[14][5][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][5][18] = (sum_out[15][5][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][5][18] = (sum_out[16][5][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][5][18] = (sum_out[17][5][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][5][18] = (sum_out[18][5][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][5][18] = (sum_out[19][5][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][5][19] = (sum_out[0][5][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][5][19] = (sum_out[1][5][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][5][19] = (sum_out[2][5][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][5][19] = (sum_out[3][5][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][5][19] = (sum_out[4][5][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][5][19] = (sum_out[5][5][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][5][19] = (sum_out[6][5][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][5][19] = (sum_out[7][5][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][5][19] = (sum_out[8][5][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][5][19] = (sum_out[9][5][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][5][19] = (sum_out[10][5][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][5][19] = (sum_out[11][5][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][5][19] = (sum_out[12][5][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][5][19] = (sum_out[13][5][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][5][19] = (sum_out[14][5][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][5][19] = (sum_out[15][5][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][5][19] = (sum_out[16][5][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][5][19] = (sum_out[17][5][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][5][19] = (sum_out[18][5][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][5][19] = (sum_out[19][5][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][5][20] = (sum_out[0][5][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][5][20] = (sum_out[1][5][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][5][20] = (sum_out[2][5][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][5][20] = (sum_out[3][5][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][5][20] = (sum_out[4][5][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][5][20] = (sum_out[5][5][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][5][20] = (sum_out[6][5][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][5][20] = (sum_out[7][5][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][5][20] = (sum_out[8][5][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][5][20] = (sum_out[9][5][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][5][20] = (sum_out[10][5][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][5][20] = (sum_out[11][5][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][5][20] = (sum_out[12][5][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][5][20] = (sum_out[13][5][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][5][20] = (sum_out[14][5][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][5][20] = (sum_out[15][5][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][5][20] = (sum_out[16][5][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][5][20] = (sum_out[17][5][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][5][20] = (sum_out[18][5][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][5][20] = (sum_out[19][5][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][5][21] = (sum_out[0][5][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][5][21] = (sum_out[1][5][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][5][21] = (sum_out[2][5][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][5][21] = (sum_out[3][5][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][5][21] = (sum_out[4][5][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][5][21] = (sum_out[5][5][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][5][21] = (sum_out[6][5][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][5][21] = (sum_out[7][5][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][5][21] = (sum_out[8][5][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][5][21] = (sum_out[9][5][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][5][21] = (sum_out[10][5][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][5][21] = (sum_out[11][5][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][5][21] = (sum_out[12][5][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][5][21] = (sum_out[13][5][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][5][21] = (sum_out[14][5][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][5][21] = (sum_out[15][5][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][5][21] = (sum_out[16][5][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][5][21] = (sum_out[17][5][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][5][21] = (sum_out[18][5][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][5][21] = (sum_out[19][5][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][5][22] = (sum_out[0][5][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][5][22] = (sum_out[1][5][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][5][22] = (sum_out[2][5][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][5][22] = (sum_out[3][5][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][5][22] = (sum_out[4][5][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][5][22] = (sum_out[5][5][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][5][22] = (sum_out[6][5][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][5][22] = (sum_out[7][5][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][5][22] = (sum_out[8][5][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][5][22] = (sum_out[9][5][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][5][22] = (sum_out[10][5][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][5][22] = (sum_out[11][5][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][5][22] = (sum_out[12][5][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][5][22] = (sum_out[13][5][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][5][22] = (sum_out[14][5][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][5][22] = (sum_out[15][5][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][5][22] = (sum_out[16][5][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][5][22] = (sum_out[17][5][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][5][22] = (sum_out[18][5][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][5][22] = (sum_out[19][5][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][5][23] = (sum_out[0][5][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][5][23] = (sum_out[1][5][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][5][23] = (sum_out[2][5][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][5][23] = (sum_out[3][5][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][5][23] = (sum_out[4][5][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][5][23] = (sum_out[5][5][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][5][23] = (sum_out[6][5][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][5][23] = (sum_out[7][5][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][5][23] = (sum_out[8][5][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][5][23] = (sum_out[9][5][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][5][23] = (sum_out[10][5][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][5][23] = (sum_out[11][5][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][5][23] = (sum_out[12][5][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][5][23] = (sum_out[13][5][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][5][23] = (sum_out[14][5][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][5][23] = (sum_out[15][5][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][5][23] = (sum_out[16][5][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][5][23] = (sum_out[17][5][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][5][23] = (sum_out[18][5][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][5][23] = (sum_out[19][5][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][6][0] = (sum_out[0][6][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][6][0] = (sum_out[1][6][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][6][0] = (sum_out[2][6][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][6][0] = (sum_out[3][6][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][6][0] = (sum_out[4][6][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][6][0] = (sum_out[5][6][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][6][0] = (sum_out[6][6][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][6][0] = (sum_out[7][6][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][6][0] = (sum_out[8][6][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][6][0] = (sum_out[9][6][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][6][0] = (sum_out[10][6][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][6][0] = (sum_out[11][6][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][6][0] = (sum_out[12][6][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][6][0] = (sum_out[13][6][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][6][0] = (sum_out[14][6][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][6][0] = (sum_out[15][6][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][6][0] = (sum_out[16][6][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][6][0] = (sum_out[17][6][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][6][0] = (sum_out[18][6][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][6][0] = (sum_out[19][6][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][6][1] = (sum_out[0][6][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][6][1] = (sum_out[1][6][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][6][1] = (sum_out[2][6][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][6][1] = (sum_out[3][6][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][6][1] = (sum_out[4][6][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][6][1] = (sum_out[5][6][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][6][1] = (sum_out[6][6][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][6][1] = (sum_out[7][6][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][6][1] = (sum_out[8][6][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][6][1] = (sum_out[9][6][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][6][1] = (sum_out[10][6][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][6][1] = (sum_out[11][6][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][6][1] = (sum_out[12][6][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][6][1] = (sum_out[13][6][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][6][1] = (sum_out[14][6][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][6][1] = (sum_out[15][6][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][6][1] = (sum_out[16][6][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][6][1] = (sum_out[17][6][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][6][1] = (sum_out[18][6][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][6][1] = (sum_out[19][6][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][6][2] = (sum_out[0][6][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][6][2] = (sum_out[1][6][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][6][2] = (sum_out[2][6][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][6][2] = (sum_out[3][6][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][6][2] = (sum_out[4][6][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][6][2] = (sum_out[5][6][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][6][2] = (sum_out[6][6][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][6][2] = (sum_out[7][6][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][6][2] = (sum_out[8][6][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][6][2] = (sum_out[9][6][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][6][2] = (sum_out[10][6][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][6][2] = (sum_out[11][6][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][6][2] = (sum_out[12][6][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][6][2] = (sum_out[13][6][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][6][2] = (sum_out[14][6][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][6][2] = (sum_out[15][6][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][6][2] = (sum_out[16][6][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][6][2] = (sum_out[17][6][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][6][2] = (sum_out[18][6][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][6][2] = (sum_out[19][6][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][6][3] = (sum_out[0][6][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][6][3] = (sum_out[1][6][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][6][3] = (sum_out[2][6][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][6][3] = (sum_out[3][6][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][6][3] = (sum_out[4][6][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][6][3] = (sum_out[5][6][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][6][3] = (sum_out[6][6][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][6][3] = (sum_out[7][6][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][6][3] = (sum_out[8][6][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][6][3] = (sum_out[9][6][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][6][3] = (sum_out[10][6][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][6][3] = (sum_out[11][6][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][6][3] = (sum_out[12][6][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][6][3] = (sum_out[13][6][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][6][3] = (sum_out[14][6][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][6][3] = (sum_out[15][6][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][6][3] = (sum_out[16][6][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][6][3] = (sum_out[17][6][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][6][3] = (sum_out[18][6][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][6][3] = (sum_out[19][6][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][6][4] = (sum_out[0][6][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][6][4] = (sum_out[1][6][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][6][4] = (sum_out[2][6][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][6][4] = (sum_out[3][6][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][6][4] = (sum_out[4][6][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][6][4] = (sum_out[5][6][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][6][4] = (sum_out[6][6][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][6][4] = (sum_out[7][6][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][6][4] = (sum_out[8][6][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][6][4] = (sum_out[9][6][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][6][4] = (sum_out[10][6][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][6][4] = (sum_out[11][6][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][6][4] = (sum_out[12][6][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][6][4] = (sum_out[13][6][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][6][4] = (sum_out[14][6][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][6][4] = (sum_out[15][6][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][6][4] = (sum_out[16][6][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][6][4] = (sum_out[17][6][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][6][4] = (sum_out[18][6][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][6][4] = (sum_out[19][6][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][6][5] = (sum_out[0][6][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][6][5] = (sum_out[1][6][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][6][5] = (sum_out[2][6][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][6][5] = (sum_out[3][6][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][6][5] = (sum_out[4][6][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][6][5] = (sum_out[5][6][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][6][5] = (sum_out[6][6][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][6][5] = (sum_out[7][6][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][6][5] = (sum_out[8][6][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][6][5] = (sum_out[9][6][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][6][5] = (sum_out[10][6][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][6][5] = (sum_out[11][6][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][6][5] = (sum_out[12][6][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][6][5] = (sum_out[13][6][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][6][5] = (sum_out[14][6][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][6][5] = (sum_out[15][6][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][6][5] = (sum_out[16][6][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][6][5] = (sum_out[17][6][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][6][5] = (sum_out[18][6][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][6][5] = (sum_out[19][6][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][6][6] = (sum_out[0][6][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][6][6] = (sum_out[1][6][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][6][6] = (sum_out[2][6][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][6][6] = (sum_out[3][6][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][6][6] = (sum_out[4][6][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][6][6] = (sum_out[5][6][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][6][6] = (sum_out[6][6][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][6][6] = (sum_out[7][6][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][6][6] = (sum_out[8][6][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][6][6] = (sum_out[9][6][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][6][6] = (sum_out[10][6][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][6][6] = (sum_out[11][6][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][6][6] = (sum_out[12][6][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][6][6] = (sum_out[13][6][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][6][6] = (sum_out[14][6][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][6][6] = (sum_out[15][6][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][6][6] = (sum_out[16][6][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][6][6] = (sum_out[17][6][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][6][6] = (sum_out[18][6][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][6][6] = (sum_out[19][6][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][6][7] = (sum_out[0][6][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][6][7] = (sum_out[1][6][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][6][7] = (sum_out[2][6][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][6][7] = (sum_out[3][6][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][6][7] = (sum_out[4][6][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][6][7] = (sum_out[5][6][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][6][7] = (sum_out[6][6][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][6][7] = (sum_out[7][6][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][6][7] = (sum_out[8][6][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][6][7] = (sum_out[9][6][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][6][7] = (sum_out[10][6][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][6][7] = (sum_out[11][6][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][6][7] = (sum_out[12][6][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][6][7] = (sum_out[13][6][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][6][7] = (sum_out[14][6][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][6][7] = (sum_out[15][6][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][6][7] = (sum_out[16][6][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][6][7] = (sum_out[17][6][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][6][7] = (sum_out[18][6][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][6][7] = (sum_out[19][6][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][6][8] = (sum_out[0][6][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][6][8] = (sum_out[1][6][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][6][8] = (sum_out[2][6][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][6][8] = (sum_out[3][6][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][6][8] = (sum_out[4][6][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][6][8] = (sum_out[5][6][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][6][8] = (sum_out[6][6][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][6][8] = (sum_out[7][6][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][6][8] = (sum_out[8][6][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][6][8] = (sum_out[9][6][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][6][8] = (sum_out[10][6][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][6][8] = (sum_out[11][6][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][6][8] = (sum_out[12][6][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][6][8] = (sum_out[13][6][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][6][8] = (sum_out[14][6][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][6][8] = (sum_out[15][6][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][6][8] = (sum_out[16][6][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][6][8] = (sum_out[17][6][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][6][8] = (sum_out[18][6][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][6][8] = (sum_out[19][6][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][6][9] = (sum_out[0][6][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][6][9] = (sum_out[1][6][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][6][9] = (sum_out[2][6][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][6][9] = (sum_out[3][6][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][6][9] = (sum_out[4][6][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][6][9] = (sum_out[5][6][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][6][9] = (sum_out[6][6][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][6][9] = (sum_out[7][6][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][6][9] = (sum_out[8][6][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][6][9] = (sum_out[9][6][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][6][9] = (sum_out[10][6][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][6][9] = (sum_out[11][6][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][6][9] = (sum_out[12][6][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][6][9] = (sum_out[13][6][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][6][9] = (sum_out[14][6][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][6][9] = (sum_out[15][6][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][6][9] = (sum_out[16][6][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][6][9] = (sum_out[17][6][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][6][9] = (sum_out[18][6][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][6][9] = (sum_out[19][6][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][6][10] = (sum_out[0][6][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][6][10] = (sum_out[1][6][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][6][10] = (sum_out[2][6][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][6][10] = (sum_out[3][6][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][6][10] = (sum_out[4][6][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][6][10] = (sum_out[5][6][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][6][10] = (sum_out[6][6][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][6][10] = (sum_out[7][6][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][6][10] = (sum_out[8][6][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][6][10] = (sum_out[9][6][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][6][10] = (sum_out[10][6][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][6][10] = (sum_out[11][6][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][6][10] = (sum_out[12][6][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][6][10] = (sum_out[13][6][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][6][10] = (sum_out[14][6][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][6][10] = (sum_out[15][6][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][6][10] = (sum_out[16][6][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][6][10] = (sum_out[17][6][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][6][10] = (sum_out[18][6][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][6][10] = (sum_out[19][6][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][6][11] = (sum_out[0][6][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][6][11] = (sum_out[1][6][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][6][11] = (sum_out[2][6][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][6][11] = (sum_out[3][6][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][6][11] = (sum_out[4][6][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][6][11] = (sum_out[5][6][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][6][11] = (sum_out[6][6][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][6][11] = (sum_out[7][6][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][6][11] = (sum_out[8][6][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][6][11] = (sum_out[9][6][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][6][11] = (sum_out[10][6][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][6][11] = (sum_out[11][6][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][6][11] = (sum_out[12][6][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][6][11] = (sum_out[13][6][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][6][11] = (sum_out[14][6][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][6][11] = (sum_out[15][6][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][6][11] = (sum_out[16][6][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][6][11] = (sum_out[17][6][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][6][11] = (sum_out[18][6][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][6][11] = (sum_out[19][6][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][6][12] = (sum_out[0][6][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][6][12] = (sum_out[1][6][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][6][12] = (sum_out[2][6][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][6][12] = (sum_out[3][6][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][6][12] = (sum_out[4][6][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][6][12] = (sum_out[5][6][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][6][12] = (sum_out[6][6][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][6][12] = (sum_out[7][6][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][6][12] = (sum_out[8][6][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][6][12] = (sum_out[9][6][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][6][12] = (sum_out[10][6][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][6][12] = (sum_out[11][6][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][6][12] = (sum_out[12][6][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][6][12] = (sum_out[13][6][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][6][12] = (sum_out[14][6][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][6][12] = (sum_out[15][6][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][6][12] = (sum_out[16][6][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][6][12] = (sum_out[17][6][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][6][12] = (sum_out[18][6][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][6][12] = (sum_out[19][6][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][6][13] = (sum_out[0][6][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][6][13] = (sum_out[1][6][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][6][13] = (sum_out[2][6][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][6][13] = (sum_out[3][6][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][6][13] = (sum_out[4][6][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][6][13] = (sum_out[5][6][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][6][13] = (sum_out[6][6][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][6][13] = (sum_out[7][6][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][6][13] = (sum_out[8][6][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][6][13] = (sum_out[9][6][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][6][13] = (sum_out[10][6][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][6][13] = (sum_out[11][6][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][6][13] = (sum_out[12][6][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][6][13] = (sum_out[13][6][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][6][13] = (sum_out[14][6][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][6][13] = (sum_out[15][6][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][6][13] = (sum_out[16][6][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][6][13] = (sum_out[17][6][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][6][13] = (sum_out[18][6][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][6][13] = (sum_out[19][6][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][6][14] = (sum_out[0][6][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][6][14] = (sum_out[1][6][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][6][14] = (sum_out[2][6][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][6][14] = (sum_out[3][6][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][6][14] = (sum_out[4][6][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][6][14] = (sum_out[5][6][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][6][14] = (sum_out[6][6][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][6][14] = (sum_out[7][6][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][6][14] = (sum_out[8][6][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][6][14] = (sum_out[9][6][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][6][14] = (sum_out[10][6][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][6][14] = (sum_out[11][6][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][6][14] = (sum_out[12][6][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][6][14] = (sum_out[13][6][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][6][14] = (sum_out[14][6][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][6][14] = (sum_out[15][6][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][6][14] = (sum_out[16][6][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][6][14] = (sum_out[17][6][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][6][14] = (sum_out[18][6][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][6][14] = (sum_out[19][6][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][6][15] = (sum_out[0][6][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][6][15] = (sum_out[1][6][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][6][15] = (sum_out[2][6][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][6][15] = (sum_out[3][6][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][6][15] = (sum_out[4][6][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][6][15] = (sum_out[5][6][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][6][15] = (sum_out[6][6][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][6][15] = (sum_out[7][6][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][6][15] = (sum_out[8][6][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][6][15] = (sum_out[9][6][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][6][15] = (sum_out[10][6][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][6][15] = (sum_out[11][6][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][6][15] = (sum_out[12][6][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][6][15] = (sum_out[13][6][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][6][15] = (sum_out[14][6][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][6][15] = (sum_out[15][6][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][6][15] = (sum_out[16][6][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][6][15] = (sum_out[17][6][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][6][15] = (sum_out[18][6][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][6][15] = (sum_out[19][6][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][6][16] = (sum_out[0][6][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][6][16] = (sum_out[1][6][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][6][16] = (sum_out[2][6][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][6][16] = (sum_out[3][6][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][6][16] = (sum_out[4][6][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][6][16] = (sum_out[5][6][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][6][16] = (sum_out[6][6][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][6][16] = (sum_out[7][6][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][6][16] = (sum_out[8][6][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][6][16] = (sum_out[9][6][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][6][16] = (sum_out[10][6][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][6][16] = (sum_out[11][6][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][6][16] = (sum_out[12][6][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][6][16] = (sum_out[13][6][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][6][16] = (sum_out[14][6][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][6][16] = (sum_out[15][6][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][6][16] = (sum_out[16][6][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][6][16] = (sum_out[17][6][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][6][16] = (sum_out[18][6][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][6][16] = (sum_out[19][6][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][6][17] = (sum_out[0][6][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][6][17] = (sum_out[1][6][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][6][17] = (sum_out[2][6][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][6][17] = (sum_out[3][6][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][6][17] = (sum_out[4][6][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][6][17] = (sum_out[5][6][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][6][17] = (sum_out[6][6][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][6][17] = (sum_out[7][6][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][6][17] = (sum_out[8][6][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][6][17] = (sum_out[9][6][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][6][17] = (sum_out[10][6][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][6][17] = (sum_out[11][6][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][6][17] = (sum_out[12][6][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][6][17] = (sum_out[13][6][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][6][17] = (sum_out[14][6][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][6][17] = (sum_out[15][6][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][6][17] = (sum_out[16][6][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][6][17] = (sum_out[17][6][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][6][17] = (sum_out[18][6][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][6][17] = (sum_out[19][6][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][6][18] = (sum_out[0][6][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][6][18] = (sum_out[1][6][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][6][18] = (sum_out[2][6][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][6][18] = (sum_out[3][6][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][6][18] = (sum_out[4][6][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][6][18] = (sum_out[5][6][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][6][18] = (sum_out[6][6][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][6][18] = (sum_out[7][6][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][6][18] = (sum_out[8][6][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][6][18] = (sum_out[9][6][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][6][18] = (sum_out[10][6][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][6][18] = (sum_out[11][6][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][6][18] = (sum_out[12][6][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][6][18] = (sum_out[13][6][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][6][18] = (sum_out[14][6][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][6][18] = (sum_out[15][6][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][6][18] = (sum_out[16][6][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][6][18] = (sum_out[17][6][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][6][18] = (sum_out[18][6][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][6][18] = (sum_out[19][6][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][6][19] = (sum_out[0][6][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][6][19] = (sum_out[1][6][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][6][19] = (sum_out[2][6][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][6][19] = (sum_out[3][6][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][6][19] = (sum_out[4][6][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][6][19] = (sum_out[5][6][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][6][19] = (sum_out[6][6][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][6][19] = (sum_out[7][6][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][6][19] = (sum_out[8][6][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][6][19] = (sum_out[9][6][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][6][19] = (sum_out[10][6][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][6][19] = (sum_out[11][6][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][6][19] = (sum_out[12][6][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][6][19] = (sum_out[13][6][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][6][19] = (sum_out[14][6][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][6][19] = (sum_out[15][6][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][6][19] = (sum_out[16][6][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][6][19] = (sum_out[17][6][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][6][19] = (sum_out[18][6][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][6][19] = (sum_out[19][6][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][6][20] = (sum_out[0][6][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][6][20] = (sum_out[1][6][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][6][20] = (sum_out[2][6][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][6][20] = (sum_out[3][6][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][6][20] = (sum_out[4][6][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][6][20] = (sum_out[5][6][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][6][20] = (sum_out[6][6][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][6][20] = (sum_out[7][6][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][6][20] = (sum_out[8][6][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][6][20] = (sum_out[9][6][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][6][20] = (sum_out[10][6][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][6][20] = (sum_out[11][6][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][6][20] = (sum_out[12][6][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][6][20] = (sum_out[13][6][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][6][20] = (sum_out[14][6][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][6][20] = (sum_out[15][6][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][6][20] = (sum_out[16][6][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][6][20] = (sum_out[17][6][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][6][20] = (sum_out[18][6][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][6][20] = (sum_out[19][6][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][6][21] = (sum_out[0][6][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][6][21] = (sum_out[1][6][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][6][21] = (sum_out[2][6][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][6][21] = (sum_out[3][6][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][6][21] = (sum_out[4][6][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][6][21] = (sum_out[5][6][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][6][21] = (sum_out[6][6][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][6][21] = (sum_out[7][6][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][6][21] = (sum_out[8][6][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][6][21] = (sum_out[9][6][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][6][21] = (sum_out[10][6][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][6][21] = (sum_out[11][6][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][6][21] = (sum_out[12][6][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][6][21] = (sum_out[13][6][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][6][21] = (sum_out[14][6][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][6][21] = (sum_out[15][6][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][6][21] = (sum_out[16][6][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][6][21] = (sum_out[17][6][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][6][21] = (sum_out[18][6][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][6][21] = (sum_out[19][6][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][6][22] = (sum_out[0][6][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][6][22] = (sum_out[1][6][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][6][22] = (sum_out[2][6][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][6][22] = (sum_out[3][6][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][6][22] = (sum_out[4][6][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][6][22] = (sum_out[5][6][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][6][22] = (sum_out[6][6][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][6][22] = (sum_out[7][6][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][6][22] = (sum_out[8][6][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][6][22] = (sum_out[9][6][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][6][22] = (sum_out[10][6][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][6][22] = (sum_out[11][6][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][6][22] = (sum_out[12][6][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][6][22] = (sum_out[13][6][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][6][22] = (sum_out[14][6][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][6][22] = (sum_out[15][6][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][6][22] = (sum_out[16][6][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][6][22] = (sum_out[17][6][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][6][22] = (sum_out[18][6][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][6][22] = (sum_out[19][6][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][6][23] = (sum_out[0][6][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][6][23] = (sum_out[1][6][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][6][23] = (sum_out[2][6][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][6][23] = (sum_out[3][6][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][6][23] = (sum_out[4][6][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][6][23] = (sum_out[5][6][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][6][23] = (sum_out[6][6][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][6][23] = (sum_out[7][6][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][6][23] = (sum_out[8][6][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][6][23] = (sum_out[9][6][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][6][23] = (sum_out[10][6][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][6][23] = (sum_out[11][6][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][6][23] = (sum_out[12][6][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][6][23] = (sum_out[13][6][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][6][23] = (sum_out[14][6][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][6][23] = (sum_out[15][6][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][6][23] = (sum_out[16][6][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][6][23] = (sum_out[17][6][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][6][23] = (sum_out[18][6][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][6][23] = (sum_out[19][6][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][7][0] = (sum_out[0][7][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][7][0] = (sum_out[1][7][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][7][0] = (sum_out[2][7][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][7][0] = (sum_out[3][7][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][7][0] = (sum_out[4][7][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][7][0] = (sum_out[5][7][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][7][0] = (sum_out[6][7][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][7][0] = (sum_out[7][7][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][7][0] = (sum_out[8][7][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][7][0] = (sum_out[9][7][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][7][0] = (sum_out[10][7][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][7][0] = (sum_out[11][7][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][7][0] = (sum_out[12][7][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][7][0] = (sum_out[13][7][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][7][0] = (sum_out[14][7][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][7][0] = (sum_out[15][7][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][7][0] = (sum_out[16][7][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][7][0] = (sum_out[17][7][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][7][0] = (sum_out[18][7][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][7][0] = (sum_out[19][7][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][7][1] = (sum_out[0][7][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][7][1] = (sum_out[1][7][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][7][1] = (sum_out[2][7][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][7][1] = (sum_out[3][7][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][7][1] = (sum_out[4][7][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][7][1] = (sum_out[5][7][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][7][1] = (sum_out[6][7][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][7][1] = (sum_out[7][7][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][7][1] = (sum_out[8][7][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][7][1] = (sum_out[9][7][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][7][1] = (sum_out[10][7][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][7][1] = (sum_out[11][7][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][7][1] = (sum_out[12][7][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][7][1] = (sum_out[13][7][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][7][1] = (sum_out[14][7][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][7][1] = (sum_out[15][7][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][7][1] = (sum_out[16][7][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][7][1] = (sum_out[17][7][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][7][1] = (sum_out[18][7][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][7][1] = (sum_out[19][7][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][7][2] = (sum_out[0][7][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][7][2] = (sum_out[1][7][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][7][2] = (sum_out[2][7][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][7][2] = (sum_out[3][7][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][7][2] = (sum_out[4][7][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][7][2] = (sum_out[5][7][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][7][2] = (sum_out[6][7][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][7][2] = (sum_out[7][7][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][7][2] = (sum_out[8][7][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][7][2] = (sum_out[9][7][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][7][2] = (sum_out[10][7][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][7][2] = (sum_out[11][7][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][7][2] = (sum_out[12][7][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][7][2] = (sum_out[13][7][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][7][2] = (sum_out[14][7][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][7][2] = (sum_out[15][7][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][7][2] = (sum_out[16][7][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][7][2] = (sum_out[17][7][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][7][2] = (sum_out[18][7][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][7][2] = (sum_out[19][7][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][7][3] = (sum_out[0][7][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][7][3] = (sum_out[1][7][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][7][3] = (sum_out[2][7][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][7][3] = (sum_out[3][7][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][7][3] = (sum_out[4][7][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][7][3] = (sum_out[5][7][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][7][3] = (sum_out[6][7][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][7][3] = (sum_out[7][7][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][7][3] = (sum_out[8][7][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][7][3] = (sum_out[9][7][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][7][3] = (sum_out[10][7][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][7][3] = (sum_out[11][7][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][7][3] = (sum_out[12][7][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][7][3] = (sum_out[13][7][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][7][3] = (sum_out[14][7][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][7][3] = (sum_out[15][7][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][7][3] = (sum_out[16][7][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][7][3] = (sum_out[17][7][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][7][3] = (sum_out[18][7][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][7][3] = (sum_out[19][7][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][7][4] = (sum_out[0][7][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][7][4] = (sum_out[1][7][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][7][4] = (sum_out[2][7][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][7][4] = (sum_out[3][7][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][7][4] = (sum_out[4][7][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][7][4] = (sum_out[5][7][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][7][4] = (sum_out[6][7][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][7][4] = (sum_out[7][7][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][7][4] = (sum_out[8][7][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][7][4] = (sum_out[9][7][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][7][4] = (sum_out[10][7][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][7][4] = (sum_out[11][7][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][7][4] = (sum_out[12][7][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][7][4] = (sum_out[13][7][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][7][4] = (sum_out[14][7][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][7][4] = (sum_out[15][7][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][7][4] = (sum_out[16][7][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][7][4] = (sum_out[17][7][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][7][4] = (sum_out[18][7][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][7][4] = (sum_out[19][7][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][7][5] = (sum_out[0][7][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][7][5] = (sum_out[1][7][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][7][5] = (sum_out[2][7][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][7][5] = (sum_out[3][7][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][7][5] = (sum_out[4][7][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][7][5] = (sum_out[5][7][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][7][5] = (sum_out[6][7][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][7][5] = (sum_out[7][7][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][7][5] = (sum_out[8][7][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][7][5] = (sum_out[9][7][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][7][5] = (sum_out[10][7][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][7][5] = (sum_out[11][7][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][7][5] = (sum_out[12][7][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][7][5] = (sum_out[13][7][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][7][5] = (sum_out[14][7][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][7][5] = (sum_out[15][7][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][7][5] = (sum_out[16][7][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][7][5] = (sum_out[17][7][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][7][5] = (sum_out[18][7][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][7][5] = (sum_out[19][7][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][7][6] = (sum_out[0][7][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][7][6] = (sum_out[1][7][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][7][6] = (sum_out[2][7][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][7][6] = (sum_out[3][7][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][7][6] = (sum_out[4][7][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][7][6] = (sum_out[5][7][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][7][6] = (sum_out[6][7][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][7][6] = (sum_out[7][7][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][7][6] = (sum_out[8][7][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][7][6] = (sum_out[9][7][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][7][6] = (sum_out[10][7][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][7][6] = (sum_out[11][7][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][7][6] = (sum_out[12][7][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][7][6] = (sum_out[13][7][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][7][6] = (sum_out[14][7][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][7][6] = (sum_out[15][7][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][7][6] = (sum_out[16][7][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][7][6] = (sum_out[17][7][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][7][6] = (sum_out[18][7][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][7][6] = (sum_out[19][7][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][7][7] = (sum_out[0][7][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][7][7] = (sum_out[1][7][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][7][7] = (sum_out[2][7][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][7][7] = (sum_out[3][7][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][7][7] = (sum_out[4][7][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][7][7] = (sum_out[5][7][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][7][7] = (sum_out[6][7][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][7][7] = (sum_out[7][7][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][7][7] = (sum_out[8][7][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][7][7] = (sum_out[9][7][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][7][7] = (sum_out[10][7][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][7][7] = (sum_out[11][7][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][7][7] = (sum_out[12][7][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][7][7] = (sum_out[13][7][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][7][7] = (sum_out[14][7][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][7][7] = (sum_out[15][7][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][7][7] = (sum_out[16][7][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][7][7] = (sum_out[17][7][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][7][7] = (sum_out[18][7][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][7][7] = (sum_out[19][7][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][7][8] = (sum_out[0][7][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][7][8] = (sum_out[1][7][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][7][8] = (sum_out[2][7][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][7][8] = (sum_out[3][7][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][7][8] = (sum_out[4][7][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][7][8] = (sum_out[5][7][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][7][8] = (sum_out[6][7][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][7][8] = (sum_out[7][7][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][7][8] = (sum_out[8][7][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][7][8] = (sum_out[9][7][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][7][8] = (sum_out[10][7][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][7][8] = (sum_out[11][7][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][7][8] = (sum_out[12][7][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][7][8] = (sum_out[13][7][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][7][8] = (sum_out[14][7][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][7][8] = (sum_out[15][7][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][7][8] = (sum_out[16][7][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][7][8] = (sum_out[17][7][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][7][8] = (sum_out[18][7][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][7][8] = (sum_out[19][7][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][7][9] = (sum_out[0][7][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][7][9] = (sum_out[1][7][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][7][9] = (sum_out[2][7][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][7][9] = (sum_out[3][7][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][7][9] = (sum_out[4][7][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][7][9] = (sum_out[5][7][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][7][9] = (sum_out[6][7][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][7][9] = (sum_out[7][7][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][7][9] = (sum_out[8][7][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][7][9] = (sum_out[9][7][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][7][9] = (sum_out[10][7][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][7][9] = (sum_out[11][7][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][7][9] = (sum_out[12][7][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][7][9] = (sum_out[13][7][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][7][9] = (sum_out[14][7][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][7][9] = (sum_out[15][7][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][7][9] = (sum_out[16][7][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][7][9] = (sum_out[17][7][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][7][9] = (sum_out[18][7][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][7][9] = (sum_out[19][7][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][7][10] = (sum_out[0][7][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][7][10] = (sum_out[1][7][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][7][10] = (sum_out[2][7][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][7][10] = (sum_out[3][7][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][7][10] = (sum_out[4][7][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][7][10] = (sum_out[5][7][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][7][10] = (sum_out[6][7][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][7][10] = (sum_out[7][7][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][7][10] = (sum_out[8][7][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][7][10] = (sum_out[9][7][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][7][10] = (sum_out[10][7][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][7][10] = (sum_out[11][7][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][7][10] = (sum_out[12][7][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][7][10] = (sum_out[13][7][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][7][10] = (sum_out[14][7][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][7][10] = (sum_out[15][7][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][7][10] = (sum_out[16][7][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][7][10] = (sum_out[17][7][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][7][10] = (sum_out[18][7][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][7][10] = (sum_out[19][7][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][7][11] = (sum_out[0][7][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][7][11] = (sum_out[1][7][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][7][11] = (sum_out[2][7][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][7][11] = (sum_out[3][7][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][7][11] = (sum_out[4][7][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][7][11] = (sum_out[5][7][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][7][11] = (sum_out[6][7][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][7][11] = (sum_out[7][7][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][7][11] = (sum_out[8][7][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][7][11] = (sum_out[9][7][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][7][11] = (sum_out[10][7][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][7][11] = (sum_out[11][7][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][7][11] = (sum_out[12][7][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][7][11] = (sum_out[13][7][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][7][11] = (sum_out[14][7][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][7][11] = (sum_out[15][7][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][7][11] = (sum_out[16][7][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][7][11] = (sum_out[17][7][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][7][11] = (sum_out[18][7][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][7][11] = (sum_out[19][7][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][7][12] = (sum_out[0][7][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][7][12] = (sum_out[1][7][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][7][12] = (sum_out[2][7][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][7][12] = (sum_out[3][7][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][7][12] = (sum_out[4][7][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][7][12] = (sum_out[5][7][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][7][12] = (sum_out[6][7][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][7][12] = (sum_out[7][7][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][7][12] = (sum_out[8][7][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][7][12] = (sum_out[9][7][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][7][12] = (sum_out[10][7][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][7][12] = (sum_out[11][7][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][7][12] = (sum_out[12][7][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][7][12] = (sum_out[13][7][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][7][12] = (sum_out[14][7][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][7][12] = (sum_out[15][7][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][7][12] = (sum_out[16][7][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][7][12] = (sum_out[17][7][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][7][12] = (sum_out[18][7][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][7][12] = (sum_out[19][7][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][7][13] = (sum_out[0][7][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][7][13] = (sum_out[1][7][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][7][13] = (sum_out[2][7][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][7][13] = (sum_out[3][7][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][7][13] = (sum_out[4][7][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][7][13] = (sum_out[5][7][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][7][13] = (sum_out[6][7][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][7][13] = (sum_out[7][7][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][7][13] = (sum_out[8][7][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][7][13] = (sum_out[9][7][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][7][13] = (sum_out[10][7][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][7][13] = (sum_out[11][7][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][7][13] = (sum_out[12][7][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][7][13] = (sum_out[13][7][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][7][13] = (sum_out[14][7][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][7][13] = (sum_out[15][7][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][7][13] = (sum_out[16][7][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][7][13] = (sum_out[17][7][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][7][13] = (sum_out[18][7][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][7][13] = (sum_out[19][7][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][7][14] = (sum_out[0][7][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][7][14] = (sum_out[1][7][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][7][14] = (sum_out[2][7][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][7][14] = (sum_out[3][7][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][7][14] = (sum_out[4][7][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][7][14] = (sum_out[5][7][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][7][14] = (sum_out[6][7][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][7][14] = (sum_out[7][7][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][7][14] = (sum_out[8][7][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][7][14] = (sum_out[9][7][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][7][14] = (sum_out[10][7][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][7][14] = (sum_out[11][7][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][7][14] = (sum_out[12][7][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][7][14] = (sum_out[13][7][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][7][14] = (sum_out[14][7][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][7][14] = (sum_out[15][7][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][7][14] = (sum_out[16][7][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][7][14] = (sum_out[17][7][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][7][14] = (sum_out[18][7][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][7][14] = (sum_out[19][7][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][7][15] = (sum_out[0][7][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][7][15] = (sum_out[1][7][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][7][15] = (sum_out[2][7][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][7][15] = (sum_out[3][7][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][7][15] = (sum_out[4][7][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][7][15] = (sum_out[5][7][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][7][15] = (sum_out[6][7][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][7][15] = (sum_out[7][7][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][7][15] = (sum_out[8][7][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][7][15] = (sum_out[9][7][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][7][15] = (sum_out[10][7][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][7][15] = (sum_out[11][7][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][7][15] = (sum_out[12][7][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][7][15] = (sum_out[13][7][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][7][15] = (sum_out[14][7][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][7][15] = (sum_out[15][7][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][7][15] = (sum_out[16][7][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][7][15] = (sum_out[17][7][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][7][15] = (sum_out[18][7][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][7][15] = (sum_out[19][7][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][7][16] = (sum_out[0][7][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][7][16] = (sum_out[1][7][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][7][16] = (sum_out[2][7][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][7][16] = (sum_out[3][7][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][7][16] = (sum_out[4][7][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][7][16] = (sum_out[5][7][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][7][16] = (sum_out[6][7][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][7][16] = (sum_out[7][7][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][7][16] = (sum_out[8][7][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][7][16] = (sum_out[9][7][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][7][16] = (sum_out[10][7][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][7][16] = (sum_out[11][7][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][7][16] = (sum_out[12][7][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][7][16] = (sum_out[13][7][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][7][16] = (sum_out[14][7][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][7][16] = (sum_out[15][7][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][7][16] = (sum_out[16][7][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][7][16] = (sum_out[17][7][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][7][16] = (sum_out[18][7][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][7][16] = (sum_out[19][7][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][7][17] = (sum_out[0][7][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][7][17] = (sum_out[1][7][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][7][17] = (sum_out[2][7][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][7][17] = (sum_out[3][7][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][7][17] = (sum_out[4][7][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][7][17] = (sum_out[5][7][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][7][17] = (sum_out[6][7][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][7][17] = (sum_out[7][7][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][7][17] = (sum_out[8][7][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][7][17] = (sum_out[9][7][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][7][17] = (sum_out[10][7][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][7][17] = (sum_out[11][7][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][7][17] = (sum_out[12][7][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][7][17] = (sum_out[13][7][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][7][17] = (sum_out[14][7][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][7][17] = (sum_out[15][7][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][7][17] = (sum_out[16][7][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][7][17] = (sum_out[17][7][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][7][17] = (sum_out[18][7][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][7][17] = (sum_out[19][7][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][7][18] = (sum_out[0][7][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][7][18] = (sum_out[1][7][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][7][18] = (sum_out[2][7][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][7][18] = (sum_out[3][7][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][7][18] = (sum_out[4][7][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][7][18] = (sum_out[5][7][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][7][18] = (sum_out[6][7][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][7][18] = (sum_out[7][7][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][7][18] = (sum_out[8][7][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][7][18] = (sum_out[9][7][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][7][18] = (sum_out[10][7][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][7][18] = (sum_out[11][7][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][7][18] = (sum_out[12][7][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][7][18] = (sum_out[13][7][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][7][18] = (sum_out[14][7][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][7][18] = (sum_out[15][7][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][7][18] = (sum_out[16][7][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][7][18] = (sum_out[17][7][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][7][18] = (sum_out[18][7][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][7][18] = (sum_out[19][7][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][7][19] = (sum_out[0][7][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][7][19] = (sum_out[1][7][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][7][19] = (sum_out[2][7][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][7][19] = (sum_out[3][7][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][7][19] = (sum_out[4][7][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][7][19] = (sum_out[5][7][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][7][19] = (sum_out[6][7][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][7][19] = (sum_out[7][7][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][7][19] = (sum_out[8][7][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][7][19] = (sum_out[9][7][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][7][19] = (sum_out[10][7][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][7][19] = (sum_out[11][7][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][7][19] = (sum_out[12][7][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][7][19] = (sum_out[13][7][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][7][19] = (sum_out[14][7][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][7][19] = (sum_out[15][7][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][7][19] = (sum_out[16][7][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][7][19] = (sum_out[17][7][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][7][19] = (sum_out[18][7][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][7][19] = (sum_out[19][7][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][7][20] = (sum_out[0][7][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][7][20] = (sum_out[1][7][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][7][20] = (sum_out[2][7][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][7][20] = (sum_out[3][7][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][7][20] = (sum_out[4][7][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][7][20] = (sum_out[5][7][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][7][20] = (sum_out[6][7][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][7][20] = (sum_out[7][7][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][7][20] = (sum_out[8][7][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][7][20] = (sum_out[9][7][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][7][20] = (sum_out[10][7][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][7][20] = (sum_out[11][7][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][7][20] = (sum_out[12][7][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][7][20] = (sum_out[13][7][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][7][20] = (sum_out[14][7][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][7][20] = (sum_out[15][7][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][7][20] = (sum_out[16][7][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][7][20] = (sum_out[17][7][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][7][20] = (sum_out[18][7][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][7][20] = (sum_out[19][7][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][7][21] = (sum_out[0][7][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][7][21] = (sum_out[1][7][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][7][21] = (sum_out[2][7][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][7][21] = (sum_out[3][7][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][7][21] = (sum_out[4][7][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][7][21] = (sum_out[5][7][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][7][21] = (sum_out[6][7][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][7][21] = (sum_out[7][7][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][7][21] = (sum_out[8][7][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][7][21] = (sum_out[9][7][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][7][21] = (sum_out[10][7][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][7][21] = (sum_out[11][7][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][7][21] = (sum_out[12][7][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][7][21] = (sum_out[13][7][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][7][21] = (sum_out[14][7][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][7][21] = (sum_out[15][7][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][7][21] = (sum_out[16][7][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][7][21] = (sum_out[17][7][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][7][21] = (sum_out[18][7][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][7][21] = (sum_out[19][7][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][7][22] = (sum_out[0][7][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][7][22] = (sum_out[1][7][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][7][22] = (sum_out[2][7][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][7][22] = (sum_out[3][7][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][7][22] = (sum_out[4][7][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][7][22] = (sum_out[5][7][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][7][22] = (sum_out[6][7][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][7][22] = (sum_out[7][7][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][7][22] = (sum_out[8][7][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][7][22] = (sum_out[9][7][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][7][22] = (sum_out[10][7][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][7][22] = (sum_out[11][7][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][7][22] = (sum_out[12][7][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][7][22] = (sum_out[13][7][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][7][22] = (sum_out[14][7][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][7][22] = (sum_out[15][7][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][7][22] = (sum_out[16][7][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][7][22] = (sum_out[17][7][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][7][22] = (sum_out[18][7][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][7][22] = (sum_out[19][7][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][7][23] = (sum_out[0][7][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][7][23] = (sum_out[1][7][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][7][23] = (sum_out[2][7][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][7][23] = (sum_out[3][7][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][7][23] = (sum_out[4][7][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][7][23] = (sum_out[5][7][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][7][23] = (sum_out[6][7][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][7][23] = (sum_out[7][7][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][7][23] = (sum_out[8][7][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][7][23] = (sum_out[9][7][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][7][23] = (sum_out[10][7][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][7][23] = (sum_out[11][7][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][7][23] = (sum_out[12][7][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][7][23] = (sum_out[13][7][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][7][23] = (sum_out[14][7][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][7][23] = (sum_out[15][7][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][7][23] = (sum_out[16][7][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][7][23] = (sum_out[17][7][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][7][23] = (sum_out[18][7][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][7][23] = (sum_out[19][7][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][8][0] = (sum_out[0][8][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][8][0] = (sum_out[1][8][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][8][0] = (sum_out[2][8][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][8][0] = (sum_out[3][8][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][8][0] = (sum_out[4][8][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][8][0] = (sum_out[5][8][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][8][0] = (sum_out[6][8][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][8][0] = (sum_out[7][8][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][8][0] = (sum_out[8][8][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][8][0] = (sum_out[9][8][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][8][0] = (sum_out[10][8][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][8][0] = (sum_out[11][8][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][8][0] = (sum_out[12][8][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][8][0] = (sum_out[13][8][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][8][0] = (sum_out[14][8][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][8][0] = (sum_out[15][8][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][8][0] = (sum_out[16][8][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][8][0] = (sum_out[17][8][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][8][0] = (sum_out[18][8][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][8][0] = (sum_out[19][8][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][8][1] = (sum_out[0][8][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][8][1] = (sum_out[1][8][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][8][1] = (sum_out[2][8][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][8][1] = (sum_out[3][8][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][8][1] = (sum_out[4][8][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][8][1] = (sum_out[5][8][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][8][1] = (sum_out[6][8][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][8][1] = (sum_out[7][8][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][8][1] = (sum_out[8][8][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][8][1] = (sum_out[9][8][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][8][1] = (sum_out[10][8][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][8][1] = (sum_out[11][8][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][8][1] = (sum_out[12][8][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][8][1] = (sum_out[13][8][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][8][1] = (sum_out[14][8][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][8][1] = (sum_out[15][8][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][8][1] = (sum_out[16][8][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][8][1] = (sum_out[17][8][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][8][1] = (sum_out[18][8][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][8][1] = (sum_out[19][8][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][8][2] = (sum_out[0][8][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][8][2] = (sum_out[1][8][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][8][2] = (sum_out[2][8][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][8][2] = (sum_out[3][8][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][8][2] = (sum_out[4][8][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][8][2] = (sum_out[5][8][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][8][2] = (sum_out[6][8][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][8][2] = (sum_out[7][8][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][8][2] = (sum_out[8][8][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][8][2] = (sum_out[9][8][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][8][2] = (sum_out[10][8][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][8][2] = (sum_out[11][8][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][8][2] = (sum_out[12][8][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][8][2] = (sum_out[13][8][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][8][2] = (sum_out[14][8][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][8][2] = (sum_out[15][8][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][8][2] = (sum_out[16][8][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][8][2] = (sum_out[17][8][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][8][2] = (sum_out[18][8][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][8][2] = (sum_out[19][8][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][8][3] = (sum_out[0][8][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][8][3] = (sum_out[1][8][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][8][3] = (sum_out[2][8][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][8][3] = (sum_out[3][8][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][8][3] = (sum_out[4][8][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][8][3] = (sum_out[5][8][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][8][3] = (sum_out[6][8][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][8][3] = (sum_out[7][8][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][8][3] = (sum_out[8][8][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][8][3] = (sum_out[9][8][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][8][3] = (sum_out[10][8][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][8][3] = (sum_out[11][8][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][8][3] = (sum_out[12][8][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][8][3] = (sum_out[13][8][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][8][3] = (sum_out[14][8][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][8][3] = (sum_out[15][8][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][8][3] = (sum_out[16][8][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][8][3] = (sum_out[17][8][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][8][3] = (sum_out[18][8][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][8][3] = (sum_out[19][8][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][8][4] = (sum_out[0][8][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][8][4] = (sum_out[1][8][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][8][4] = (sum_out[2][8][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][8][4] = (sum_out[3][8][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][8][4] = (sum_out[4][8][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][8][4] = (sum_out[5][8][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][8][4] = (sum_out[6][8][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][8][4] = (sum_out[7][8][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][8][4] = (sum_out[8][8][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][8][4] = (sum_out[9][8][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][8][4] = (sum_out[10][8][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][8][4] = (sum_out[11][8][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][8][4] = (sum_out[12][8][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][8][4] = (sum_out[13][8][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][8][4] = (sum_out[14][8][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][8][4] = (sum_out[15][8][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][8][4] = (sum_out[16][8][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][8][4] = (sum_out[17][8][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][8][4] = (sum_out[18][8][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][8][4] = (sum_out[19][8][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][8][5] = (sum_out[0][8][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][8][5] = (sum_out[1][8][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][8][5] = (sum_out[2][8][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][8][5] = (sum_out[3][8][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][8][5] = (sum_out[4][8][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][8][5] = (sum_out[5][8][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][8][5] = (sum_out[6][8][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][8][5] = (sum_out[7][8][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][8][5] = (sum_out[8][8][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][8][5] = (sum_out[9][8][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][8][5] = (sum_out[10][8][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][8][5] = (sum_out[11][8][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][8][5] = (sum_out[12][8][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][8][5] = (sum_out[13][8][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][8][5] = (sum_out[14][8][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][8][5] = (sum_out[15][8][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][8][5] = (sum_out[16][8][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][8][5] = (sum_out[17][8][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][8][5] = (sum_out[18][8][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][8][5] = (sum_out[19][8][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][8][6] = (sum_out[0][8][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][8][6] = (sum_out[1][8][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][8][6] = (sum_out[2][8][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][8][6] = (sum_out[3][8][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][8][6] = (sum_out[4][8][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][8][6] = (sum_out[5][8][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][8][6] = (sum_out[6][8][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][8][6] = (sum_out[7][8][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][8][6] = (sum_out[8][8][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][8][6] = (sum_out[9][8][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][8][6] = (sum_out[10][8][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][8][6] = (sum_out[11][8][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][8][6] = (sum_out[12][8][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][8][6] = (sum_out[13][8][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][8][6] = (sum_out[14][8][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][8][6] = (sum_out[15][8][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][8][6] = (sum_out[16][8][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][8][6] = (sum_out[17][8][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][8][6] = (sum_out[18][8][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][8][6] = (sum_out[19][8][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][8][7] = (sum_out[0][8][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][8][7] = (sum_out[1][8][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][8][7] = (sum_out[2][8][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][8][7] = (sum_out[3][8][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][8][7] = (sum_out[4][8][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][8][7] = (sum_out[5][8][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][8][7] = (sum_out[6][8][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][8][7] = (sum_out[7][8][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][8][7] = (sum_out[8][8][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][8][7] = (sum_out[9][8][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][8][7] = (sum_out[10][8][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][8][7] = (sum_out[11][8][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][8][7] = (sum_out[12][8][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][8][7] = (sum_out[13][8][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][8][7] = (sum_out[14][8][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][8][7] = (sum_out[15][8][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][8][7] = (sum_out[16][8][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][8][7] = (sum_out[17][8][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][8][7] = (sum_out[18][8][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][8][7] = (sum_out[19][8][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][8][8] = (sum_out[0][8][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][8][8] = (sum_out[1][8][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][8][8] = (sum_out[2][8][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][8][8] = (sum_out[3][8][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][8][8] = (sum_out[4][8][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][8][8] = (sum_out[5][8][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][8][8] = (sum_out[6][8][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][8][8] = (sum_out[7][8][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][8][8] = (sum_out[8][8][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][8][8] = (sum_out[9][8][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][8][8] = (sum_out[10][8][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][8][8] = (sum_out[11][8][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][8][8] = (sum_out[12][8][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][8][8] = (sum_out[13][8][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][8][8] = (sum_out[14][8][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][8][8] = (sum_out[15][8][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][8][8] = (sum_out[16][8][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][8][8] = (sum_out[17][8][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][8][8] = (sum_out[18][8][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][8][8] = (sum_out[19][8][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][8][9] = (sum_out[0][8][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][8][9] = (sum_out[1][8][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][8][9] = (sum_out[2][8][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][8][9] = (sum_out[3][8][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][8][9] = (sum_out[4][8][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][8][9] = (sum_out[5][8][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][8][9] = (sum_out[6][8][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][8][9] = (sum_out[7][8][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][8][9] = (sum_out[8][8][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][8][9] = (sum_out[9][8][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][8][9] = (sum_out[10][8][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][8][9] = (sum_out[11][8][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][8][9] = (sum_out[12][8][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][8][9] = (sum_out[13][8][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][8][9] = (sum_out[14][8][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][8][9] = (sum_out[15][8][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][8][9] = (sum_out[16][8][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][8][9] = (sum_out[17][8][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][8][9] = (sum_out[18][8][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][8][9] = (sum_out[19][8][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][8][10] = (sum_out[0][8][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][8][10] = (sum_out[1][8][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][8][10] = (sum_out[2][8][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][8][10] = (sum_out[3][8][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][8][10] = (sum_out[4][8][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][8][10] = (sum_out[5][8][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][8][10] = (sum_out[6][8][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][8][10] = (sum_out[7][8][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][8][10] = (sum_out[8][8][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][8][10] = (sum_out[9][8][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][8][10] = (sum_out[10][8][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][8][10] = (sum_out[11][8][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][8][10] = (sum_out[12][8][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][8][10] = (sum_out[13][8][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][8][10] = (sum_out[14][8][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][8][10] = (sum_out[15][8][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][8][10] = (sum_out[16][8][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][8][10] = (sum_out[17][8][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][8][10] = (sum_out[18][8][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][8][10] = (sum_out[19][8][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][8][11] = (sum_out[0][8][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][8][11] = (sum_out[1][8][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][8][11] = (sum_out[2][8][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][8][11] = (sum_out[3][8][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][8][11] = (sum_out[4][8][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][8][11] = (sum_out[5][8][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][8][11] = (sum_out[6][8][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][8][11] = (sum_out[7][8][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][8][11] = (sum_out[8][8][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][8][11] = (sum_out[9][8][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][8][11] = (sum_out[10][8][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][8][11] = (sum_out[11][8][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][8][11] = (sum_out[12][8][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][8][11] = (sum_out[13][8][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][8][11] = (sum_out[14][8][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][8][11] = (sum_out[15][8][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][8][11] = (sum_out[16][8][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][8][11] = (sum_out[17][8][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][8][11] = (sum_out[18][8][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][8][11] = (sum_out[19][8][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][8][12] = (sum_out[0][8][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][8][12] = (sum_out[1][8][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][8][12] = (sum_out[2][8][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][8][12] = (sum_out[3][8][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][8][12] = (sum_out[4][8][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][8][12] = (sum_out[5][8][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][8][12] = (sum_out[6][8][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][8][12] = (sum_out[7][8][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][8][12] = (sum_out[8][8][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][8][12] = (sum_out[9][8][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][8][12] = (sum_out[10][8][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][8][12] = (sum_out[11][8][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][8][12] = (sum_out[12][8][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][8][12] = (sum_out[13][8][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][8][12] = (sum_out[14][8][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][8][12] = (sum_out[15][8][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][8][12] = (sum_out[16][8][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][8][12] = (sum_out[17][8][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][8][12] = (sum_out[18][8][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][8][12] = (sum_out[19][8][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][8][13] = (sum_out[0][8][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][8][13] = (sum_out[1][8][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][8][13] = (sum_out[2][8][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][8][13] = (sum_out[3][8][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][8][13] = (sum_out[4][8][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][8][13] = (sum_out[5][8][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][8][13] = (sum_out[6][8][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][8][13] = (sum_out[7][8][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][8][13] = (sum_out[8][8][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][8][13] = (sum_out[9][8][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][8][13] = (sum_out[10][8][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][8][13] = (sum_out[11][8][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][8][13] = (sum_out[12][8][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][8][13] = (sum_out[13][8][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][8][13] = (sum_out[14][8][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][8][13] = (sum_out[15][8][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][8][13] = (sum_out[16][8][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][8][13] = (sum_out[17][8][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][8][13] = (sum_out[18][8][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][8][13] = (sum_out[19][8][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][8][14] = (sum_out[0][8][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][8][14] = (sum_out[1][8][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][8][14] = (sum_out[2][8][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][8][14] = (sum_out[3][8][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][8][14] = (sum_out[4][8][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][8][14] = (sum_out[5][8][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][8][14] = (sum_out[6][8][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][8][14] = (sum_out[7][8][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][8][14] = (sum_out[8][8][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][8][14] = (sum_out[9][8][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][8][14] = (sum_out[10][8][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][8][14] = (sum_out[11][8][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][8][14] = (sum_out[12][8][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][8][14] = (sum_out[13][8][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][8][14] = (sum_out[14][8][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][8][14] = (sum_out[15][8][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][8][14] = (sum_out[16][8][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][8][14] = (sum_out[17][8][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][8][14] = (sum_out[18][8][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][8][14] = (sum_out[19][8][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][8][15] = (sum_out[0][8][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][8][15] = (sum_out[1][8][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][8][15] = (sum_out[2][8][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][8][15] = (sum_out[3][8][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][8][15] = (sum_out[4][8][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][8][15] = (sum_out[5][8][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][8][15] = (sum_out[6][8][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][8][15] = (sum_out[7][8][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][8][15] = (sum_out[8][8][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][8][15] = (sum_out[9][8][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][8][15] = (sum_out[10][8][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][8][15] = (sum_out[11][8][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][8][15] = (sum_out[12][8][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][8][15] = (sum_out[13][8][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][8][15] = (sum_out[14][8][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][8][15] = (sum_out[15][8][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][8][15] = (sum_out[16][8][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][8][15] = (sum_out[17][8][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][8][15] = (sum_out[18][8][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][8][15] = (sum_out[19][8][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][8][16] = (sum_out[0][8][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][8][16] = (sum_out[1][8][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][8][16] = (sum_out[2][8][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][8][16] = (sum_out[3][8][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][8][16] = (sum_out[4][8][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][8][16] = (sum_out[5][8][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][8][16] = (sum_out[6][8][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][8][16] = (sum_out[7][8][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][8][16] = (sum_out[8][8][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][8][16] = (sum_out[9][8][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][8][16] = (sum_out[10][8][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][8][16] = (sum_out[11][8][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][8][16] = (sum_out[12][8][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][8][16] = (sum_out[13][8][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][8][16] = (sum_out[14][8][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][8][16] = (sum_out[15][8][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][8][16] = (sum_out[16][8][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][8][16] = (sum_out[17][8][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][8][16] = (sum_out[18][8][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][8][16] = (sum_out[19][8][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][8][17] = (sum_out[0][8][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][8][17] = (sum_out[1][8][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][8][17] = (sum_out[2][8][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][8][17] = (sum_out[3][8][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][8][17] = (sum_out[4][8][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][8][17] = (sum_out[5][8][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][8][17] = (sum_out[6][8][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][8][17] = (sum_out[7][8][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][8][17] = (sum_out[8][8][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][8][17] = (sum_out[9][8][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][8][17] = (sum_out[10][8][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][8][17] = (sum_out[11][8][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][8][17] = (sum_out[12][8][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][8][17] = (sum_out[13][8][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][8][17] = (sum_out[14][8][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][8][17] = (sum_out[15][8][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][8][17] = (sum_out[16][8][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][8][17] = (sum_out[17][8][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][8][17] = (sum_out[18][8][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][8][17] = (sum_out[19][8][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][8][18] = (sum_out[0][8][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][8][18] = (sum_out[1][8][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][8][18] = (sum_out[2][8][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][8][18] = (sum_out[3][8][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][8][18] = (sum_out[4][8][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][8][18] = (sum_out[5][8][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][8][18] = (sum_out[6][8][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][8][18] = (sum_out[7][8][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][8][18] = (sum_out[8][8][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][8][18] = (sum_out[9][8][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][8][18] = (sum_out[10][8][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][8][18] = (sum_out[11][8][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][8][18] = (sum_out[12][8][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][8][18] = (sum_out[13][8][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][8][18] = (sum_out[14][8][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][8][18] = (sum_out[15][8][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][8][18] = (sum_out[16][8][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][8][18] = (sum_out[17][8][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][8][18] = (sum_out[18][8][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][8][18] = (sum_out[19][8][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][8][19] = (sum_out[0][8][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][8][19] = (sum_out[1][8][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][8][19] = (sum_out[2][8][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][8][19] = (sum_out[3][8][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][8][19] = (sum_out[4][8][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][8][19] = (sum_out[5][8][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][8][19] = (sum_out[6][8][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][8][19] = (sum_out[7][8][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][8][19] = (sum_out[8][8][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][8][19] = (sum_out[9][8][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][8][19] = (sum_out[10][8][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][8][19] = (sum_out[11][8][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][8][19] = (sum_out[12][8][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][8][19] = (sum_out[13][8][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][8][19] = (sum_out[14][8][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][8][19] = (sum_out[15][8][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][8][19] = (sum_out[16][8][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][8][19] = (sum_out[17][8][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][8][19] = (sum_out[18][8][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][8][19] = (sum_out[19][8][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][8][20] = (sum_out[0][8][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][8][20] = (sum_out[1][8][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][8][20] = (sum_out[2][8][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][8][20] = (sum_out[3][8][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][8][20] = (sum_out[4][8][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][8][20] = (sum_out[5][8][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][8][20] = (sum_out[6][8][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][8][20] = (sum_out[7][8][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][8][20] = (sum_out[8][8][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][8][20] = (sum_out[9][8][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][8][20] = (sum_out[10][8][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][8][20] = (sum_out[11][8][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][8][20] = (sum_out[12][8][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][8][20] = (sum_out[13][8][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][8][20] = (sum_out[14][8][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][8][20] = (sum_out[15][8][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][8][20] = (sum_out[16][8][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][8][20] = (sum_out[17][8][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][8][20] = (sum_out[18][8][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][8][20] = (sum_out[19][8][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][8][21] = (sum_out[0][8][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][8][21] = (sum_out[1][8][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][8][21] = (sum_out[2][8][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][8][21] = (sum_out[3][8][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][8][21] = (sum_out[4][8][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][8][21] = (sum_out[5][8][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][8][21] = (sum_out[6][8][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][8][21] = (sum_out[7][8][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][8][21] = (sum_out[8][8][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][8][21] = (sum_out[9][8][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][8][21] = (sum_out[10][8][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][8][21] = (sum_out[11][8][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][8][21] = (sum_out[12][8][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][8][21] = (sum_out[13][8][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][8][21] = (sum_out[14][8][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][8][21] = (sum_out[15][8][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][8][21] = (sum_out[16][8][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][8][21] = (sum_out[17][8][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][8][21] = (sum_out[18][8][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][8][21] = (sum_out[19][8][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][8][22] = (sum_out[0][8][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][8][22] = (sum_out[1][8][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][8][22] = (sum_out[2][8][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][8][22] = (sum_out[3][8][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][8][22] = (sum_out[4][8][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][8][22] = (sum_out[5][8][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][8][22] = (sum_out[6][8][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][8][22] = (sum_out[7][8][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][8][22] = (sum_out[8][8][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][8][22] = (sum_out[9][8][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][8][22] = (sum_out[10][8][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][8][22] = (sum_out[11][8][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][8][22] = (sum_out[12][8][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][8][22] = (sum_out[13][8][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][8][22] = (sum_out[14][8][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][8][22] = (sum_out[15][8][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][8][22] = (sum_out[16][8][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][8][22] = (sum_out[17][8][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][8][22] = (sum_out[18][8][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][8][22] = (sum_out[19][8][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][8][23] = (sum_out[0][8][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][8][23] = (sum_out[1][8][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][8][23] = (sum_out[2][8][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][8][23] = (sum_out[3][8][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][8][23] = (sum_out[4][8][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][8][23] = (sum_out[5][8][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][8][23] = (sum_out[6][8][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][8][23] = (sum_out[7][8][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][8][23] = (sum_out[8][8][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][8][23] = (sum_out[9][8][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][8][23] = (sum_out[10][8][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][8][23] = (sum_out[11][8][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][8][23] = (sum_out[12][8][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][8][23] = (sum_out[13][8][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][8][23] = (sum_out[14][8][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][8][23] = (sum_out[15][8][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][8][23] = (sum_out[16][8][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][8][23] = (sum_out[17][8][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][8][23] = (sum_out[18][8][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][8][23] = (sum_out[19][8][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][9][0] = (sum_out[0][9][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][9][0] = (sum_out[1][9][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][9][0] = (sum_out[2][9][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][9][0] = (sum_out[3][9][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][9][0] = (sum_out[4][9][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][9][0] = (sum_out[5][9][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][9][0] = (sum_out[6][9][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][9][0] = (sum_out[7][9][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][9][0] = (sum_out[8][9][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][9][0] = (sum_out[9][9][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][9][0] = (sum_out[10][9][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][9][0] = (sum_out[11][9][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][9][0] = (sum_out[12][9][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][9][0] = (sum_out[13][9][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][9][0] = (sum_out[14][9][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][9][0] = (sum_out[15][9][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][9][0] = (sum_out[16][9][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][9][0] = (sum_out[17][9][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][9][0] = (sum_out[18][9][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][9][0] = (sum_out[19][9][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][9][1] = (sum_out[0][9][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][9][1] = (sum_out[1][9][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][9][1] = (sum_out[2][9][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][9][1] = (sum_out[3][9][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][9][1] = (sum_out[4][9][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][9][1] = (sum_out[5][9][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][9][1] = (sum_out[6][9][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][9][1] = (sum_out[7][9][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][9][1] = (sum_out[8][9][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][9][1] = (sum_out[9][9][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][9][1] = (sum_out[10][9][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][9][1] = (sum_out[11][9][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][9][1] = (sum_out[12][9][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][9][1] = (sum_out[13][9][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][9][1] = (sum_out[14][9][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][9][1] = (sum_out[15][9][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][9][1] = (sum_out[16][9][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][9][1] = (sum_out[17][9][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][9][1] = (sum_out[18][9][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][9][1] = (sum_out[19][9][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][9][2] = (sum_out[0][9][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][9][2] = (sum_out[1][9][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][9][2] = (sum_out[2][9][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][9][2] = (sum_out[3][9][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][9][2] = (sum_out[4][9][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][9][2] = (sum_out[5][9][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][9][2] = (sum_out[6][9][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][9][2] = (sum_out[7][9][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][9][2] = (sum_out[8][9][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][9][2] = (sum_out[9][9][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][9][2] = (sum_out[10][9][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][9][2] = (sum_out[11][9][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][9][2] = (sum_out[12][9][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][9][2] = (sum_out[13][9][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][9][2] = (sum_out[14][9][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][9][2] = (sum_out[15][9][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][9][2] = (sum_out[16][9][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][9][2] = (sum_out[17][9][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][9][2] = (sum_out[18][9][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][9][2] = (sum_out[19][9][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][9][3] = (sum_out[0][9][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][9][3] = (sum_out[1][9][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][9][3] = (sum_out[2][9][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][9][3] = (sum_out[3][9][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][9][3] = (sum_out[4][9][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][9][3] = (sum_out[5][9][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][9][3] = (sum_out[6][9][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][9][3] = (sum_out[7][9][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][9][3] = (sum_out[8][9][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][9][3] = (sum_out[9][9][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][9][3] = (sum_out[10][9][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][9][3] = (sum_out[11][9][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][9][3] = (sum_out[12][9][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][9][3] = (sum_out[13][9][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][9][3] = (sum_out[14][9][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][9][3] = (sum_out[15][9][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][9][3] = (sum_out[16][9][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][9][3] = (sum_out[17][9][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][9][3] = (sum_out[18][9][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][9][3] = (sum_out[19][9][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][9][4] = (sum_out[0][9][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][9][4] = (sum_out[1][9][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][9][4] = (sum_out[2][9][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][9][4] = (sum_out[3][9][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][9][4] = (sum_out[4][9][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][9][4] = (sum_out[5][9][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][9][4] = (sum_out[6][9][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][9][4] = (sum_out[7][9][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][9][4] = (sum_out[8][9][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][9][4] = (sum_out[9][9][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][9][4] = (sum_out[10][9][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][9][4] = (sum_out[11][9][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][9][4] = (sum_out[12][9][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][9][4] = (sum_out[13][9][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][9][4] = (sum_out[14][9][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][9][4] = (sum_out[15][9][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][9][4] = (sum_out[16][9][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][9][4] = (sum_out[17][9][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][9][4] = (sum_out[18][9][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][9][4] = (sum_out[19][9][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][9][5] = (sum_out[0][9][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][9][5] = (sum_out[1][9][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][9][5] = (sum_out[2][9][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][9][5] = (sum_out[3][9][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][9][5] = (sum_out[4][9][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][9][5] = (sum_out[5][9][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][9][5] = (sum_out[6][9][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][9][5] = (sum_out[7][9][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][9][5] = (sum_out[8][9][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][9][5] = (sum_out[9][9][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][9][5] = (sum_out[10][9][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][9][5] = (sum_out[11][9][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][9][5] = (sum_out[12][9][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][9][5] = (sum_out[13][9][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][9][5] = (sum_out[14][9][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][9][5] = (sum_out[15][9][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][9][5] = (sum_out[16][9][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][9][5] = (sum_out[17][9][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][9][5] = (sum_out[18][9][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][9][5] = (sum_out[19][9][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][9][6] = (sum_out[0][9][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][9][6] = (sum_out[1][9][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][9][6] = (sum_out[2][9][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][9][6] = (sum_out[3][9][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][9][6] = (sum_out[4][9][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][9][6] = (sum_out[5][9][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][9][6] = (sum_out[6][9][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][9][6] = (sum_out[7][9][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][9][6] = (sum_out[8][9][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][9][6] = (sum_out[9][9][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][9][6] = (sum_out[10][9][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][9][6] = (sum_out[11][9][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][9][6] = (sum_out[12][9][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][9][6] = (sum_out[13][9][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][9][6] = (sum_out[14][9][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][9][6] = (sum_out[15][9][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][9][6] = (sum_out[16][9][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][9][6] = (sum_out[17][9][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][9][6] = (sum_out[18][9][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][9][6] = (sum_out[19][9][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][9][7] = (sum_out[0][9][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][9][7] = (sum_out[1][9][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][9][7] = (sum_out[2][9][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][9][7] = (sum_out[3][9][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][9][7] = (sum_out[4][9][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][9][7] = (sum_out[5][9][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][9][7] = (sum_out[6][9][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][9][7] = (sum_out[7][9][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][9][7] = (sum_out[8][9][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][9][7] = (sum_out[9][9][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][9][7] = (sum_out[10][9][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][9][7] = (sum_out[11][9][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][9][7] = (sum_out[12][9][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][9][7] = (sum_out[13][9][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][9][7] = (sum_out[14][9][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][9][7] = (sum_out[15][9][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][9][7] = (sum_out[16][9][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][9][7] = (sum_out[17][9][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][9][7] = (sum_out[18][9][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][9][7] = (sum_out[19][9][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][9][8] = (sum_out[0][9][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][9][8] = (sum_out[1][9][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][9][8] = (sum_out[2][9][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][9][8] = (sum_out[3][9][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][9][8] = (sum_out[4][9][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][9][8] = (sum_out[5][9][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][9][8] = (sum_out[6][9][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][9][8] = (sum_out[7][9][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][9][8] = (sum_out[8][9][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][9][8] = (sum_out[9][9][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][9][8] = (sum_out[10][9][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][9][8] = (sum_out[11][9][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][9][8] = (sum_out[12][9][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][9][8] = (sum_out[13][9][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][9][8] = (sum_out[14][9][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][9][8] = (sum_out[15][9][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][9][8] = (sum_out[16][9][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][9][8] = (sum_out[17][9][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][9][8] = (sum_out[18][9][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][9][8] = (sum_out[19][9][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][9][9] = (sum_out[0][9][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][9][9] = (sum_out[1][9][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][9][9] = (sum_out[2][9][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][9][9] = (sum_out[3][9][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][9][9] = (sum_out[4][9][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][9][9] = (sum_out[5][9][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][9][9] = (sum_out[6][9][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][9][9] = (sum_out[7][9][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][9][9] = (sum_out[8][9][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][9][9] = (sum_out[9][9][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][9][9] = (sum_out[10][9][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][9][9] = (sum_out[11][9][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][9][9] = (sum_out[12][9][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][9][9] = (sum_out[13][9][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][9][9] = (sum_out[14][9][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][9][9] = (sum_out[15][9][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][9][9] = (sum_out[16][9][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][9][9] = (sum_out[17][9][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][9][9] = (sum_out[18][9][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][9][9] = (sum_out[19][9][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][9][10] = (sum_out[0][9][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][9][10] = (sum_out[1][9][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][9][10] = (sum_out[2][9][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][9][10] = (sum_out[3][9][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][9][10] = (sum_out[4][9][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][9][10] = (sum_out[5][9][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][9][10] = (sum_out[6][9][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][9][10] = (sum_out[7][9][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][9][10] = (sum_out[8][9][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][9][10] = (sum_out[9][9][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][9][10] = (sum_out[10][9][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][9][10] = (sum_out[11][9][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][9][10] = (sum_out[12][9][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][9][10] = (sum_out[13][9][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][9][10] = (sum_out[14][9][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][9][10] = (sum_out[15][9][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][9][10] = (sum_out[16][9][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][9][10] = (sum_out[17][9][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][9][10] = (sum_out[18][9][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][9][10] = (sum_out[19][9][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][9][11] = (sum_out[0][9][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][9][11] = (sum_out[1][9][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][9][11] = (sum_out[2][9][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][9][11] = (sum_out[3][9][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][9][11] = (sum_out[4][9][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][9][11] = (sum_out[5][9][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][9][11] = (sum_out[6][9][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][9][11] = (sum_out[7][9][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][9][11] = (sum_out[8][9][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][9][11] = (sum_out[9][9][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][9][11] = (sum_out[10][9][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][9][11] = (sum_out[11][9][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][9][11] = (sum_out[12][9][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][9][11] = (sum_out[13][9][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][9][11] = (sum_out[14][9][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][9][11] = (sum_out[15][9][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][9][11] = (sum_out[16][9][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][9][11] = (sum_out[17][9][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][9][11] = (sum_out[18][9][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][9][11] = (sum_out[19][9][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][9][12] = (sum_out[0][9][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][9][12] = (sum_out[1][9][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][9][12] = (sum_out[2][9][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][9][12] = (sum_out[3][9][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][9][12] = (sum_out[4][9][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][9][12] = (sum_out[5][9][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][9][12] = (sum_out[6][9][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][9][12] = (sum_out[7][9][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][9][12] = (sum_out[8][9][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][9][12] = (sum_out[9][9][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][9][12] = (sum_out[10][9][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][9][12] = (sum_out[11][9][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][9][12] = (sum_out[12][9][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][9][12] = (sum_out[13][9][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][9][12] = (sum_out[14][9][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][9][12] = (sum_out[15][9][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][9][12] = (sum_out[16][9][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][9][12] = (sum_out[17][9][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][9][12] = (sum_out[18][9][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][9][12] = (sum_out[19][9][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][9][13] = (sum_out[0][9][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][9][13] = (sum_out[1][9][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][9][13] = (sum_out[2][9][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][9][13] = (sum_out[3][9][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][9][13] = (sum_out[4][9][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][9][13] = (sum_out[5][9][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][9][13] = (sum_out[6][9][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][9][13] = (sum_out[7][9][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][9][13] = (sum_out[8][9][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][9][13] = (sum_out[9][9][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][9][13] = (sum_out[10][9][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][9][13] = (sum_out[11][9][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][9][13] = (sum_out[12][9][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][9][13] = (sum_out[13][9][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][9][13] = (sum_out[14][9][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][9][13] = (sum_out[15][9][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][9][13] = (sum_out[16][9][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][9][13] = (sum_out[17][9][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][9][13] = (sum_out[18][9][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][9][13] = (sum_out[19][9][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][9][14] = (sum_out[0][9][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][9][14] = (sum_out[1][9][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][9][14] = (sum_out[2][9][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][9][14] = (sum_out[3][9][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][9][14] = (sum_out[4][9][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][9][14] = (sum_out[5][9][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][9][14] = (sum_out[6][9][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][9][14] = (sum_out[7][9][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][9][14] = (sum_out[8][9][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][9][14] = (sum_out[9][9][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][9][14] = (sum_out[10][9][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][9][14] = (sum_out[11][9][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][9][14] = (sum_out[12][9][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][9][14] = (sum_out[13][9][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][9][14] = (sum_out[14][9][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][9][14] = (sum_out[15][9][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][9][14] = (sum_out[16][9][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][9][14] = (sum_out[17][9][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][9][14] = (sum_out[18][9][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][9][14] = (sum_out[19][9][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][9][15] = (sum_out[0][9][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][9][15] = (sum_out[1][9][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][9][15] = (sum_out[2][9][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][9][15] = (sum_out[3][9][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][9][15] = (sum_out[4][9][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][9][15] = (sum_out[5][9][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][9][15] = (sum_out[6][9][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][9][15] = (sum_out[7][9][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][9][15] = (sum_out[8][9][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][9][15] = (sum_out[9][9][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][9][15] = (sum_out[10][9][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][9][15] = (sum_out[11][9][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][9][15] = (sum_out[12][9][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][9][15] = (sum_out[13][9][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][9][15] = (sum_out[14][9][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][9][15] = (sum_out[15][9][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][9][15] = (sum_out[16][9][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][9][15] = (sum_out[17][9][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][9][15] = (sum_out[18][9][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][9][15] = (sum_out[19][9][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][9][16] = (sum_out[0][9][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][9][16] = (sum_out[1][9][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][9][16] = (sum_out[2][9][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][9][16] = (sum_out[3][9][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][9][16] = (sum_out[4][9][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][9][16] = (sum_out[5][9][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][9][16] = (sum_out[6][9][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][9][16] = (sum_out[7][9][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][9][16] = (sum_out[8][9][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][9][16] = (sum_out[9][9][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][9][16] = (sum_out[10][9][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][9][16] = (sum_out[11][9][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][9][16] = (sum_out[12][9][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][9][16] = (sum_out[13][9][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][9][16] = (sum_out[14][9][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][9][16] = (sum_out[15][9][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][9][16] = (sum_out[16][9][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][9][16] = (sum_out[17][9][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][9][16] = (sum_out[18][9][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][9][16] = (sum_out[19][9][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][9][17] = (sum_out[0][9][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][9][17] = (sum_out[1][9][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][9][17] = (sum_out[2][9][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][9][17] = (sum_out[3][9][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][9][17] = (sum_out[4][9][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][9][17] = (sum_out[5][9][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][9][17] = (sum_out[6][9][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][9][17] = (sum_out[7][9][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][9][17] = (sum_out[8][9][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][9][17] = (sum_out[9][9][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][9][17] = (sum_out[10][9][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][9][17] = (sum_out[11][9][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][9][17] = (sum_out[12][9][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][9][17] = (sum_out[13][9][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][9][17] = (sum_out[14][9][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][9][17] = (sum_out[15][9][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][9][17] = (sum_out[16][9][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][9][17] = (sum_out[17][9][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][9][17] = (sum_out[18][9][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][9][17] = (sum_out[19][9][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][9][18] = (sum_out[0][9][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][9][18] = (sum_out[1][9][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][9][18] = (sum_out[2][9][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][9][18] = (sum_out[3][9][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][9][18] = (sum_out[4][9][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][9][18] = (sum_out[5][9][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][9][18] = (sum_out[6][9][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][9][18] = (sum_out[7][9][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][9][18] = (sum_out[8][9][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][9][18] = (sum_out[9][9][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][9][18] = (sum_out[10][9][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][9][18] = (sum_out[11][9][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][9][18] = (sum_out[12][9][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][9][18] = (sum_out[13][9][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][9][18] = (sum_out[14][9][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][9][18] = (sum_out[15][9][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][9][18] = (sum_out[16][9][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][9][18] = (sum_out[17][9][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][9][18] = (sum_out[18][9][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][9][18] = (sum_out[19][9][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][9][19] = (sum_out[0][9][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][9][19] = (sum_out[1][9][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][9][19] = (sum_out[2][9][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][9][19] = (sum_out[3][9][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][9][19] = (sum_out[4][9][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][9][19] = (sum_out[5][9][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][9][19] = (sum_out[6][9][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][9][19] = (sum_out[7][9][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][9][19] = (sum_out[8][9][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][9][19] = (sum_out[9][9][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][9][19] = (sum_out[10][9][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][9][19] = (sum_out[11][9][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][9][19] = (sum_out[12][9][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][9][19] = (sum_out[13][9][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][9][19] = (sum_out[14][9][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][9][19] = (sum_out[15][9][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][9][19] = (sum_out[16][9][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][9][19] = (sum_out[17][9][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][9][19] = (sum_out[18][9][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][9][19] = (sum_out[19][9][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][9][20] = (sum_out[0][9][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][9][20] = (sum_out[1][9][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][9][20] = (sum_out[2][9][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][9][20] = (sum_out[3][9][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][9][20] = (sum_out[4][9][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][9][20] = (sum_out[5][9][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][9][20] = (sum_out[6][9][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][9][20] = (sum_out[7][9][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][9][20] = (sum_out[8][9][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][9][20] = (sum_out[9][9][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][9][20] = (sum_out[10][9][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][9][20] = (sum_out[11][9][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][9][20] = (sum_out[12][9][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][9][20] = (sum_out[13][9][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][9][20] = (sum_out[14][9][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][9][20] = (sum_out[15][9][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][9][20] = (sum_out[16][9][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][9][20] = (sum_out[17][9][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][9][20] = (sum_out[18][9][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][9][20] = (sum_out[19][9][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][9][21] = (sum_out[0][9][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][9][21] = (sum_out[1][9][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][9][21] = (sum_out[2][9][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][9][21] = (sum_out[3][9][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][9][21] = (sum_out[4][9][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][9][21] = (sum_out[5][9][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][9][21] = (sum_out[6][9][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][9][21] = (sum_out[7][9][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][9][21] = (sum_out[8][9][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][9][21] = (sum_out[9][9][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][9][21] = (sum_out[10][9][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][9][21] = (sum_out[11][9][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][9][21] = (sum_out[12][9][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][9][21] = (sum_out[13][9][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][9][21] = (sum_out[14][9][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][9][21] = (sum_out[15][9][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][9][21] = (sum_out[16][9][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][9][21] = (sum_out[17][9][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][9][21] = (sum_out[18][9][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][9][21] = (sum_out[19][9][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][9][22] = (sum_out[0][9][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][9][22] = (sum_out[1][9][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][9][22] = (sum_out[2][9][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][9][22] = (sum_out[3][9][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][9][22] = (sum_out[4][9][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][9][22] = (sum_out[5][9][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][9][22] = (sum_out[6][9][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][9][22] = (sum_out[7][9][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][9][22] = (sum_out[8][9][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][9][22] = (sum_out[9][9][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][9][22] = (sum_out[10][9][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][9][22] = (sum_out[11][9][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][9][22] = (sum_out[12][9][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][9][22] = (sum_out[13][9][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][9][22] = (sum_out[14][9][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][9][22] = (sum_out[15][9][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][9][22] = (sum_out[16][9][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][9][22] = (sum_out[17][9][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][9][22] = (sum_out[18][9][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][9][22] = (sum_out[19][9][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][9][23] = (sum_out[0][9][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][9][23] = (sum_out[1][9][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][9][23] = (sum_out[2][9][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][9][23] = (sum_out[3][9][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][9][23] = (sum_out[4][9][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][9][23] = (sum_out[5][9][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][9][23] = (sum_out[6][9][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][9][23] = (sum_out[7][9][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][9][23] = (sum_out[8][9][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][9][23] = (sum_out[9][9][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][9][23] = (sum_out[10][9][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][9][23] = (sum_out[11][9][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][9][23] = (sum_out[12][9][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][9][23] = (sum_out[13][9][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][9][23] = (sum_out[14][9][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][9][23] = (sum_out[15][9][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][9][23] = (sum_out[16][9][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][9][23] = (sum_out[17][9][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][9][23] = (sum_out[18][9][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][9][23] = (sum_out[19][9][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][10][0] = (sum_out[0][10][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][10][0] = (sum_out[1][10][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][10][0] = (sum_out[2][10][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][10][0] = (sum_out[3][10][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][10][0] = (sum_out[4][10][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][10][0] = (sum_out[5][10][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][10][0] = (sum_out[6][10][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][10][0] = (sum_out[7][10][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][10][0] = (sum_out[8][10][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][10][0] = (sum_out[9][10][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][10][0] = (sum_out[10][10][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][10][0] = (sum_out[11][10][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][10][0] = (sum_out[12][10][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][10][0] = (sum_out[13][10][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][10][0] = (sum_out[14][10][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][10][0] = (sum_out[15][10][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][10][0] = (sum_out[16][10][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][10][0] = (sum_out[17][10][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][10][0] = (sum_out[18][10][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][10][0] = (sum_out[19][10][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][10][1] = (sum_out[0][10][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][10][1] = (sum_out[1][10][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][10][1] = (sum_out[2][10][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][10][1] = (sum_out[3][10][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][10][1] = (sum_out[4][10][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][10][1] = (sum_out[5][10][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][10][1] = (sum_out[6][10][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][10][1] = (sum_out[7][10][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][10][1] = (sum_out[8][10][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][10][1] = (sum_out[9][10][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][10][1] = (sum_out[10][10][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][10][1] = (sum_out[11][10][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][10][1] = (sum_out[12][10][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][10][1] = (sum_out[13][10][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][10][1] = (sum_out[14][10][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][10][1] = (sum_out[15][10][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][10][1] = (sum_out[16][10][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][10][1] = (sum_out[17][10][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][10][1] = (sum_out[18][10][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][10][1] = (sum_out[19][10][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][10][2] = (sum_out[0][10][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][10][2] = (sum_out[1][10][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][10][2] = (sum_out[2][10][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][10][2] = (sum_out[3][10][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][10][2] = (sum_out[4][10][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][10][2] = (sum_out[5][10][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][10][2] = (sum_out[6][10][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][10][2] = (sum_out[7][10][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][10][2] = (sum_out[8][10][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][10][2] = (sum_out[9][10][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][10][2] = (sum_out[10][10][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][10][2] = (sum_out[11][10][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][10][2] = (sum_out[12][10][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][10][2] = (sum_out[13][10][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][10][2] = (sum_out[14][10][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][10][2] = (sum_out[15][10][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][10][2] = (sum_out[16][10][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][10][2] = (sum_out[17][10][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][10][2] = (sum_out[18][10][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][10][2] = (sum_out[19][10][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][10][3] = (sum_out[0][10][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][10][3] = (sum_out[1][10][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][10][3] = (sum_out[2][10][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][10][3] = (sum_out[3][10][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][10][3] = (sum_out[4][10][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][10][3] = (sum_out[5][10][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][10][3] = (sum_out[6][10][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][10][3] = (sum_out[7][10][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][10][3] = (sum_out[8][10][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][10][3] = (sum_out[9][10][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][10][3] = (sum_out[10][10][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][10][3] = (sum_out[11][10][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][10][3] = (sum_out[12][10][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][10][3] = (sum_out[13][10][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][10][3] = (sum_out[14][10][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][10][3] = (sum_out[15][10][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][10][3] = (sum_out[16][10][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][10][3] = (sum_out[17][10][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][10][3] = (sum_out[18][10][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][10][3] = (sum_out[19][10][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][10][4] = (sum_out[0][10][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][10][4] = (sum_out[1][10][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][10][4] = (sum_out[2][10][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][10][4] = (sum_out[3][10][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][10][4] = (sum_out[4][10][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][10][4] = (sum_out[5][10][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][10][4] = (sum_out[6][10][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][10][4] = (sum_out[7][10][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][10][4] = (sum_out[8][10][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][10][4] = (sum_out[9][10][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][10][4] = (sum_out[10][10][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][10][4] = (sum_out[11][10][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][10][4] = (sum_out[12][10][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][10][4] = (sum_out[13][10][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][10][4] = (sum_out[14][10][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][10][4] = (sum_out[15][10][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][10][4] = (sum_out[16][10][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][10][4] = (sum_out[17][10][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][10][4] = (sum_out[18][10][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][10][4] = (sum_out[19][10][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][10][5] = (sum_out[0][10][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][10][5] = (sum_out[1][10][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][10][5] = (sum_out[2][10][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][10][5] = (sum_out[3][10][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][10][5] = (sum_out[4][10][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][10][5] = (sum_out[5][10][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][10][5] = (sum_out[6][10][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][10][5] = (sum_out[7][10][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][10][5] = (sum_out[8][10][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][10][5] = (sum_out[9][10][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][10][5] = (sum_out[10][10][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][10][5] = (sum_out[11][10][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][10][5] = (sum_out[12][10][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][10][5] = (sum_out[13][10][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][10][5] = (sum_out[14][10][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][10][5] = (sum_out[15][10][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][10][5] = (sum_out[16][10][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][10][5] = (sum_out[17][10][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][10][5] = (sum_out[18][10][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][10][5] = (sum_out[19][10][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][10][6] = (sum_out[0][10][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][10][6] = (sum_out[1][10][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][10][6] = (sum_out[2][10][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][10][6] = (sum_out[3][10][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][10][6] = (sum_out[4][10][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][10][6] = (sum_out[5][10][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][10][6] = (sum_out[6][10][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][10][6] = (sum_out[7][10][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][10][6] = (sum_out[8][10][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][10][6] = (sum_out[9][10][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][10][6] = (sum_out[10][10][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][10][6] = (sum_out[11][10][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][10][6] = (sum_out[12][10][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][10][6] = (sum_out[13][10][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][10][6] = (sum_out[14][10][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][10][6] = (sum_out[15][10][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][10][6] = (sum_out[16][10][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][10][6] = (sum_out[17][10][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][10][6] = (sum_out[18][10][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][10][6] = (sum_out[19][10][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][10][7] = (sum_out[0][10][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][10][7] = (sum_out[1][10][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][10][7] = (sum_out[2][10][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][10][7] = (sum_out[3][10][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][10][7] = (sum_out[4][10][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][10][7] = (sum_out[5][10][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][10][7] = (sum_out[6][10][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][10][7] = (sum_out[7][10][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][10][7] = (sum_out[8][10][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][10][7] = (sum_out[9][10][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][10][7] = (sum_out[10][10][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][10][7] = (sum_out[11][10][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][10][7] = (sum_out[12][10][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][10][7] = (sum_out[13][10][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][10][7] = (sum_out[14][10][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][10][7] = (sum_out[15][10][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][10][7] = (sum_out[16][10][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][10][7] = (sum_out[17][10][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][10][7] = (sum_out[18][10][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][10][7] = (sum_out[19][10][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][10][8] = (sum_out[0][10][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][10][8] = (sum_out[1][10][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][10][8] = (sum_out[2][10][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][10][8] = (sum_out[3][10][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][10][8] = (sum_out[4][10][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][10][8] = (sum_out[5][10][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][10][8] = (sum_out[6][10][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][10][8] = (sum_out[7][10][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][10][8] = (sum_out[8][10][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][10][8] = (sum_out[9][10][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][10][8] = (sum_out[10][10][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][10][8] = (sum_out[11][10][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][10][8] = (sum_out[12][10][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][10][8] = (sum_out[13][10][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][10][8] = (sum_out[14][10][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][10][8] = (sum_out[15][10][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][10][8] = (sum_out[16][10][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][10][8] = (sum_out[17][10][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][10][8] = (sum_out[18][10][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][10][8] = (sum_out[19][10][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][10][9] = (sum_out[0][10][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][10][9] = (sum_out[1][10][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][10][9] = (sum_out[2][10][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][10][9] = (sum_out[3][10][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][10][9] = (sum_out[4][10][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][10][9] = (sum_out[5][10][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][10][9] = (sum_out[6][10][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][10][9] = (sum_out[7][10][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][10][9] = (sum_out[8][10][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][10][9] = (sum_out[9][10][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][10][9] = (sum_out[10][10][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][10][9] = (sum_out[11][10][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][10][9] = (sum_out[12][10][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][10][9] = (sum_out[13][10][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][10][9] = (sum_out[14][10][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][10][9] = (sum_out[15][10][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][10][9] = (sum_out[16][10][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][10][9] = (sum_out[17][10][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][10][9] = (sum_out[18][10][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][10][9] = (sum_out[19][10][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][10][10] = (sum_out[0][10][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][10][10] = (sum_out[1][10][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][10][10] = (sum_out[2][10][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][10][10] = (sum_out[3][10][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][10][10] = (sum_out[4][10][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][10][10] = (sum_out[5][10][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][10][10] = (sum_out[6][10][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][10][10] = (sum_out[7][10][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][10][10] = (sum_out[8][10][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][10][10] = (sum_out[9][10][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][10][10] = (sum_out[10][10][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][10][10] = (sum_out[11][10][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][10][10] = (sum_out[12][10][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][10][10] = (sum_out[13][10][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][10][10] = (sum_out[14][10][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][10][10] = (sum_out[15][10][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][10][10] = (sum_out[16][10][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][10][10] = (sum_out[17][10][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][10][10] = (sum_out[18][10][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][10][10] = (sum_out[19][10][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][10][11] = (sum_out[0][10][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][10][11] = (sum_out[1][10][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][10][11] = (sum_out[2][10][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][10][11] = (sum_out[3][10][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][10][11] = (sum_out[4][10][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][10][11] = (sum_out[5][10][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][10][11] = (sum_out[6][10][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][10][11] = (sum_out[7][10][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][10][11] = (sum_out[8][10][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][10][11] = (sum_out[9][10][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][10][11] = (sum_out[10][10][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][10][11] = (sum_out[11][10][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][10][11] = (sum_out[12][10][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][10][11] = (sum_out[13][10][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][10][11] = (sum_out[14][10][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][10][11] = (sum_out[15][10][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][10][11] = (sum_out[16][10][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][10][11] = (sum_out[17][10][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][10][11] = (sum_out[18][10][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][10][11] = (sum_out[19][10][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][10][12] = (sum_out[0][10][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][10][12] = (sum_out[1][10][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][10][12] = (sum_out[2][10][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][10][12] = (sum_out[3][10][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][10][12] = (sum_out[4][10][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][10][12] = (sum_out[5][10][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][10][12] = (sum_out[6][10][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][10][12] = (sum_out[7][10][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][10][12] = (sum_out[8][10][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][10][12] = (sum_out[9][10][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][10][12] = (sum_out[10][10][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][10][12] = (sum_out[11][10][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][10][12] = (sum_out[12][10][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][10][12] = (sum_out[13][10][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][10][12] = (sum_out[14][10][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][10][12] = (sum_out[15][10][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][10][12] = (sum_out[16][10][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][10][12] = (sum_out[17][10][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][10][12] = (sum_out[18][10][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][10][12] = (sum_out[19][10][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][10][13] = (sum_out[0][10][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][10][13] = (sum_out[1][10][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][10][13] = (sum_out[2][10][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][10][13] = (sum_out[3][10][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][10][13] = (sum_out[4][10][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][10][13] = (sum_out[5][10][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][10][13] = (sum_out[6][10][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][10][13] = (sum_out[7][10][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][10][13] = (sum_out[8][10][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][10][13] = (sum_out[9][10][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][10][13] = (sum_out[10][10][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][10][13] = (sum_out[11][10][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][10][13] = (sum_out[12][10][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][10][13] = (sum_out[13][10][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][10][13] = (sum_out[14][10][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][10][13] = (sum_out[15][10][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][10][13] = (sum_out[16][10][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][10][13] = (sum_out[17][10][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][10][13] = (sum_out[18][10][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][10][13] = (sum_out[19][10][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][10][14] = (sum_out[0][10][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][10][14] = (sum_out[1][10][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][10][14] = (sum_out[2][10][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][10][14] = (sum_out[3][10][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][10][14] = (sum_out[4][10][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][10][14] = (sum_out[5][10][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][10][14] = (sum_out[6][10][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][10][14] = (sum_out[7][10][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][10][14] = (sum_out[8][10][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][10][14] = (sum_out[9][10][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][10][14] = (sum_out[10][10][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][10][14] = (sum_out[11][10][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][10][14] = (sum_out[12][10][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][10][14] = (sum_out[13][10][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][10][14] = (sum_out[14][10][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][10][14] = (sum_out[15][10][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][10][14] = (sum_out[16][10][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][10][14] = (sum_out[17][10][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][10][14] = (sum_out[18][10][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][10][14] = (sum_out[19][10][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][10][15] = (sum_out[0][10][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][10][15] = (sum_out[1][10][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][10][15] = (sum_out[2][10][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][10][15] = (sum_out[3][10][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][10][15] = (sum_out[4][10][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][10][15] = (sum_out[5][10][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][10][15] = (sum_out[6][10][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][10][15] = (sum_out[7][10][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][10][15] = (sum_out[8][10][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][10][15] = (sum_out[9][10][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][10][15] = (sum_out[10][10][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][10][15] = (sum_out[11][10][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][10][15] = (sum_out[12][10][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][10][15] = (sum_out[13][10][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][10][15] = (sum_out[14][10][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][10][15] = (sum_out[15][10][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][10][15] = (sum_out[16][10][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][10][15] = (sum_out[17][10][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][10][15] = (sum_out[18][10][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][10][15] = (sum_out[19][10][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][10][16] = (sum_out[0][10][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][10][16] = (sum_out[1][10][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][10][16] = (sum_out[2][10][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][10][16] = (sum_out[3][10][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][10][16] = (sum_out[4][10][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][10][16] = (sum_out[5][10][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][10][16] = (sum_out[6][10][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][10][16] = (sum_out[7][10][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][10][16] = (sum_out[8][10][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][10][16] = (sum_out[9][10][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][10][16] = (sum_out[10][10][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][10][16] = (sum_out[11][10][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][10][16] = (sum_out[12][10][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][10][16] = (sum_out[13][10][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][10][16] = (sum_out[14][10][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][10][16] = (sum_out[15][10][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][10][16] = (sum_out[16][10][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][10][16] = (sum_out[17][10][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][10][16] = (sum_out[18][10][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][10][16] = (sum_out[19][10][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][10][17] = (sum_out[0][10][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][10][17] = (sum_out[1][10][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][10][17] = (sum_out[2][10][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][10][17] = (sum_out[3][10][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][10][17] = (sum_out[4][10][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][10][17] = (sum_out[5][10][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][10][17] = (sum_out[6][10][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][10][17] = (sum_out[7][10][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][10][17] = (sum_out[8][10][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][10][17] = (sum_out[9][10][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][10][17] = (sum_out[10][10][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][10][17] = (sum_out[11][10][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][10][17] = (sum_out[12][10][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][10][17] = (sum_out[13][10][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][10][17] = (sum_out[14][10][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][10][17] = (sum_out[15][10][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][10][17] = (sum_out[16][10][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][10][17] = (sum_out[17][10][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][10][17] = (sum_out[18][10][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][10][17] = (sum_out[19][10][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][10][18] = (sum_out[0][10][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][10][18] = (sum_out[1][10][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][10][18] = (sum_out[2][10][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][10][18] = (sum_out[3][10][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][10][18] = (sum_out[4][10][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][10][18] = (sum_out[5][10][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][10][18] = (sum_out[6][10][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][10][18] = (sum_out[7][10][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][10][18] = (sum_out[8][10][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][10][18] = (sum_out[9][10][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][10][18] = (sum_out[10][10][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][10][18] = (sum_out[11][10][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][10][18] = (sum_out[12][10][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][10][18] = (sum_out[13][10][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][10][18] = (sum_out[14][10][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][10][18] = (sum_out[15][10][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][10][18] = (sum_out[16][10][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][10][18] = (sum_out[17][10][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][10][18] = (sum_out[18][10][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][10][18] = (sum_out[19][10][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][10][19] = (sum_out[0][10][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][10][19] = (sum_out[1][10][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][10][19] = (sum_out[2][10][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][10][19] = (sum_out[3][10][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][10][19] = (sum_out[4][10][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][10][19] = (sum_out[5][10][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][10][19] = (sum_out[6][10][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][10][19] = (sum_out[7][10][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][10][19] = (sum_out[8][10][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][10][19] = (sum_out[9][10][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][10][19] = (sum_out[10][10][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][10][19] = (sum_out[11][10][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][10][19] = (sum_out[12][10][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][10][19] = (sum_out[13][10][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][10][19] = (sum_out[14][10][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][10][19] = (sum_out[15][10][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][10][19] = (sum_out[16][10][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][10][19] = (sum_out[17][10][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][10][19] = (sum_out[18][10][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][10][19] = (sum_out[19][10][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][10][20] = (sum_out[0][10][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][10][20] = (sum_out[1][10][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][10][20] = (sum_out[2][10][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][10][20] = (sum_out[3][10][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][10][20] = (sum_out[4][10][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][10][20] = (sum_out[5][10][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][10][20] = (sum_out[6][10][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][10][20] = (sum_out[7][10][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][10][20] = (sum_out[8][10][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][10][20] = (sum_out[9][10][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][10][20] = (sum_out[10][10][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][10][20] = (sum_out[11][10][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][10][20] = (sum_out[12][10][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][10][20] = (sum_out[13][10][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][10][20] = (sum_out[14][10][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][10][20] = (sum_out[15][10][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][10][20] = (sum_out[16][10][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][10][20] = (sum_out[17][10][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][10][20] = (sum_out[18][10][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][10][20] = (sum_out[19][10][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][10][21] = (sum_out[0][10][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][10][21] = (sum_out[1][10][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][10][21] = (sum_out[2][10][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][10][21] = (sum_out[3][10][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][10][21] = (sum_out[4][10][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][10][21] = (sum_out[5][10][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][10][21] = (sum_out[6][10][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][10][21] = (sum_out[7][10][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][10][21] = (sum_out[8][10][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][10][21] = (sum_out[9][10][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][10][21] = (sum_out[10][10][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][10][21] = (sum_out[11][10][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][10][21] = (sum_out[12][10][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][10][21] = (sum_out[13][10][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][10][21] = (sum_out[14][10][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][10][21] = (sum_out[15][10][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][10][21] = (sum_out[16][10][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][10][21] = (sum_out[17][10][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][10][21] = (sum_out[18][10][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][10][21] = (sum_out[19][10][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][10][22] = (sum_out[0][10][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][10][22] = (sum_out[1][10][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][10][22] = (sum_out[2][10][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][10][22] = (sum_out[3][10][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][10][22] = (sum_out[4][10][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][10][22] = (sum_out[5][10][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][10][22] = (sum_out[6][10][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][10][22] = (sum_out[7][10][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][10][22] = (sum_out[8][10][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][10][22] = (sum_out[9][10][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][10][22] = (sum_out[10][10][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][10][22] = (sum_out[11][10][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][10][22] = (sum_out[12][10][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][10][22] = (sum_out[13][10][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][10][22] = (sum_out[14][10][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][10][22] = (sum_out[15][10][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][10][22] = (sum_out[16][10][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][10][22] = (sum_out[17][10][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][10][22] = (sum_out[18][10][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][10][22] = (sum_out[19][10][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][10][23] = (sum_out[0][10][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][10][23] = (sum_out[1][10][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][10][23] = (sum_out[2][10][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][10][23] = (sum_out[3][10][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][10][23] = (sum_out[4][10][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][10][23] = (sum_out[5][10][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][10][23] = (sum_out[6][10][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][10][23] = (sum_out[7][10][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][10][23] = (sum_out[8][10][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][10][23] = (sum_out[9][10][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][10][23] = (sum_out[10][10][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][10][23] = (sum_out[11][10][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][10][23] = (sum_out[12][10][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][10][23] = (sum_out[13][10][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][10][23] = (sum_out[14][10][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][10][23] = (sum_out[15][10][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][10][23] = (sum_out[16][10][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][10][23] = (sum_out[17][10][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][10][23] = (sum_out[18][10][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][10][23] = (sum_out[19][10][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][11][0] = (sum_out[0][11][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][11][0] = (sum_out[1][11][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][11][0] = (sum_out[2][11][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][11][0] = (sum_out[3][11][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][11][0] = (sum_out[4][11][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][11][0] = (sum_out[5][11][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][11][0] = (sum_out[6][11][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][11][0] = (sum_out[7][11][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][11][0] = (sum_out[8][11][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][11][0] = (sum_out[9][11][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][11][0] = (sum_out[10][11][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][11][0] = (sum_out[11][11][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][11][0] = (sum_out[12][11][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][11][0] = (sum_out[13][11][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][11][0] = (sum_out[14][11][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][11][0] = (sum_out[15][11][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][11][0] = (sum_out[16][11][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][11][0] = (sum_out[17][11][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][11][0] = (sum_out[18][11][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][11][0] = (sum_out[19][11][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][11][1] = (sum_out[0][11][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][11][1] = (sum_out[1][11][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][11][1] = (sum_out[2][11][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][11][1] = (sum_out[3][11][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][11][1] = (sum_out[4][11][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][11][1] = (sum_out[5][11][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][11][1] = (sum_out[6][11][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][11][1] = (sum_out[7][11][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][11][1] = (sum_out[8][11][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][11][1] = (sum_out[9][11][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][11][1] = (sum_out[10][11][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][11][1] = (sum_out[11][11][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][11][1] = (sum_out[12][11][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][11][1] = (sum_out[13][11][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][11][1] = (sum_out[14][11][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][11][1] = (sum_out[15][11][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][11][1] = (sum_out[16][11][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][11][1] = (sum_out[17][11][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][11][1] = (sum_out[18][11][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][11][1] = (sum_out[19][11][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][11][2] = (sum_out[0][11][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][11][2] = (sum_out[1][11][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][11][2] = (sum_out[2][11][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][11][2] = (sum_out[3][11][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][11][2] = (sum_out[4][11][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][11][2] = (sum_out[5][11][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][11][2] = (sum_out[6][11][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][11][2] = (sum_out[7][11][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][11][2] = (sum_out[8][11][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][11][2] = (sum_out[9][11][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][11][2] = (sum_out[10][11][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][11][2] = (sum_out[11][11][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][11][2] = (sum_out[12][11][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][11][2] = (sum_out[13][11][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][11][2] = (sum_out[14][11][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][11][2] = (sum_out[15][11][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][11][2] = (sum_out[16][11][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][11][2] = (sum_out[17][11][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][11][2] = (sum_out[18][11][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][11][2] = (sum_out[19][11][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][11][3] = (sum_out[0][11][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][11][3] = (sum_out[1][11][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][11][3] = (sum_out[2][11][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][11][3] = (sum_out[3][11][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][11][3] = (sum_out[4][11][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][11][3] = (sum_out[5][11][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][11][3] = (sum_out[6][11][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][11][3] = (sum_out[7][11][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][11][3] = (sum_out[8][11][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][11][3] = (sum_out[9][11][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][11][3] = (sum_out[10][11][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][11][3] = (sum_out[11][11][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][11][3] = (sum_out[12][11][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][11][3] = (sum_out[13][11][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][11][3] = (sum_out[14][11][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][11][3] = (sum_out[15][11][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][11][3] = (sum_out[16][11][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][11][3] = (sum_out[17][11][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][11][3] = (sum_out[18][11][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][11][3] = (sum_out[19][11][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][11][4] = (sum_out[0][11][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][11][4] = (sum_out[1][11][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][11][4] = (sum_out[2][11][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][11][4] = (sum_out[3][11][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][11][4] = (sum_out[4][11][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][11][4] = (sum_out[5][11][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][11][4] = (sum_out[6][11][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][11][4] = (sum_out[7][11][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][11][4] = (sum_out[8][11][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][11][4] = (sum_out[9][11][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][11][4] = (sum_out[10][11][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][11][4] = (sum_out[11][11][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][11][4] = (sum_out[12][11][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][11][4] = (sum_out[13][11][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][11][4] = (sum_out[14][11][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][11][4] = (sum_out[15][11][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][11][4] = (sum_out[16][11][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][11][4] = (sum_out[17][11][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][11][4] = (sum_out[18][11][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][11][4] = (sum_out[19][11][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][11][5] = (sum_out[0][11][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][11][5] = (sum_out[1][11][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][11][5] = (sum_out[2][11][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][11][5] = (sum_out[3][11][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][11][5] = (sum_out[4][11][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][11][5] = (sum_out[5][11][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][11][5] = (sum_out[6][11][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][11][5] = (sum_out[7][11][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][11][5] = (sum_out[8][11][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][11][5] = (sum_out[9][11][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][11][5] = (sum_out[10][11][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][11][5] = (sum_out[11][11][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][11][5] = (sum_out[12][11][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][11][5] = (sum_out[13][11][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][11][5] = (sum_out[14][11][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][11][5] = (sum_out[15][11][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][11][5] = (sum_out[16][11][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][11][5] = (sum_out[17][11][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][11][5] = (sum_out[18][11][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][11][5] = (sum_out[19][11][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][11][6] = (sum_out[0][11][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][11][6] = (sum_out[1][11][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][11][6] = (sum_out[2][11][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][11][6] = (sum_out[3][11][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][11][6] = (sum_out[4][11][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][11][6] = (sum_out[5][11][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][11][6] = (sum_out[6][11][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][11][6] = (sum_out[7][11][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][11][6] = (sum_out[8][11][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][11][6] = (sum_out[9][11][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][11][6] = (sum_out[10][11][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][11][6] = (sum_out[11][11][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][11][6] = (sum_out[12][11][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][11][6] = (sum_out[13][11][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][11][6] = (sum_out[14][11][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][11][6] = (sum_out[15][11][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][11][6] = (sum_out[16][11][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][11][6] = (sum_out[17][11][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][11][6] = (sum_out[18][11][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][11][6] = (sum_out[19][11][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][11][7] = (sum_out[0][11][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][11][7] = (sum_out[1][11][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][11][7] = (sum_out[2][11][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][11][7] = (sum_out[3][11][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][11][7] = (sum_out[4][11][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][11][7] = (sum_out[5][11][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][11][7] = (sum_out[6][11][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][11][7] = (sum_out[7][11][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][11][7] = (sum_out[8][11][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][11][7] = (sum_out[9][11][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][11][7] = (sum_out[10][11][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][11][7] = (sum_out[11][11][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][11][7] = (sum_out[12][11][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][11][7] = (sum_out[13][11][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][11][7] = (sum_out[14][11][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][11][7] = (sum_out[15][11][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][11][7] = (sum_out[16][11][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][11][7] = (sum_out[17][11][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][11][7] = (sum_out[18][11][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][11][7] = (sum_out[19][11][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][11][8] = (sum_out[0][11][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][11][8] = (sum_out[1][11][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][11][8] = (sum_out[2][11][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][11][8] = (sum_out[3][11][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][11][8] = (sum_out[4][11][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][11][8] = (sum_out[5][11][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][11][8] = (sum_out[6][11][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][11][8] = (sum_out[7][11][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][11][8] = (sum_out[8][11][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][11][8] = (sum_out[9][11][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][11][8] = (sum_out[10][11][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][11][8] = (sum_out[11][11][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][11][8] = (sum_out[12][11][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][11][8] = (sum_out[13][11][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][11][8] = (sum_out[14][11][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][11][8] = (sum_out[15][11][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][11][8] = (sum_out[16][11][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][11][8] = (sum_out[17][11][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][11][8] = (sum_out[18][11][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][11][8] = (sum_out[19][11][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][11][9] = (sum_out[0][11][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][11][9] = (sum_out[1][11][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][11][9] = (sum_out[2][11][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][11][9] = (sum_out[3][11][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][11][9] = (sum_out[4][11][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][11][9] = (sum_out[5][11][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][11][9] = (sum_out[6][11][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][11][9] = (sum_out[7][11][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][11][9] = (sum_out[8][11][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][11][9] = (sum_out[9][11][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][11][9] = (sum_out[10][11][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][11][9] = (sum_out[11][11][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][11][9] = (sum_out[12][11][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][11][9] = (sum_out[13][11][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][11][9] = (sum_out[14][11][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][11][9] = (sum_out[15][11][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][11][9] = (sum_out[16][11][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][11][9] = (sum_out[17][11][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][11][9] = (sum_out[18][11][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][11][9] = (sum_out[19][11][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][11][10] = (sum_out[0][11][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][11][10] = (sum_out[1][11][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][11][10] = (sum_out[2][11][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][11][10] = (sum_out[3][11][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][11][10] = (sum_out[4][11][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][11][10] = (sum_out[5][11][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][11][10] = (sum_out[6][11][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][11][10] = (sum_out[7][11][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][11][10] = (sum_out[8][11][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][11][10] = (sum_out[9][11][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][11][10] = (sum_out[10][11][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][11][10] = (sum_out[11][11][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][11][10] = (sum_out[12][11][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][11][10] = (sum_out[13][11][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][11][10] = (sum_out[14][11][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][11][10] = (sum_out[15][11][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][11][10] = (sum_out[16][11][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][11][10] = (sum_out[17][11][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][11][10] = (sum_out[18][11][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][11][10] = (sum_out[19][11][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][11][11] = (sum_out[0][11][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][11][11] = (sum_out[1][11][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][11][11] = (sum_out[2][11][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][11][11] = (sum_out[3][11][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][11][11] = (sum_out[4][11][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][11][11] = (sum_out[5][11][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][11][11] = (sum_out[6][11][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][11][11] = (sum_out[7][11][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][11][11] = (sum_out[8][11][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][11][11] = (sum_out[9][11][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][11][11] = (sum_out[10][11][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][11][11] = (sum_out[11][11][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][11][11] = (sum_out[12][11][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][11][11] = (sum_out[13][11][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][11][11] = (sum_out[14][11][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][11][11] = (sum_out[15][11][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][11][11] = (sum_out[16][11][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][11][11] = (sum_out[17][11][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][11][11] = (sum_out[18][11][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][11][11] = (sum_out[19][11][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][11][12] = (sum_out[0][11][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][11][12] = (sum_out[1][11][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][11][12] = (sum_out[2][11][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][11][12] = (sum_out[3][11][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][11][12] = (sum_out[4][11][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][11][12] = (sum_out[5][11][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][11][12] = (sum_out[6][11][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][11][12] = (sum_out[7][11][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][11][12] = (sum_out[8][11][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][11][12] = (sum_out[9][11][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][11][12] = (sum_out[10][11][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][11][12] = (sum_out[11][11][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][11][12] = (sum_out[12][11][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][11][12] = (sum_out[13][11][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][11][12] = (sum_out[14][11][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][11][12] = (sum_out[15][11][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][11][12] = (sum_out[16][11][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][11][12] = (sum_out[17][11][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][11][12] = (sum_out[18][11][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][11][12] = (sum_out[19][11][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][11][13] = (sum_out[0][11][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][11][13] = (sum_out[1][11][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][11][13] = (sum_out[2][11][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][11][13] = (sum_out[3][11][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][11][13] = (sum_out[4][11][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][11][13] = (sum_out[5][11][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][11][13] = (sum_out[6][11][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][11][13] = (sum_out[7][11][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][11][13] = (sum_out[8][11][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][11][13] = (sum_out[9][11][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][11][13] = (sum_out[10][11][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][11][13] = (sum_out[11][11][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][11][13] = (sum_out[12][11][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][11][13] = (sum_out[13][11][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][11][13] = (sum_out[14][11][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][11][13] = (sum_out[15][11][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][11][13] = (sum_out[16][11][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][11][13] = (sum_out[17][11][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][11][13] = (sum_out[18][11][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][11][13] = (sum_out[19][11][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][11][14] = (sum_out[0][11][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][11][14] = (sum_out[1][11][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][11][14] = (sum_out[2][11][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][11][14] = (sum_out[3][11][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][11][14] = (sum_out[4][11][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][11][14] = (sum_out[5][11][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][11][14] = (sum_out[6][11][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][11][14] = (sum_out[7][11][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][11][14] = (sum_out[8][11][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][11][14] = (sum_out[9][11][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][11][14] = (sum_out[10][11][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][11][14] = (sum_out[11][11][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][11][14] = (sum_out[12][11][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][11][14] = (sum_out[13][11][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][11][14] = (sum_out[14][11][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][11][14] = (sum_out[15][11][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][11][14] = (sum_out[16][11][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][11][14] = (sum_out[17][11][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][11][14] = (sum_out[18][11][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][11][14] = (sum_out[19][11][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][11][15] = (sum_out[0][11][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][11][15] = (sum_out[1][11][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][11][15] = (sum_out[2][11][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][11][15] = (sum_out[3][11][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][11][15] = (sum_out[4][11][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][11][15] = (sum_out[5][11][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][11][15] = (sum_out[6][11][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][11][15] = (sum_out[7][11][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][11][15] = (sum_out[8][11][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][11][15] = (sum_out[9][11][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][11][15] = (sum_out[10][11][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][11][15] = (sum_out[11][11][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][11][15] = (sum_out[12][11][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][11][15] = (sum_out[13][11][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][11][15] = (sum_out[14][11][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][11][15] = (sum_out[15][11][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][11][15] = (sum_out[16][11][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][11][15] = (sum_out[17][11][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][11][15] = (sum_out[18][11][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][11][15] = (sum_out[19][11][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][11][16] = (sum_out[0][11][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][11][16] = (sum_out[1][11][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][11][16] = (sum_out[2][11][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][11][16] = (sum_out[3][11][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][11][16] = (sum_out[4][11][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][11][16] = (sum_out[5][11][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][11][16] = (sum_out[6][11][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][11][16] = (sum_out[7][11][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][11][16] = (sum_out[8][11][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][11][16] = (sum_out[9][11][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][11][16] = (sum_out[10][11][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][11][16] = (sum_out[11][11][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][11][16] = (sum_out[12][11][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][11][16] = (sum_out[13][11][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][11][16] = (sum_out[14][11][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][11][16] = (sum_out[15][11][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][11][16] = (sum_out[16][11][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][11][16] = (sum_out[17][11][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][11][16] = (sum_out[18][11][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][11][16] = (sum_out[19][11][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][11][17] = (sum_out[0][11][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][11][17] = (sum_out[1][11][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][11][17] = (sum_out[2][11][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][11][17] = (sum_out[3][11][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][11][17] = (sum_out[4][11][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][11][17] = (sum_out[5][11][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][11][17] = (sum_out[6][11][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][11][17] = (sum_out[7][11][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][11][17] = (sum_out[8][11][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][11][17] = (sum_out[9][11][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][11][17] = (sum_out[10][11][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][11][17] = (sum_out[11][11][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][11][17] = (sum_out[12][11][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][11][17] = (sum_out[13][11][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][11][17] = (sum_out[14][11][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][11][17] = (sum_out[15][11][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][11][17] = (sum_out[16][11][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][11][17] = (sum_out[17][11][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][11][17] = (sum_out[18][11][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][11][17] = (sum_out[19][11][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][11][18] = (sum_out[0][11][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][11][18] = (sum_out[1][11][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][11][18] = (sum_out[2][11][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][11][18] = (sum_out[3][11][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][11][18] = (sum_out[4][11][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][11][18] = (sum_out[5][11][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][11][18] = (sum_out[6][11][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][11][18] = (sum_out[7][11][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][11][18] = (sum_out[8][11][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][11][18] = (sum_out[9][11][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][11][18] = (sum_out[10][11][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][11][18] = (sum_out[11][11][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][11][18] = (sum_out[12][11][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][11][18] = (sum_out[13][11][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][11][18] = (sum_out[14][11][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][11][18] = (sum_out[15][11][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][11][18] = (sum_out[16][11][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][11][18] = (sum_out[17][11][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][11][18] = (sum_out[18][11][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][11][18] = (sum_out[19][11][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][11][19] = (sum_out[0][11][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][11][19] = (sum_out[1][11][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][11][19] = (sum_out[2][11][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][11][19] = (sum_out[3][11][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][11][19] = (sum_out[4][11][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][11][19] = (sum_out[5][11][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][11][19] = (sum_out[6][11][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][11][19] = (sum_out[7][11][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][11][19] = (sum_out[8][11][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][11][19] = (sum_out[9][11][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][11][19] = (sum_out[10][11][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][11][19] = (sum_out[11][11][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][11][19] = (sum_out[12][11][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][11][19] = (sum_out[13][11][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][11][19] = (sum_out[14][11][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][11][19] = (sum_out[15][11][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][11][19] = (sum_out[16][11][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][11][19] = (sum_out[17][11][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][11][19] = (sum_out[18][11][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][11][19] = (sum_out[19][11][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][11][20] = (sum_out[0][11][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][11][20] = (sum_out[1][11][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][11][20] = (sum_out[2][11][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][11][20] = (sum_out[3][11][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][11][20] = (sum_out[4][11][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][11][20] = (sum_out[5][11][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][11][20] = (sum_out[6][11][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][11][20] = (sum_out[7][11][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][11][20] = (sum_out[8][11][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][11][20] = (sum_out[9][11][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][11][20] = (sum_out[10][11][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][11][20] = (sum_out[11][11][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][11][20] = (sum_out[12][11][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][11][20] = (sum_out[13][11][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][11][20] = (sum_out[14][11][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][11][20] = (sum_out[15][11][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][11][20] = (sum_out[16][11][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][11][20] = (sum_out[17][11][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][11][20] = (sum_out[18][11][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][11][20] = (sum_out[19][11][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][11][21] = (sum_out[0][11][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][11][21] = (sum_out[1][11][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][11][21] = (sum_out[2][11][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][11][21] = (sum_out[3][11][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][11][21] = (sum_out[4][11][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][11][21] = (sum_out[5][11][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][11][21] = (sum_out[6][11][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][11][21] = (sum_out[7][11][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][11][21] = (sum_out[8][11][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][11][21] = (sum_out[9][11][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][11][21] = (sum_out[10][11][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][11][21] = (sum_out[11][11][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][11][21] = (sum_out[12][11][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][11][21] = (sum_out[13][11][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][11][21] = (sum_out[14][11][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][11][21] = (sum_out[15][11][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][11][21] = (sum_out[16][11][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][11][21] = (sum_out[17][11][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][11][21] = (sum_out[18][11][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][11][21] = (sum_out[19][11][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][11][22] = (sum_out[0][11][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][11][22] = (sum_out[1][11][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][11][22] = (sum_out[2][11][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][11][22] = (sum_out[3][11][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][11][22] = (sum_out[4][11][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][11][22] = (sum_out[5][11][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][11][22] = (sum_out[6][11][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][11][22] = (sum_out[7][11][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][11][22] = (sum_out[8][11][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][11][22] = (sum_out[9][11][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][11][22] = (sum_out[10][11][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][11][22] = (sum_out[11][11][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][11][22] = (sum_out[12][11][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][11][22] = (sum_out[13][11][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][11][22] = (sum_out[14][11][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][11][22] = (sum_out[15][11][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][11][22] = (sum_out[16][11][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][11][22] = (sum_out[17][11][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][11][22] = (sum_out[18][11][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][11][22] = (sum_out[19][11][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][11][23] = (sum_out[0][11][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][11][23] = (sum_out[1][11][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][11][23] = (sum_out[2][11][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][11][23] = (sum_out[3][11][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][11][23] = (sum_out[4][11][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][11][23] = (sum_out[5][11][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][11][23] = (sum_out[6][11][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][11][23] = (sum_out[7][11][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][11][23] = (sum_out[8][11][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][11][23] = (sum_out[9][11][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][11][23] = (sum_out[10][11][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][11][23] = (sum_out[11][11][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][11][23] = (sum_out[12][11][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][11][23] = (sum_out[13][11][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][11][23] = (sum_out[14][11][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][11][23] = (sum_out[15][11][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][11][23] = (sum_out[16][11][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][11][23] = (sum_out[17][11][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][11][23] = (sum_out[18][11][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][11][23] = (sum_out[19][11][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][12][0] = (sum_out[0][12][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][12][0] = (sum_out[1][12][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][12][0] = (sum_out[2][12][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][12][0] = (sum_out[3][12][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][12][0] = (sum_out[4][12][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][12][0] = (sum_out[5][12][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][12][0] = (sum_out[6][12][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][12][0] = (sum_out[7][12][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][12][0] = (sum_out[8][12][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][12][0] = (sum_out[9][12][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][12][0] = (sum_out[10][12][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][12][0] = (sum_out[11][12][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][12][0] = (sum_out[12][12][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][12][0] = (sum_out[13][12][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][12][0] = (sum_out[14][12][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][12][0] = (sum_out[15][12][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][12][0] = (sum_out[16][12][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][12][0] = (sum_out[17][12][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][12][0] = (sum_out[18][12][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][12][0] = (sum_out[19][12][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][12][1] = (sum_out[0][12][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][12][1] = (sum_out[1][12][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][12][1] = (sum_out[2][12][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][12][1] = (sum_out[3][12][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][12][1] = (sum_out[4][12][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][12][1] = (sum_out[5][12][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][12][1] = (sum_out[6][12][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][12][1] = (sum_out[7][12][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][12][1] = (sum_out[8][12][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][12][1] = (sum_out[9][12][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][12][1] = (sum_out[10][12][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][12][1] = (sum_out[11][12][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][12][1] = (sum_out[12][12][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][12][1] = (sum_out[13][12][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][12][1] = (sum_out[14][12][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][12][1] = (sum_out[15][12][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][12][1] = (sum_out[16][12][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][12][1] = (sum_out[17][12][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][12][1] = (sum_out[18][12][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][12][1] = (sum_out[19][12][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][12][2] = (sum_out[0][12][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][12][2] = (sum_out[1][12][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][12][2] = (sum_out[2][12][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][12][2] = (sum_out[3][12][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][12][2] = (sum_out[4][12][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][12][2] = (sum_out[5][12][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][12][2] = (sum_out[6][12][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][12][2] = (sum_out[7][12][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][12][2] = (sum_out[8][12][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][12][2] = (sum_out[9][12][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][12][2] = (sum_out[10][12][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][12][2] = (sum_out[11][12][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][12][2] = (sum_out[12][12][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][12][2] = (sum_out[13][12][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][12][2] = (sum_out[14][12][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][12][2] = (sum_out[15][12][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][12][2] = (sum_out[16][12][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][12][2] = (sum_out[17][12][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][12][2] = (sum_out[18][12][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][12][2] = (sum_out[19][12][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][12][3] = (sum_out[0][12][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][12][3] = (sum_out[1][12][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][12][3] = (sum_out[2][12][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][12][3] = (sum_out[3][12][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][12][3] = (sum_out[4][12][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][12][3] = (sum_out[5][12][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][12][3] = (sum_out[6][12][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][12][3] = (sum_out[7][12][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][12][3] = (sum_out[8][12][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][12][3] = (sum_out[9][12][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][12][3] = (sum_out[10][12][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][12][3] = (sum_out[11][12][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][12][3] = (sum_out[12][12][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][12][3] = (sum_out[13][12][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][12][3] = (sum_out[14][12][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][12][3] = (sum_out[15][12][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][12][3] = (sum_out[16][12][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][12][3] = (sum_out[17][12][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][12][3] = (sum_out[18][12][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][12][3] = (sum_out[19][12][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][12][4] = (sum_out[0][12][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][12][4] = (sum_out[1][12][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][12][4] = (sum_out[2][12][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][12][4] = (sum_out[3][12][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][12][4] = (sum_out[4][12][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][12][4] = (sum_out[5][12][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][12][4] = (sum_out[6][12][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][12][4] = (sum_out[7][12][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][12][4] = (sum_out[8][12][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][12][4] = (sum_out[9][12][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][12][4] = (sum_out[10][12][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][12][4] = (sum_out[11][12][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][12][4] = (sum_out[12][12][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][12][4] = (sum_out[13][12][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][12][4] = (sum_out[14][12][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][12][4] = (sum_out[15][12][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][12][4] = (sum_out[16][12][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][12][4] = (sum_out[17][12][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][12][4] = (sum_out[18][12][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][12][4] = (sum_out[19][12][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][12][5] = (sum_out[0][12][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][12][5] = (sum_out[1][12][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][12][5] = (sum_out[2][12][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][12][5] = (sum_out[3][12][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][12][5] = (sum_out[4][12][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][12][5] = (sum_out[5][12][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][12][5] = (sum_out[6][12][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][12][5] = (sum_out[7][12][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][12][5] = (sum_out[8][12][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][12][5] = (sum_out[9][12][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][12][5] = (sum_out[10][12][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][12][5] = (sum_out[11][12][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][12][5] = (sum_out[12][12][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][12][5] = (sum_out[13][12][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][12][5] = (sum_out[14][12][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][12][5] = (sum_out[15][12][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][12][5] = (sum_out[16][12][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][12][5] = (sum_out[17][12][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][12][5] = (sum_out[18][12][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][12][5] = (sum_out[19][12][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][12][6] = (sum_out[0][12][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][12][6] = (sum_out[1][12][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][12][6] = (sum_out[2][12][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][12][6] = (sum_out[3][12][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][12][6] = (sum_out[4][12][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][12][6] = (sum_out[5][12][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][12][6] = (sum_out[6][12][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][12][6] = (sum_out[7][12][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][12][6] = (sum_out[8][12][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][12][6] = (sum_out[9][12][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][12][6] = (sum_out[10][12][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][12][6] = (sum_out[11][12][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][12][6] = (sum_out[12][12][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][12][6] = (sum_out[13][12][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][12][6] = (sum_out[14][12][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][12][6] = (sum_out[15][12][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][12][6] = (sum_out[16][12][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][12][6] = (sum_out[17][12][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][12][6] = (sum_out[18][12][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][12][6] = (sum_out[19][12][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][12][7] = (sum_out[0][12][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][12][7] = (sum_out[1][12][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][12][7] = (sum_out[2][12][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][12][7] = (sum_out[3][12][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][12][7] = (sum_out[4][12][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][12][7] = (sum_out[5][12][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][12][7] = (sum_out[6][12][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][12][7] = (sum_out[7][12][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][12][7] = (sum_out[8][12][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][12][7] = (sum_out[9][12][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][12][7] = (sum_out[10][12][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][12][7] = (sum_out[11][12][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][12][7] = (sum_out[12][12][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][12][7] = (sum_out[13][12][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][12][7] = (sum_out[14][12][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][12][7] = (sum_out[15][12][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][12][7] = (sum_out[16][12][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][12][7] = (sum_out[17][12][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][12][7] = (sum_out[18][12][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][12][7] = (sum_out[19][12][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][12][8] = (sum_out[0][12][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][12][8] = (sum_out[1][12][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][12][8] = (sum_out[2][12][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][12][8] = (sum_out[3][12][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][12][8] = (sum_out[4][12][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][12][8] = (sum_out[5][12][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][12][8] = (sum_out[6][12][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][12][8] = (sum_out[7][12][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][12][8] = (sum_out[8][12][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][12][8] = (sum_out[9][12][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][12][8] = (sum_out[10][12][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][12][8] = (sum_out[11][12][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][12][8] = (sum_out[12][12][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][12][8] = (sum_out[13][12][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][12][8] = (sum_out[14][12][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][12][8] = (sum_out[15][12][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][12][8] = (sum_out[16][12][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][12][8] = (sum_out[17][12][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][12][8] = (sum_out[18][12][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][12][8] = (sum_out[19][12][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][12][9] = (sum_out[0][12][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][12][9] = (sum_out[1][12][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][12][9] = (sum_out[2][12][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][12][9] = (sum_out[3][12][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][12][9] = (sum_out[4][12][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][12][9] = (sum_out[5][12][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][12][9] = (sum_out[6][12][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][12][9] = (sum_out[7][12][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][12][9] = (sum_out[8][12][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][12][9] = (sum_out[9][12][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][12][9] = (sum_out[10][12][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][12][9] = (sum_out[11][12][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][12][9] = (sum_out[12][12][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][12][9] = (sum_out[13][12][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][12][9] = (sum_out[14][12][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][12][9] = (sum_out[15][12][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][12][9] = (sum_out[16][12][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][12][9] = (sum_out[17][12][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][12][9] = (sum_out[18][12][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][12][9] = (sum_out[19][12][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][12][10] = (sum_out[0][12][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][12][10] = (sum_out[1][12][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][12][10] = (sum_out[2][12][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][12][10] = (sum_out[3][12][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][12][10] = (sum_out[4][12][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][12][10] = (sum_out[5][12][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][12][10] = (sum_out[6][12][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][12][10] = (sum_out[7][12][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][12][10] = (sum_out[8][12][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][12][10] = (sum_out[9][12][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][12][10] = (sum_out[10][12][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][12][10] = (sum_out[11][12][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][12][10] = (sum_out[12][12][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][12][10] = (sum_out[13][12][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][12][10] = (sum_out[14][12][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][12][10] = (sum_out[15][12][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][12][10] = (sum_out[16][12][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][12][10] = (sum_out[17][12][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][12][10] = (sum_out[18][12][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][12][10] = (sum_out[19][12][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][12][11] = (sum_out[0][12][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][12][11] = (sum_out[1][12][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][12][11] = (sum_out[2][12][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][12][11] = (sum_out[3][12][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][12][11] = (sum_out[4][12][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][12][11] = (sum_out[5][12][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][12][11] = (sum_out[6][12][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][12][11] = (sum_out[7][12][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][12][11] = (sum_out[8][12][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][12][11] = (sum_out[9][12][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][12][11] = (sum_out[10][12][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][12][11] = (sum_out[11][12][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][12][11] = (sum_out[12][12][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][12][11] = (sum_out[13][12][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][12][11] = (sum_out[14][12][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][12][11] = (sum_out[15][12][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][12][11] = (sum_out[16][12][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][12][11] = (sum_out[17][12][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][12][11] = (sum_out[18][12][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][12][11] = (sum_out[19][12][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][12][12] = (sum_out[0][12][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][12][12] = (sum_out[1][12][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][12][12] = (sum_out[2][12][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][12][12] = (sum_out[3][12][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][12][12] = (sum_out[4][12][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][12][12] = (sum_out[5][12][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][12][12] = (sum_out[6][12][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][12][12] = (sum_out[7][12][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][12][12] = (sum_out[8][12][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][12][12] = (sum_out[9][12][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][12][12] = (sum_out[10][12][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][12][12] = (sum_out[11][12][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][12][12] = (sum_out[12][12][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][12][12] = (sum_out[13][12][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][12][12] = (sum_out[14][12][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][12][12] = (sum_out[15][12][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][12][12] = (sum_out[16][12][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][12][12] = (sum_out[17][12][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][12][12] = (sum_out[18][12][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][12][12] = (sum_out[19][12][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][12][13] = (sum_out[0][12][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][12][13] = (sum_out[1][12][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][12][13] = (sum_out[2][12][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][12][13] = (sum_out[3][12][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][12][13] = (sum_out[4][12][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][12][13] = (sum_out[5][12][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][12][13] = (sum_out[6][12][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][12][13] = (sum_out[7][12][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][12][13] = (sum_out[8][12][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][12][13] = (sum_out[9][12][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][12][13] = (sum_out[10][12][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][12][13] = (sum_out[11][12][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][12][13] = (sum_out[12][12][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][12][13] = (sum_out[13][12][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][12][13] = (sum_out[14][12][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][12][13] = (sum_out[15][12][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][12][13] = (sum_out[16][12][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][12][13] = (sum_out[17][12][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][12][13] = (sum_out[18][12][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][12][13] = (sum_out[19][12][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][12][14] = (sum_out[0][12][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][12][14] = (sum_out[1][12][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][12][14] = (sum_out[2][12][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][12][14] = (sum_out[3][12][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][12][14] = (sum_out[4][12][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][12][14] = (sum_out[5][12][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][12][14] = (sum_out[6][12][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][12][14] = (sum_out[7][12][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][12][14] = (sum_out[8][12][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][12][14] = (sum_out[9][12][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][12][14] = (sum_out[10][12][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][12][14] = (sum_out[11][12][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][12][14] = (sum_out[12][12][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][12][14] = (sum_out[13][12][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][12][14] = (sum_out[14][12][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][12][14] = (sum_out[15][12][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][12][14] = (sum_out[16][12][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][12][14] = (sum_out[17][12][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][12][14] = (sum_out[18][12][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][12][14] = (sum_out[19][12][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][12][15] = (sum_out[0][12][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][12][15] = (sum_out[1][12][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][12][15] = (sum_out[2][12][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][12][15] = (sum_out[3][12][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][12][15] = (sum_out[4][12][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][12][15] = (sum_out[5][12][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][12][15] = (sum_out[6][12][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][12][15] = (sum_out[7][12][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][12][15] = (sum_out[8][12][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][12][15] = (sum_out[9][12][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][12][15] = (sum_out[10][12][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][12][15] = (sum_out[11][12][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][12][15] = (sum_out[12][12][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][12][15] = (sum_out[13][12][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][12][15] = (sum_out[14][12][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][12][15] = (sum_out[15][12][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][12][15] = (sum_out[16][12][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][12][15] = (sum_out[17][12][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][12][15] = (sum_out[18][12][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][12][15] = (sum_out[19][12][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][12][16] = (sum_out[0][12][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][12][16] = (sum_out[1][12][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][12][16] = (sum_out[2][12][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][12][16] = (sum_out[3][12][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][12][16] = (sum_out[4][12][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][12][16] = (sum_out[5][12][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][12][16] = (sum_out[6][12][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][12][16] = (sum_out[7][12][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][12][16] = (sum_out[8][12][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][12][16] = (sum_out[9][12][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][12][16] = (sum_out[10][12][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][12][16] = (sum_out[11][12][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][12][16] = (sum_out[12][12][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][12][16] = (sum_out[13][12][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][12][16] = (sum_out[14][12][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][12][16] = (sum_out[15][12][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][12][16] = (sum_out[16][12][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][12][16] = (sum_out[17][12][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][12][16] = (sum_out[18][12][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][12][16] = (sum_out[19][12][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][12][17] = (sum_out[0][12][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][12][17] = (sum_out[1][12][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][12][17] = (sum_out[2][12][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][12][17] = (sum_out[3][12][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][12][17] = (sum_out[4][12][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][12][17] = (sum_out[5][12][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][12][17] = (sum_out[6][12][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][12][17] = (sum_out[7][12][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][12][17] = (sum_out[8][12][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][12][17] = (sum_out[9][12][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][12][17] = (sum_out[10][12][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][12][17] = (sum_out[11][12][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][12][17] = (sum_out[12][12][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][12][17] = (sum_out[13][12][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][12][17] = (sum_out[14][12][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][12][17] = (sum_out[15][12][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][12][17] = (sum_out[16][12][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][12][17] = (sum_out[17][12][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][12][17] = (sum_out[18][12][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][12][17] = (sum_out[19][12][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][12][18] = (sum_out[0][12][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][12][18] = (sum_out[1][12][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][12][18] = (sum_out[2][12][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][12][18] = (sum_out[3][12][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][12][18] = (sum_out[4][12][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][12][18] = (sum_out[5][12][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][12][18] = (sum_out[6][12][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][12][18] = (sum_out[7][12][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][12][18] = (sum_out[8][12][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][12][18] = (sum_out[9][12][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][12][18] = (sum_out[10][12][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][12][18] = (sum_out[11][12][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][12][18] = (sum_out[12][12][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][12][18] = (sum_out[13][12][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][12][18] = (sum_out[14][12][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][12][18] = (sum_out[15][12][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][12][18] = (sum_out[16][12][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][12][18] = (sum_out[17][12][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][12][18] = (sum_out[18][12][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][12][18] = (sum_out[19][12][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][12][19] = (sum_out[0][12][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][12][19] = (sum_out[1][12][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][12][19] = (sum_out[2][12][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][12][19] = (sum_out[3][12][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][12][19] = (sum_out[4][12][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][12][19] = (sum_out[5][12][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][12][19] = (sum_out[6][12][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][12][19] = (sum_out[7][12][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][12][19] = (sum_out[8][12][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][12][19] = (sum_out[9][12][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][12][19] = (sum_out[10][12][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][12][19] = (sum_out[11][12][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][12][19] = (sum_out[12][12][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][12][19] = (sum_out[13][12][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][12][19] = (sum_out[14][12][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][12][19] = (sum_out[15][12][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][12][19] = (sum_out[16][12][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][12][19] = (sum_out[17][12][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][12][19] = (sum_out[18][12][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][12][19] = (sum_out[19][12][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][12][20] = (sum_out[0][12][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][12][20] = (sum_out[1][12][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][12][20] = (sum_out[2][12][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][12][20] = (sum_out[3][12][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][12][20] = (sum_out[4][12][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][12][20] = (sum_out[5][12][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][12][20] = (sum_out[6][12][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][12][20] = (sum_out[7][12][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][12][20] = (sum_out[8][12][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][12][20] = (sum_out[9][12][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][12][20] = (sum_out[10][12][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][12][20] = (sum_out[11][12][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][12][20] = (sum_out[12][12][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][12][20] = (sum_out[13][12][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][12][20] = (sum_out[14][12][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][12][20] = (sum_out[15][12][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][12][20] = (sum_out[16][12][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][12][20] = (sum_out[17][12][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][12][20] = (sum_out[18][12][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][12][20] = (sum_out[19][12][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][12][21] = (sum_out[0][12][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][12][21] = (sum_out[1][12][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][12][21] = (sum_out[2][12][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][12][21] = (sum_out[3][12][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][12][21] = (sum_out[4][12][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][12][21] = (sum_out[5][12][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][12][21] = (sum_out[6][12][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][12][21] = (sum_out[7][12][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][12][21] = (sum_out[8][12][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][12][21] = (sum_out[9][12][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][12][21] = (sum_out[10][12][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][12][21] = (sum_out[11][12][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][12][21] = (sum_out[12][12][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][12][21] = (sum_out[13][12][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][12][21] = (sum_out[14][12][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][12][21] = (sum_out[15][12][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][12][21] = (sum_out[16][12][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][12][21] = (sum_out[17][12][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][12][21] = (sum_out[18][12][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][12][21] = (sum_out[19][12][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][12][22] = (sum_out[0][12][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][12][22] = (sum_out[1][12][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][12][22] = (sum_out[2][12][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][12][22] = (sum_out[3][12][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][12][22] = (sum_out[4][12][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][12][22] = (sum_out[5][12][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][12][22] = (sum_out[6][12][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][12][22] = (sum_out[7][12][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][12][22] = (sum_out[8][12][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][12][22] = (sum_out[9][12][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][12][22] = (sum_out[10][12][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][12][22] = (sum_out[11][12][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][12][22] = (sum_out[12][12][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][12][22] = (sum_out[13][12][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][12][22] = (sum_out[14][12][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][12][22] = (sum_out[15][12][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][12][22] = (sum_out[16][12][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][12][22] = (sum_out[17][12][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][12][22] = (sum_out[18][12][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][12][22] = (sum_out[19][12][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][12][23] = (sum_out[0][12][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][12][23] = (sum_out[1][12][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][12][23] = (sum_out[2][12][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][12][23] = (sum_out[3][12][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][12][23] = (sum_out[4][12][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][12][23] = (sum_out[5][12][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][12][23] = (sum_out[6][12][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][12][23] = (sum_out[7][12][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][12][23] = (sum_out[8][12][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][12][23] = (sum_out[9][12][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][12][23] = (sum_out[10][12][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][12][23] = (sum_out[11][12][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][12][23] = (sum_out[12][12][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][12][23] = (sum_out[13][12][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][12][23] = (sum_out[14][12][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][12][23] = (sum_out[15][12][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][12][23] = (sum_out[16][12][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][12][23] = (sum_out[17][12][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][12][23] = (sum_out[18][12][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][12][23] = (sum_out[19][12][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][13][0] = (sum_out[0][13][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][13][0] = (sum_out[1][13][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][13][0] = (sum_out[2][13][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][13][0] = (sum_out[3][13][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][13][0] = (sum_out[4][13][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][13][0] = (sum_out[5][13][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][13][0] = (sum_out[6][13][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][13][0] = (sum_out[7][13][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][13][0] = (sum_out[8][13][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][13][0] = (sum_out[9][13][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][13][0] = (sum_out[10][13][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][13][0] = (sum_out[11][13][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][13][0] = (sum_out[12][13][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][13][0] = (sum_out[13][13][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][13][0] = (sum_out[14][13][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][13][0] = (sum_out[15][13][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][13][0] = (sum_out[16][13][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][13][0] = (sum_out[17][13][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][13][0] = (sum_out[18][13][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][13][0] = (sum_out[19][13][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][13][1] = (sum_out[0][13][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][13][1] = (sum_out[1][13][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][13][1] = (sum_out[2][13][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][13][1] = (sum_out[3][13][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][13][1] = (sum_out[4][13][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][13][1] = (sum_out[5][13][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][13][1] = (sum_out[6][13][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][13][1] = (sum_out[7][13][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][13][1] = (sum_out[8][13][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][13][1] = (sum_out[9][13][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][13][1] = (sum_out[10][13][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][13][1] = (sum_out[11][13][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][13][1] = (sum_out[12][13][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][13][1] = (sum_out[13][13][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][13][1] = (sum_out[14][13][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][13][1] = (sum_out[15][13][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][13][1] = (sum_out[16][13][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][13][1] = (sum_out[17][13][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][13][1] = (sum_out[18][13][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][13][1] = (sum_out[19][13][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][13][2] = (sum_out[0][13][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][13][2] = (sum_out[1][13][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][13][2] = (sum_out[2][13][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][13][2] = (sum_out[3][13][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][13][2] = (sum_out[4][13][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][13][2] = (sum_out[5][13][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][13][2] = (sum_out[6][13][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][13][2] = (sum_out[7][13][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][13][2] = (sum_out[8][13][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][13][2] = (sum_out[9][13][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][13][2] = (sum_out[10][13][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][13][2] = (sum_out[11][13][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][13][2] = (sum_out[12][13][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][13][2] = (sum_out[13][13][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][13][2] = (sum_out[14][13][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][13][2] = (sum_out[15][13][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][13][2] = (sum_out[16][13][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][13][2] = (sum_out[17][13][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][13][2] = (sum_out[18][13][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][13][2] = (sum_out[19][13][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][13][3] = (sum_out[0][13][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][13][3] = (sum_out[1][13][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][13][3] = (sum_out[2][13][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][13][3] = (sum_out[3][13][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][13][3] = (sum_out[4][13][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][13][3] = (sum_out[5][13][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][13][3] = (sum_out[6][13][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][13][3] = (sum_out[7][13][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][13][3] = (sum_out[8][13][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][13][3] = (sum_out[9][13][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][13][3] = (sum_out[10][13][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][13][3] = (sum_out[11][13][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][13][3] = (sum_out[12][13][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][13][3] = (sum_out[13][13][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][13][3] = (sum_out[14][13][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][13][3] = (sum_out[15][13][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][13][3] = (sum_out[16][13][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][13][3] = (sum_out[17][13][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][13][3] = (sum_out[18][13][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][13][3] = (sum_out[19][13][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][13][4] = (sum_out[0][13][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][13][4] = (sum_out[1][13][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][13][4] = (sum_out[2][13][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][13][4] = (sum_out[3][13][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][13][4] = (sum_out[4][13][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][13][4] = (sum_out[5][13][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][13][4] = (sum_out[6][13][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][13][4] = (sum_out[7][13][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][13][4] = (sum_out[8][13][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][13][4] = (sum_out[9][13][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][13][4] = (sum_out[10][13][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][13][4] = (sum_out[11][13][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][13][4] = (sum_out[12][13][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][13][4] = (sum_out[13][13][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][13][4] = (sum_out[14][13][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][13][4] = (sum_out[15][13][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][13][4] = (sum_out[16][13][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][13][4] = (sum_out[17][13][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][13][4] = (sum_out[18][13][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][13][4] = (sum_out[19][13][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][13][5] = (sum_out[0][13][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][13][5] = (sum_out[1][13][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][13][5] = (sum_out[2][13][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][13][5] = (sum_out[3][13][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][13][5] = (sum_out[4][13][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][13][5] = (sum_out[5][13][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][13][5] = (sum_out[6][13][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][13][5] = (sum_out[7][13][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][13][5] = (sum_out[8][13][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][13][5] = (sum_out[9][13][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][13][5] = (sum_out[10][13][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][13][5] = (sum_out[11][13][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][13][5] = (sum_out[12][13][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][13][5] = (sum_out[13][13][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][13][5] = (sum_out[14][13][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][13][5] = (sum_out[15][13][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][13][5] = (sum_out[16][13][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][13][5] = (sum_out[17][13][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][13][5] = (sum_out[18][13][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][13][5] = (sum_out[19][13][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][13][6] = (sum_out[0][13][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][13][6] = (sum_out[1][13][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][13][6] = (sum_out[2][13][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][13][6] = (sum_out[3][13][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][13][6] = (sum_out[4][13][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][13][6] = (sum_out[5][13][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][13][6] = (sum_out[6][13][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][13][6] = (sum_out[7][13][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][13][6] = (sum_out[8][13][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][13][6] = (sum_out[9][13][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][13][6] = (sum_out[10][13][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][13][6] = (sum_out[11][13][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][13][6] = (sum_out[12][13][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][13][6] = (sum_out[13][13][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][13][6] = (sum_out[14][13][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][13][6] = (sum_out[15][13][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][13][6] = (sum_out[16][13][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][13][6] = (sum_out[17][13][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][13][6] = (sum_out[18][13][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][13][6] = (sum_out[19][13][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][13][7] = (sum_out[0][13][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][13][7] = (sum_out[1][13][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][13][7] = (sum_out[2][13][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][13][7] = (sum_out[3][13][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][13][7] = (sum_out[4][13][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][13][7] = (sum_out[5][13][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][13][7] = (sum_out[6][13][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][13][7] = (sum_out[7][13][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][13][7] = (sum_out[8][13][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][13][7] = (sum_out[9][13][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][13][7] = (sum_out[10][13][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][13][7] = (sum_out[11][13][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][13][7] = (sum_out[12][13][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][13][7] = (sum_out[13][13][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][13][7] = (sum_out[14][13][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][13][7] = (sum_out[15][13][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][13][7] = (sum_out[16][13][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][13][7] = (sum_out[17][13][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][13][7] = (sum_out[18][13][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][13][7] = (sum_out[19][13][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][13][8] = (sum_out[0][13][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][13][8] = (sum_out[1][13][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][13][8] = (sum_out[2][13][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][13][8] = (sum_out[3][13][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][13][8] = (sum_out[4][13][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][13][8] = (sum_out[5][13][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][13][8] = (sum_out[6][13][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][13][8] = (sum_out[7][13][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][13][8] = (sum_out[8][13][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][13][8] = (sum_out[9][13][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][13][8] = (sum_out[10][13][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][13][8] = (sum_out[11][13][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][13][8] = (sum_out[12][13][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][13][8] = (sum_out[13][13][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][13][8] = (sum_out[14][13][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][13][8] = (sum_out[15][13][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][13][8] = (sum_out[16][13][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][13][8] = (sum_out[17][13][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][13][8] = (sum_out[18][13][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][13][8] = (sum_out[19][13][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][13][9] = (sum_out[0][13][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][13][9] = (sum_out[1][13][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][13][9] = (sum_out[2][13][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][13][9] = (sum_out[3][13][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][13][9] = (sum_out[4][13][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][13][9] = (sum_out[5][13][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][13][9] = (sum_out[6][13][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][13][9] = (sum_out[7][13][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][13][9] = (sum_out[8][13][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][13][9] = (sum_out[9][13][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][13][9] = (sum_out[10][13][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][13][9] = (sum_out[11][13][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][13][9] = (sum_out[12][13][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][13][9] = (sum_out[13][13][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][13][9] = (sum_out[14][13][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][13][9] = (sum_out[15][13][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][13][9] = (sum_out[16][13][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][13][9] = (sum_out[17][13][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][13][9] = (sum_out[18][13][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][13][9] = (sum_out[19][13][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][13][10] = (sum_out[0][13][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][13][10] = (sum_out[1][13][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][13][10] = (sum_out[2][13][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][13][10] = (sum_out[3][13][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][13][10] = (sum_out[4][13][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][13][10] = (sum_out[5][13][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][13][10] = (sum_out[6][13][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][13][10] = (sum_out[7][13][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][13][10] = (sum_out[8][13][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][13][10] = (sum_out[9][13][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][13][10] = (sum_out[10][13][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][13][10] = (sum_out[11][13][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][13][10] = (sum_out[12][13][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][13][10] = (sum_out[13][13][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][13][10] = (sum_out[14][13][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][13][10] = (sum_out[15][13][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][13][10] = (sum_out[16][13][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][13][10] = (sum_out[17][13][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][13][10] = (sum_out[18][13][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][13][10] = (sum_out[19][13][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][13][11] = (sum_out[0][13][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][13][11] = (sum_out[1][13][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][13][11] = (sum_out[2][13][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][13][11] = (sum_out[3][13][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][13][11] = (sum_out[4][13][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][13][11] = (sum_out[5][13][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][13][11] = (sum_out[6][13][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][13][11] = (sum_out[7][13][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][13][11] = (sum_out[8][13][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][13][11] = (sum_out[9][13][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][13][11] = (sum_out[10][13][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][13][11] = (sum_out[11][13][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][13][11] = (sum_out[12][13][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][13][11] = (sum_out[13][13][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][13][11] = (sum_out[14][13][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][13][11] = (sum_out[15][13][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][13][11] = (sum_out[16][13][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][13][11] = (sum_out[17][13][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][13][11] = (sum_out[18][13][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][13][11] = (sum_out[19][13][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][13][12] = (sum_out[0][13][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][13][12] = (sum_out[1][13][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][13][12] = (sum_out[2][13][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][13][12] = (sum_out[3][13][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][13][12] = (sum_out[4][13][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][13][12] = (sum_out[5][13][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][13][12] = (sum_out[6][13][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][13][12] = (sum_out[7][13][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][13][12] = (sum_out[8][13][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][13][12] = (sum_out[9][13][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][13][12] = (sum_out[10][13][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][13][12] = (sum_out[11][13][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][13][12] = (sum_out[12][13][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][13][12] = (sum_out[13][13][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][13][12] = (sum_out[14][13][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][13][12] = (sum_out[15][13][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][13][12] = (sum_out[16][13][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][13][12] = (sum_out[17][13][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][13][12] = (sum_out[18][13][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][13][12] = (sum_out[19][13][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][13][13] = (sum_out[0][13][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][13][13] = (sum_out[1][13][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][13][13] = (sum_out[2][13][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][13][13] = (sum_out[3][13][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][13][13] = (sum_out[4][13][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][13][13] = (sum_out[5][13][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][13][13] = (sum_out[6][13][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][13][13] = (sum_out[7][13][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][13][13] = (sum_out[8][13][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][13][13] = (sum_out[9][13][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][13][13] = (sum_out[10][13][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][13][13] = (sum_out[11][13][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][13][13] = (sum_out[12][13][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][13][13] = (sum_out[13][13][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][13][13] = (sum_out[14][13][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][13][13] = (sum_out[15][13][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][13][13] = (sum_out[16][13][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][13][13] = (sum_out[17][13][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][13][13] = (sum_out[18][13][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][13][13] = (sum_out[19][13][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][13][14] = (sum_out[0][13][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][13][14] = (sum_out[1][13][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][13][14] = (sum_out[2][13][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][13][14] = (sum_out[3][13][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][13][14] = (sum_out[4][13][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][13][14] = (sum_out[5][13][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][13][14] = (sum_out[6][13][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][13][14] = (sum_out[7][13][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][13][14] = (sum_out[8][13][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][13][14] = (sum_out[9][13][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][13][14] = (sum_out[10][13][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][13][14] = (sum_out[11][13][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][13][14] = (sum_out[12][13][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][13][14] = (sum_out[13][13][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][13][14] = (sum_out[14][13][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][13][14] = (sum_out[15][13][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][13][14] = (sum_out[16][13][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][13][14] = (sum_out[17][13][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][13][14] = (sum_out[18][13][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][13][14] = (sum_out[19][13][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][13][15] = (sum_out[0][13][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][13][15] = (sum_out[1][13][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][13][15] = (sum_out[2][13][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][13][15] = (sum_out[3][13][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][13][15] = (sum_out[4][13][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][13][15] = (sum_out[5][13][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][13][15] = (sum_out[6][13][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][13][15] = (sum_out[7][13][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][13][15] = (sum_out[8][13][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][13][15] = (sum_out[9][13][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][13][15] = (sum_out[10][13][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][13][15] = (sum_out[11][13][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][13][15] = (sum_out[12][13][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][13][15] = (sum_out[13][13][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][13][15] = (sum_out[14][13][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][13][15] = (sum_out[15][13][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][13][15] = (sum_out[16][13][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][13][15] = (sum_out[17][13][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][13][15] = (sum_out[18][13][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][13][15] = (sum_out[19][13][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][13][16] = (sum_out[0][13][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][13][16] = (sum_out[1][13][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][13][16] = (sum_out[2][13][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][13][16] = (sum_out[3][13][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][13][16] = (sum_out[4][13][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][13][16] = (sum_out[5][13][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][13][16] = (sum_out[6][13][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][13][16] = (sum_out[7][13][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][13][16] = (sum_out[8][13][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][13][16] = (sum_out[9][13][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][13][16] = (sum_out[10][13][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][13][16] = (sum_out[11][13][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][13][16] = (sum_out[12][13][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][13][16] = (sum_out[13][13][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][13][16] = (sum_out[14][13][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][13][16] = (sum_out[15][13][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][13][16] = (sum_out[16][13][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][13][16] = (sum_out[17][13][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][13][16] = (sum_out[18][13][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][13][16] = (sum_out[19][13][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][13][17] = (sum_out[0][13][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][13][17] = (sum_out[1][13][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][13][17] = (sum_out[2][13][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][13][17] = (sum_out[3][13][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][13][17] = (sum_out[4][13][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][13][17] = (sum_out[5][13][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][13][17] = (sum_out[6][13][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][13][17] = (sum_out[7][13][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][13][17] = (sum_out[8][13][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][13][17] = (sum_out[9][13][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][13][17] = (sum_out[10][13][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][13][17] = (sum_out[11][13][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][13][17] = (sum_out[12][13][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][13][17] = (sum_out[13][13][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][13][17] = (sum_out[14][13][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][13][17] = (sum_out[15][13][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][13][17] = (sum_out[16][13][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][13][17] = (sum_out[17][13][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][13][17] = (sum_out[18][13][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][13][17] = (sum_out[19][13][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][13][18] = (sum_out[0][13][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][13][18] = (sum_out[1][13][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][13][18] = (sum_out[2][13][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][13][18] = (sum_out[3][13][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][13][18] = (sum_out[4][13][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][13][18] = (sum_out[5][13][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][13][18] = (sum_out[6][13][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][13][18] = (sum_out[7][13][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][13][18] = (sum_out[8][13][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][13][18] = (sum_out[9][13][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][13][18] = (sum_out[10][13][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][13][18] = (sum_out[11][13][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][13][18] = (sum_out[12][13][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][13][18] = (sum_out[13][13][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][13][18] = (sum_out[14][13][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][13][18] = (sum_out[15][13][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][13][18] = (sum_out[16][13][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][13][18] = (sum_out[17][13][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][13][18] = (sum_out[18][13][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][13][18] = (sum_out[19][13][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][13][19] = (sum_out[0][13][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][13][19] = (sum_out[1][13][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][13][19] = (sum_out[2][13][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][13][19] = (sum_out[3][13][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][13][19] = (sum_out[4][13][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][13][19] = (sum_out[5][13][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][13][19] = (sum_out[6][13][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][13][19] = (sum_out[7][13][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][13][19] = (sum_out[8][13][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][13][19] = (sum_out[9][13][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][13][19] = (sum_out[10][13][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][13][19] = (sum_out[11][13][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][13][19] = (sum_out[12][13][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][13][19] = (sum_out[13][13][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][13][19] = (sum_out[14][13][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][13][19] = (sum_out[15][13][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][13][19] = (sum_out[16][13][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][13][19] = (sum_out[17][13][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][13][19] = (sum_out[18][13][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][13][19] = (sum_out[19][13][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][13][20] = (sum_out[0][13][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][13][20] = (sum_out[1][13][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][13][20] = (sum_out[2][13][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][13][20] = (sum_out[3][13][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][13][20] = (sum_out[4][13][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][13][20] = (sum_out[5][13][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][13][20] = (sum_out[6][13][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][13][20] = (sum_out[7][13][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][13][20] = (sum_out[8][13][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][13][20] = (sum_out[9][13][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][13][20] = (sum_out[10][13][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][13][20] = (sum_out[11][13][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][13][20] = (sum_out[12][13][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][13][20] = (sum_out[13][13][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][13][20] = (sum_out[14][13][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][13][20] = (sum_out[15][13][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][13][20] = (sum_out[16][13][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][13][20] = (sum_out[17][13][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][13][20] = (sum_out[18][13][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][13][20] = (sum_out[19][13][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][13][21] = (sum_out[0][13][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][13][21] = (sum_out[1][13][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][13][21] = (sum_out[2][13][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][13][21] = (sum_out[3][13][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][13][21] = (sum_out[4][13][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][13][21] = (sum_out[5][13][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][13][21] = (sum_out[6][13][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][13][21] = (sum_out[7][13][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][13][21] = (sum_out[8][13][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][13][21] = (sum_out[9][13][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][13][21] = (sum_out[10][13][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][13][21] = (sum_out[11][13][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][13][21] = (sum_out[12][13][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][13][21] = (sum_out[13][13][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][13][21] = (sum_out[14][13][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][13][21] = (sum_out[15][13][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][13][21] = (sum_out[16][13][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][13][21] = (sum_out[17][13][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][13][21] = (sum_out[18][13][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][13][21] = (sum_out[19][13][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][13][22] = (sum_out[0][13][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][13][22] = (sum_out[1][13][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][13][22] = (sum_out[2][13][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][13][22] = (sum_out[3][13][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][13][22] = (sum_out[4][13][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][13][22] = (sum_out[5][13][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][13][22] = (sum_out[6][13][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][13][22] = (sum_out[7][13][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][13][22] = (sum_out[8][13][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][13][22] = (sum_out[9][13][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][13][22] = (sum_out[10][13][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][13][22] = (sum_out[11][13][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][13][22] = (sum_out[12][13][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][13][22] = (sum_out[13][13][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][13][22] = (sum_out[14][13][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][13][22] = (sum_out[15][13][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][13][22] = (sum_out[16][13][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][13][22] = (sum_out[17][13][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][13][22] = (sum_out[18][13][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][13][22] = (sum_out[19][13][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][13][23] = (sum_out[0][13][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][13][23] = (sum_out[1][13][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][13][23] = (sum_out[2][13][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][13][23] = (sum_out[3][13][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][13][23] = (sum_out[4][13][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][13][23] = (sum_out[5][13][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][13][23] = (sum_out[6][13][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][13][23] = (sum_out[7][13][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][13][23] = (sum_out[8][13][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][13][23] = (sum_out[9][13][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][13][23] = (sum_out[10][13][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][13][23] = (sum_out[11][13][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][13][23] = (sum_out[12][13][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][13][23] = (sum_out[13][13][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][13][23] = (sum_out[14][13][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][13][23] = (sum_out[15][13][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][13][23] = (sum_out[16][13][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][13][23] = (sum_out[17][13][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][13][23] = (sum_out[18][13][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][13][23] = (sum_out[19][13][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][14][0] = (sum_out[0][14][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][14][0] = (sum_out[1][14][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][14][0] = (sum_out[2][14][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][14][0] = (sum_out[3][14][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][14][0] = (sum_out[4][14][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][14][0] = (sum_out[5][14][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][14][0] = (sum_out[6][14][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][14][0] = (sum_out[7][14][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][14][0] = (sum_out[8][14][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][14][0] = (sum_out[9][14][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][14][0] = (sum_out[10][14][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][14][0] = (sum_out[11][14][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][14][0] = (sum_out[12][14][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][14][0] = (sum_out[13][14][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][14][0] = (sum_out[14][14][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][14][0] = (sum_out[15][14][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][14][0] = (sum_out[16][14][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][14][0] = (sum_out[17][14][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][14][0] = (sum_out[18][14][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][14][0] = (sum_out[19][14][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][14][1] = (sum_out[0][14][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][14][1] = (sum_out[1][14][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][14][1] = (sum_out[2][14][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][14][1] = (sum_out[3][14][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][14][1] = (sum_out[4][14][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][14][1] = (sum_out[5][14][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][14][1] = (sum_out[6][14][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][14][1] = (sum_out[7][14][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][14][1] = (sum_out[8][14][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][14][1] = (sum_out[9][14][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][14][1] = (sum_out[10][14][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][14][1] = (sum_out[11][14][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][14][1] = (sum_out[12][14][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][14][1] = (sum_out[13][14][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][14][1] = (sum_out[14][14][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][14][1] = (sum_out[15][14][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][14][1] = (sum_out[16][14][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][14][1] = (sum_out[17][14][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][14][1] = (sum_out[18][14][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][14][1] = (sum_out[19][14][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][14][2] = (sum_out[0][14][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][14][2] = (sum_out[1][14][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][14][2] = (sum_out[2][14][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][14][2] = (sum_out[3][14][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][14][2] = (sum_out[4][14][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][14][2] = (sum_out[5][14][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][14][2] = (sum_out[6][14][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][14][2] = (sum_out[7][14][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][14][2] = (sum_out[8][14][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][14][2] = (sum_out[9][14][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][14][2] = (sum_out[10][14][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][14][2] = (sum_out[11][14][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][14][2] = (sum_out[12][14][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][14][2] = (sum_out[13][14][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][14][2] = (sum_out[14][14][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][14][2] = (sum_out[15][14][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][14][2] = (sum_out[16][14][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][14][2] = (sum_out[17][14][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][14][2] = (sum_out[18][14][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][14][2] = (sum_out[19][14][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][14][3] = (sum_out[0][14][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][14][3] = (sum_out[1][14][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][14][3] = (sum_out[2][14][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][14][3] = (sum_out[3][14][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][14][3] = (sum_out[4][14][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][14][3] = (sum_out[5][14][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][14][3] = (sum_out[6][14][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][14][3] = (sum_out[7][14][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][14][3] = (sum_out[8][14][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][14][3] = (sum_out[9][14][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][14][3] = (sum_out[10][14][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][14][3] = (sum_out[11][14][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][14][3] = (sum_out[12][14][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][14][3] = (sum_out[13][14][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][14][3] = (sum_out[14][14][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][14][3] = (sum_out[15][14][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][14][3] = (sum_out[16][14][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][14][3] = (sum_out[17][14][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][14][3] = (sum_out[18][14][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][14][3] = (sum_out[19][14][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][14][4] = (sum_out[0][14][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][14][4] = (sum_out[1][14][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][14][4] = (sum_out[2][14][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][14][4] = (sum_out[3][14][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][14][4] = (sum_out[4][14][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][14][4] = (sum_out[5][14][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][14][4] = (sum_out[6][14][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][14][4] = (sum_out[7][14][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][14][4] = (sum_out[8][14][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][14][4] = (sum_out[9][14][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][14][4] = (sum_out[10][14][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][14][4] = (sum_out[11][14][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][14][4] = (sum_out[12][14][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][14][4] = (sum_out[13][14][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][14][4] = (sum_out[14][14][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][14][4] = (sum_out[15][14][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][14][4] = (sum_out[16][14][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][14][4] = (sum_out[17][14][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][14][4] = (sum_out[18][14][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][14][4] = (sum_out[19][14][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][14][5] = (sum_out[0][14][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][14][5] = (sum_out[1][14][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][14][5] = (sum_out[2][14][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][14][5] = (sum_out[3][14][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][14][5] = (sum_out[4][14][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][14][5] = (sum_out[5][14][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][14][5] = (sum_out[6][14][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][14][5] = (sum_out[7][14][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][14][5] = (sum_out[8][14][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][14][5] = (sum_out[9][14][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][14][5] = (sum_out[10][14][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][14][5] = (sum_out[11][14][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][14][5] = (sum_out[12][14][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][14][5] = (sum_out[13][14][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][14][5] = (sum_out[14][14][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][14][5] = (sum_out[15][14][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][14][5] = (sum_out[16][14][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][14][5] = (sum_out[17][14][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][14][5] = (sum_out[18][14][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][14][5] = (sum_out[19][14][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][14][6] = (sum_out[0][14][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][14][6] = (sum_out[1][14][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][14][6] = (sum_out[2][14][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][14][6] = (sum_out[3][14][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][14][6] = (sum_out[4][14][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][14][6] = (sum_out[5][14][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][14][6] = (sum_out[6][14][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][14][6] = (sum_out[7][14][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][14][6] = (sum_out[8][14][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][14][6] = (sum_out[9][14][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][14][6] = (sum_out[10][14][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][14][6] = (sum_out[11][14][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][14][6] = (sum_out[12][14][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][14][6] = (sum_out[13][14][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][14][6] = (sum_out[14][14][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][14][6] = (sum_out[15][14][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][14][6] = (sum_out[16][14][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][14][6] = (sum_out[17][14][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][14][6] = (sum_out[18][14][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][14][6] = (sum_out[19][14][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][14][7] = (sum_out[0][14][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][14][7] = (sum_out[1][14][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][14][7] = (sum_out[2][14][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][14][7] = (sum_out[3][14][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][14][7] = (sum_out[4][14][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][14][7] = (sum_out[5][14][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][14][7] = (sum_out[6][14][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][14][7] = (sum_out[7][14][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][14][7] = (sum_out[8][14][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][14][7] = (sum_out[9][14][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][14][7] = (sum_out[10][14][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][14][7] = (sum_out[11][14][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][14][7] = (sum_out[12][14][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][14][7] = (sum_out[13][14][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][14][7] = (sum_out[14][14][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][14][7] = (sum_out[15][14][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][14][7] = (sum_out[16][14][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][14][7] = (sum_out[17][14][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][14][7] = (sum_out[18][14][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][14][7] = (sum_out[19][14][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][14][8] = (sum_out[0][14][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][14][8] = (sum_out[1][14][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][14][8] = (sum_out[2][14][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][14][8] = (sum_out[3][14][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][14][8] = (sum_out[4][14][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][14][8] = (sum_out[5][14][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][14][8] = (sum_out[6][14][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][14][8] = (sum_out[7][14][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][14][8] = (sum_out[8][14][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][14][8] = (sum_out[9][14][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][14][8] = (sum_out[10][14][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][14][8] = (sum_out[11][14][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][14][8] = (sum_out[12][14][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][14][8] = (sum_out[13][14][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][14][8] = (sum_out[14][14][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][14][8] = (sum_out[15][14][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][14][8] = (sum_out[16][14][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][14][8] = (sum_out[17][14][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][14][8] = (sum_out[18][14][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][14][8] = (sum_out[19][14][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][14][9] = (sum_out[0][14][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][14][9] = (sum_out[1][14][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][14][9] = (sum_out[2][14][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][14][9] = (sum_out[3][14][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][14][9] = (sum_out[4][14][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][14][9] = (sum_out[5][14][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][14][9] = (sum_out[6][14][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][14][9] = (sum_out[7][14][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][14][9] = (sum_out[8][14][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][14][9] = (sum_out[9][14][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][14][9] = (sum_out[10][14][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][14][9] = (sum_out[11][14][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][14][9] = (sum_out[12][14][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][14][9] = (sum_out[13][14][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][14][9] = (sum_out[14][14][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][14][9] = (sum_out[15][14][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][14][9] = (sum_out[16][14][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][14][9] = (sum_out[17][14][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][14][9] = (sum_out[18][14][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][14][9] = (sum_out[19][14][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][14][10] = (sum_out[0][14][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][14][10] = (sum_out[1][14][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][14][10] = (sum_out[2][14][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][14][10] = (sum_out[3][14][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][14][10] = (sum_out[4][14][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][14][10] = (sum_out[5][14][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][14][10] = (sum_out[6][14][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][14][10] = (sum_out[7][14][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][14][10] = (sum_out[8][14][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][14][10] = (sum_out[9][14][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][14][10] = (sum_out[10][14][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][14][10] = (sum_out[11][14][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][14][10] = (sum_out[12][14][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][14][10] = (sum_out[13][14][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][14][10] = (sum_out[14][14][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][14][10] = (sum_out[15][14][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][14][10] = (sum_out[16][14][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][14][10] = (sum_out[17][14][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][14][10] = (sum_out[18][14][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][14][10] = (sum_out[19][14][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][14][11] = (sum_out[0][14][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][14][11] = (sum_out[1][14][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][14][11] = (sum_out[2][14][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][14][11] = (sum_out[3][14][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][14][11] = (sum_out[4][14][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][14][11] = (sum_out[5][14][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][14][11] = (sum_out[6][14][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][14][11] = (sum_out[7][14][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][14][11] = (sum_out[8][14][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][14][11] = (sum_out[9][14][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][14][11] = (sum_out[10][14][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][14][11] = (sum_out[11][14][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][14][11] = (sum_out[12][14][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][14][11] = (sum_out[13][14][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][14][11] = (sum_out[14][14][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][14][11] = (sum_out[15][14][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][14][11] = (sum_out[16][14][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][14][11] = (sum_out[17][14][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][14][11] = (sum_out[18][14][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][14][11] = (sum_out[19][14][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][14][12] = (sum_out[0][14][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][14][12] = (sum_out[1][14][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][14][12] = (sum_out[2][14][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][14][12] = (sum_out[3][14][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][14][12] = (sum_out[4][14][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][14][12] = (sum_out[5][14][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][14][12] = (sum_out[6][14][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][14][12] = (sum_out[7][14][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][14][12] = (sum_out[8][14][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][14][12] = (sum_out[9][14][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][14][12] = (sum_out[10][14][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][14][12] = (sum_out[11][14][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][14][12] = (sum_out[12][14][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][14][12] = (sum_out[13][14][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][14][12] = (sum_out[14][14][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][14][12] = (sum_out[15][14][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][14][12] = (sum_out[16][14][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][14][12] = (sum_out[17][14][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][14][12] = (sum_out[18][14][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][14][12] = (sum_out[19][14][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][14][13] = (sum_out[0][14][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][14][13] = (sum_out[1][14][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][14][13] = (sum_out[2][14][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][14][13] = (sum_out[3][14][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][14][13] = (sum_out[4][14][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][14][13] = (sum_out[5][14][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][14][13] = (sum_out[6][14][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][14][13] = (sum_out[7][14][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][14][13] = (sum_out[8][14][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][14][13] = (sum_out[9][14][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][14][13] = (sum_out[10][14][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][14][13] = (sum_out[11][14][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][14][13] = (sum_out[12][14][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][14][13] = (sum_out[13][14][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][14][13] = (sum_out[14][14][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][14][13] = (sum_out[15][14][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][14][13] = (sum_out[16][14][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][14][13] = (sum_out[17][14][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][14][13] = (sum_out[18][14][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][14][13] = (sum_out[19][14][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][14][14] = (sum_out[0][14][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][14][14] = (sum_out[1][14][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][14][14] = (sum_out[2][14][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][14][14] = (sum_out[3][14][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][14][14] = (sum_out[4][14][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][14][14] = (sum_out[5][14][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][14][14] = (sum_out[6][14][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][14][14] = (sum_out[7][14][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][14][14] = (sum_out[8][14][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][14][14] = (sum_out[9][14][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][14][14] = (sum_out[10][14][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][14][14] = (sum_out[11][14][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][14][14] = (sum_out[12][14][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][14][14] = (sum_out[13][14][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][14][14] = (sum_out[14][14][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][14][14] = (sum_out[15][14][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][14][14] = (sum_out[16][14][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][14][14] = (sum_out[17][14][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][14][14] = (sum_out[18][14][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][14][14] = (sum_out[19][14][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][14][15] = (sum_out[0][14][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][14][15] = (sum_out[1][14][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][14][15] = (sum_out[2][14][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][14][15] = (sum_out[3][14][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][14][15] = (sum_out[4][14][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][14][15] = (sum_out[5][14][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][14][15] = (sum_out[6][14][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][14][15] = (sum_out[7][14][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][14][15] = (sum_out[8][14][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][14][15] = (sum_out[9][14][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][14][15] = (sum_out[10][14][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][14][15] = (sum_out[11][14][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][14][15] = (sum_out[12][14][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][14][15] = (sum_out[13][14][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][14][15] = (sum_out[14][14][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][14][15] = (sum_out[15][14][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][14][15] = (sum_out[16][14][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][14][15] = (sum_out[17][14][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][14][15] = (sum_out[18][14][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][14][15] = (sum_out[19][14][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][14][16] = (sum_out[0][14][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][14][16] = (sum_out[1][14][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][14][16] = (sum_out[2][14][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][14][16] = (sum_out[3][14][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][14][16] = (sum_out[4][14][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][14][16] = (sum_out[5][14][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][14][16] = (sum_out[6][14][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][14][16] = (sum_out[7][14][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][14][16] = (sum_out[8][14][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][14][16] = (sum_out[9][14][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][14][16] = (sum_out[10][14][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][14][16] = (sum_out[11][14][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][14][16] = (sum_out[12][14][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][14][16] = (sum_out[13][14][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][14][16] = (sum_out[14][14][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][14][16] = (sum_out[15][14][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][14][16] = (sum_out[16][14][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][14][16] = (sum_out[17][14][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][14][16] = (sum_out[18][14][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][14][16] = (sum_out[19][14][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][14][17] = (sum_out[0][14][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][14][17] = (sum_out[1][14][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][14][17] = (sum_out[2][14][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][14][17] = (sum_out[3][14][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][14][17] = (sum_out[4][14][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][14][17] = (sum_out[5][14][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][14][17] = (sum_out[6][14][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][14][17] = (sum_out[7][14][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][14][17] = (sum_out[8][14][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][14][17] = (sum_out[9][14][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][14][17] = (sum_out[10][14][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][14][17] = (sum_out[11][14][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][14][17] = (sum_out[12][14][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][14][17] = (sum_out[13][14][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][14][17] = (sum_out[14][14][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][14][17] = (sum_out[15][14][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][14][17] = (sum_out[16][14][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][14][17] = (sum_out[17][14][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][14][17] = (sum_out[18][14][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][14][17] = (sum_out[19][14][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][14][18] = (sum_out[0][14][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][14][18] = (sum_out[1][14][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][14][18] = (sum_out[2][14][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][14][18] = (sum_out[3][14][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][14][18] = (sum_out[4][14][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][14][18] = (sum_out[5][14][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][14][18] = (sum_out[6][14][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][14][18] = (sum_out[7][14][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][14][18] = (sum_out[8][14][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][14][18] = (sum_out[9][14][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][14][18] = (sum_out[10][14][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][14][18] = (sum_out[11][14][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][14][18] = (sum_out[12][14][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][14][18] = (sum_out[13][14][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][14][18] = (sum_out[14][14][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][14][18] = (sum_out[15][14][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][14][18] = (sum_out[16][14][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][14][18] = (sum_out[17][14][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][14][18] = (sum_out[18][14][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][14][18] = (sum_out[19][14][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][14][19] = (sum_out[0][14][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][14][19] = (sum_out[1][14][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][14][19] = (sum_out[2][14][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][14][19] = (sum_out[3][14][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][14][19] = (sum_out[4][14][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][14][19] = (sum_out[5][14][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][14][19] = (sum_out[6][14][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][14][19] = (sum_out[7][14][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][14][19] = (sum_out[8][14][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][14][19] = (sum_out[9][14][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][14][19] = (sum_out[10][14][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][14][19] = (sum_out[11][14][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][14][19] = (sum_out[12][14][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][14][19] = (sum_out[13][14][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][14][19] = (sum_out[14][14][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][14][19] = (sum_out[15][14][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][14][19] = (sum_out[16][14][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][14][19] = (sum_out[17][14][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][14][19] = (sum_out[18][14][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][14][19] = (sum_out[19][14][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][14][20] = (sum_out[0][14][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][14][20] = (sum_out[1][14][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][14][20] = (sum_out[2][14][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][14][20] = (sum_out[3][14][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][14][20] = (sum_out[4][14][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][14][20] = (sum_out[5][14][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][14][20] = (sum_out[6][14][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][14][20] = (sum_out[7][14][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][14][20] = (sum_out[8][14][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][14][20] = (sum_out[9][14][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][14][20] = (sum_out[10][14][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][14][20] = (sum_out[11][14][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][14][20] = (sum_out[12][14][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][14][20] = (sum_out[13][14][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][14][20] = (sum_out[14][14][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][14][20] = (sum_out[15][14][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][14][20] = (sum_out[16][14][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][14][20] = (sum_out[17][14][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][14][20] = (sum_out[18][14][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][14][20] = (sum_out[19][14][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][14][21] = (sum_out[0][14][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][14][21] = (sum_out[1][14][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][14][21] = (sum_out[2][14][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][14][21] = (sum_out[3][14][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][14][21] = (sum_out[4][14][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][14][21] = (sum_out[5][14][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][14][21] = (sum_out[6][14][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][14][21] = (sum_out[7][14][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][14][21] = (sum_out[8][14][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][14][21] = (sum_out[9][14][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][14][21] = (sum_out[10][14][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][14][21] = (sum_out[11][14][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][14][21] = (sum_out[12][14][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][14][21] = (sum_out[13][14][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][14][21] = (sum_out[14][14][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][14][21] = (sum_out[15][14][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][14][21] = (sum_out[16][14][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][14][21] = (sum_out[17][14][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][14][21] = (sum_out[18][14][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][14][21] = (sum_out[19][14][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][14][22] = (sum_out[0][14][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][14][22] = (sum_out[1][14][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][14][22] = (sum_out[2][14][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][14][22] = (sum_out[3][14][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][14][22] = (sum_out[4][14][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][14][22] = (sum_out[5][14][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][14][22] = (sum_out[6][14][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][14][22] = (sum_out[7][14][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][14][22] = (sum_out[8][14][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][14][22] = (sum_out[9][14][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][14][22] = (sum_out[10][14][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][14][22] = (sum_out[11][14][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][14][22] = (sum_out[12][14][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][14][22] = (sum_out[13][14][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][14][22] = (sum_out[14][14][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][14][22] = (sum_out[15][14][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][14][22] = (sum_out[16][14][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][14][22] = (sum_out[17][14][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][14][22] = (sum_out[18][14][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][14][22] = (sum_out[19][14][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][14][23] = (sum_out[0][14][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][14][23] = (sum_out[1][14][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][14][23] = (sum_out[2][14][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][14][23] = (sum_out[3][14][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][14][23] = (sum_out[4][14][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][14][23] = (sum_out[5][14][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][14][23] = (sum_out[6][14][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][14][23] = (sum_out[7][14][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][14][23] = (sum_out[8][14][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][14][23] = (sum_out[9][14][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][14][23] = (sum_out[10][14][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][14][23] = (sum_out[11][14][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][14][23] = (sum_out[12][14][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][14][23] = (sum_out[13][14][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][14][23] = (sum_out[14][14][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][14][23] = (sum_out[15][14][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][14][23] = (sum_out[16][14][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][14][23] = (sum_out[17][14][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][14][23] = (sum_out[18][14][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][14][23] = (sum_out[19][14][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][15][0] = (sum_out[0][15][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][15][0] = (sum_out[1][15][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][15][0] = (sum_out[2][15][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][15][0] = (sum_out[3][15][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][15][0] = (sum_out[4][15][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][15][0] = (sum_out[5][15][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][15][0] = (sum_out[6][15][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][15][0] = (sum_out[7][15][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][15][0] = (sum_out[8][15][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][15][0] = (sum_out[9][15][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][15][0] = (sum_out[10][15][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][15][0] = (sum_out[11][15][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][15][0] = (sum_out[12][15][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][15][0] = (sum_out[13][15][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][15][0] = (sum_out[14][15][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][15][0] = (sum_out[15][15][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][15][0] = (sum_out[16][15][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][15][0] = (sum_out[17][15][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][15][0] = (sum_out[18][15][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][15][0] = (sum_out[19][15][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][15][1] = (sum_out[0][15][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][15][1] = (sum_out[1][15][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][15][1] = (sum_out[2][15][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][15][1] = (sum_out[3][15][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][15][1] = (sum_out[4][15][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][15][1] = (sum_out[5][15][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][15][1] = (sum_out[6][15][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][15][1] = (sum_out[7][15][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][15][1] = (sum_out[8][15][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][15][1] = (sum_out[9][15][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][15][1] = (sum_out[10][15][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][15][1] = (sum_out[11][15][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][15][1] = (sum_out[12][15][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][15][1] = (sum_out[13][15][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][15][1] = (sum_out[14][15][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][15][1] = (sum_out[15][15][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][15][1] = (sum_out[16][15][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][15][1] = (sum_out[17][15][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][15][1] = (sum_out[18][15][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][15][1] = (sum_out[19][15][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][15][2] = (sum_out[0][15][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][15][2] = (sum_out[1][15][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][15][2] = (sum_out[2][15][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][15][2] = (sum_out[3][15][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][15][2] = (sum_out[4][15][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][15][2] = (sum_out[5][15][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][15][2] = (sum_out[6][15][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][15][2] = (sum_out[7][15][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][15][2] = (sum_out[8][15][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][15][2] = (sum_out[9][15][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][15][2] = (sum_out[10][15][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][15][2] = (sum_out[11][15][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][15][2] = (sum_out[12][15][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][15][2] = (sum_out[13][15][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][15][2] = (sum_out[14][15][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][15][2] = (sum_out[15][15][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][15][2] = (sum_out[16][15][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][15][2] = (sum_out[17][15][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][15][2] = (sum_out[18][15][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][15][2] = (sum_out[19][15][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][15][3] = (sum_out[0][15][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][15][3] = (sum_out[1][15][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][15][3] = (sum_out[2][15][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][15][3] = (sum_out[3][15][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][15][3] = (sum_out[4][15][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][15][3] = (sum_out[5][15][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][15][3] = (sum_out[6][15][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][15][3] = (sum_out[7][15][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][15][3] = (sum_out[8][15][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][15][3] = (sum_out[9][15][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][15][3] = (sum_out[10][15][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][15][3] = (sum_out[11][15][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][15][3] = (sum_out[12][15][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][15][3] = (sum_out[13][15][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][15][3] = (sum_out[14][15][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][15][3] = (sum_out[15][15][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][15][3] = (sum_out[16][15][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][15][3] = (sum_out[17][15][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][15][3] = (sum_out[18][15][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][15][3] = (sum_out[19][15][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][15][4] = (sum_out[0][15][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][15][4] = (sum_out[1][15][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][15][4] = (sum_out[2][15][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][15][4] = (sum_out[3][15][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][15][4] = (sum_out[4][15][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][15][4] = (sum_out[5][15][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][15][4] = (sum_out[6][15][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][15][4] = (sum_out[7][15][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][15][4] = (sum_out[8][15][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][15][4] = (sum_out[9][15][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][15][4] = (sum_out[10][15][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][15][4] = (sum_out[11][15][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][15][4] = (sum_out[12][15][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][15][4] = (sum_out[13][15][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][15][4] = (sum_out[14][15][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][15][4] = (sum_out[15][15][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][15][4] = (sum_out[16][15][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][15][4] = (sum_out[17][15][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][15][4] = (sum_out[18][15][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][15][4] = (sum_out[19][15][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][15][5] = (sum_out[0][15][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][15][5] = (sum_out[1][15][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][15][5] = (sum_out[2][15][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][15][5] = (sum_out[3][15][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][15][5] = (sum_out[4][15][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][15][5] = (sum_out[5][15][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][15][5] = (sum_out[6][15][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][15][5] = (sum_out[7][15][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][15][5] = (sum_out[8][15][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][15][5] = (sum_out[9][15][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][15][5] = (sum_out[10][15][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][15][5] = (sum_out[11][15][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][15][5] = (sum_out[12][15][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][15][5] = (sum_out[13][15][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][15][5] = (sum_out[14][15][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][15][5] = (sum_out[15][15][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][15][5] = (sum_out[16][15][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][15][5] = (sum_out[17][15][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][15][5] = (sum_out[18][15][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][15][5] = (sum_out[19][15][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][15][6] = (sum_out[0][15][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][15][6] = (sum_out[1][15][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][15][6] = (sum_out[2][15][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][15][6] = (sum_out[3][15][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][15][6] = (sum_out[4][15][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][15][6] = (sum_out[5][15][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][15][6] = (sum_out[6][15][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][15][6] = (sum_out[7][15][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][15][6] = (sum_out[8][15][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][15][6] = (sum_out[9][15][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][15][6] = (sum_out[10][15][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][15][6] = (sum_out[11][15][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][15][6] = (sum_out[12][15][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][15][6] = (sum_out[13][15][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][15][6] = (sum_out[14][15][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][15][6] = (sum_out[15][15][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][15][6] = (sum_out[16][15][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][15][6] = (sum_out[17][15][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][15][6] = (sum_out[18][15][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][15][6] = (sum_out[19][15][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][15][7] = (sum_out[0][15][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][15][7] = (sum_out[1][15][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][15][7] = (sum_out[2][15][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][15][7] = (sum_out[3][15][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][15][7] = (sum_out[4][15][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][15][7] = (sum_out[5][15][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][15][7] = (sum_out[6][15][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][15][7] = (sum_out[7][15][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][15][7] = (sum_out[8][15][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][15][7] = (sum_out[9][15][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][15][7] = (sum_out[10][15][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][15][7] = (sum_out[11][15][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][15][7] = (sum_out[12][15][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][15][7] = (sum_out[13][15][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][15][7] = (sum_out[14][15][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][15][7] = (sum_out[15][15][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][15][7] = (sum_out[16][15][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][15][7] = (sum_out[17][15][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][15][7] = (sum_out[18][15][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][15][7] = (sum_out[19][15][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][15][8] = (sum_out[0][15][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][15][8] = (sum_out[1][15][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][15][8] = (sum_out[2][15][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][15][8] = (sum_out[3][15][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][15][8] = (sum_out[4][15][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][15][8] = (sum_out[5][15][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][15][8] = (sum_out[6][15][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][15][8] = (sum_out[7][15][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][15][8] = (sum_out[8][15][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][15][8] = (sum_out[9][15][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][15][8] = (sum_out[10][15][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][15][8] = (sum_out[11][15][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][15][8] = (sum_out[12][15][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][15][8] = (sum_out[13][15][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][15][8] = (sum_out[14][15][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][15][8] = (sum_out[15][15][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][15][8] = (sum_out[16][15][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][15][8] = (sum_out[17][15][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][15][8] = (sum_out[18][15][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][15][8] = (sum_out[19][15][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][15][9] = (sum_out[0][15][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][15][9] = (sum_out[1][15][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][15][9] = (sum_out[2][15][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][15][9] = (sum_out[3][15][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][15][9] = (sum_out[4][15][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][15][9] = (sum_out[5][15][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][15][9] = (sum_out[6][15][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][15][9] = (sum_out[7][15][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][15][9] = (sum_out[8][15][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][15][9] = (sum_out[9][15][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][15][9] = (sum_out[10][15][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][15][9] = (sum_out[11][15][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][15][9] = (sum_out[12][15][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][15][9] = (sum_out[13][15][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][15][9] = (sum_out[14][15][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][15][9] = (sum_out[15][15][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][15][9] = (sum_out[16][15][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][15][9] = (sum_out[17][15][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][15][9] = (sum_out[18][15][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][15][9] = (sum_out[19][15][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][15][10] = (sum_out[0][15][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][15][10] = (sum_out[1][15][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][15][10] = (sum_out[2][15][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][15][10] = (sum_out[3][15][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][15][10] = (sum_out[4][15][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][15][10] = (sum_out[5][15][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][15][10] = (sum_out[6][15][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][15][10] = (sum_out[7][15][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][15][10] = (sum_out[8][15][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][15][10] = (sum_out[9][15][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][15][10] = (sum_out[10][15][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][15][10] = (sum_out[11][15][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][15][10] = (sum_out[12][15][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][15][10] = (sum_out[13][15][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][15][10] = (sum_out[14][15][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][15][10] = (sum_out[15][15][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][15][10] = (sum_out[16][15][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][15][10] = (sum_out[17][15][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][15][10] = (sum_out[18][15][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][15][10] = (sum_out[19][15][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][15][11] = (sum_out[0][15][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][15][11] = (sum_out[1][15][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][15][11] = (sum_out[2][15][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][15][11] = (sum_out[3][15][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][15][11] = (sum_out[4][15][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][15][11] = (sum_out[5][15][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][15][11] = (sum_out[6][15][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][15][11] = (sum_out[7][15][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][15][11] = (sum_out[8][15][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][15][11] = (sum_out[9][15][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][15][11] = (sum_out[10][15][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][15][11] = (sum_out[11][15][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][15][11] = (sum_out[12][15][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][15][11] = (sum_out[13][15][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][15][11] = (sum_out[14][15][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][15][11] = (sum_out[15][15][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][15][11] = (sum_out[16][15][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][15][11] = (sum_out[17][15][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][15][11] = (sum_out[18][15][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][15][11] = (sum_out[19][15][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][15][12] = (sum_out[0][15][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][15][12] = (sum_out[1][15][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][15][12] = (sum_out[2][15][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][15][12] = (sum_out[3][15][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][15][12] = (sum_out[4][15][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][15][12] = (sum_out[5][15][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][15][12] = (sum_out[6][15][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][15][12] = (sum_out[7][15][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][15][12] = (sum_out[8][15][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][15][12] = (sum_out[9][15][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][15][12] = (sum_out[10][15][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][15][12] = (sum_out[11][15][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][15][12] = (sum_out[12][15][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][15][12] = (sum_out[13][15][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][15][12] = (sum_out[14][15][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][15][12] = (sum_out[15][15][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][15][12] = (sum_out[16][15][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][15][12] = (sum_out[17][15][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][15][12] = (sum_out[18][15][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][15][12] = (sum_out[19][15][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][15][13] = (sum_out[0][15][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][15][13] = (sum_out[1][15][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][15][13] = (sum_out[2][15][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][15][13] = (sum_out[3][15][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][15][13] = (sum_out[4][15][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][15][13] = (sum_out[5][15][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][15][13] = (sum_out[6][15][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][15][13] = (sum_out[7][15][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][15][13] = (sum_out[8][15][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][15][13] = (sum_out[9][15][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][15][13] = (sum_out[10][15][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][15][13] = (sum_out[11][15][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][15][13] = (sum_out[12][15][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][15][13] = (sum_out[13][15][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][15][13] = (sum_out[14][15][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][15][13] = (sum_out[15][15][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][15][13] = (sum_out[16][15][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][15][13] = (sum_out[17][15][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][15][13] = (sum_out[18][15][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][15][13] = (sum_out[19][15][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][15][14] = (sum_out[0][15][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][15][14] = (sum_out[1][15][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][15][14] = (sum_out[2][15][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][15][14] = (sum_out[3][15][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][15][14] = (sum_out[4][15][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][15][14] = (sum_out[5][15][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][15][14] = (sum_out[6][15][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][15][14] = (sum_out[7][15][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][15][14] = (sum_out[8][15][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][15][14] = (sum_out[9][15][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][15][14] = (sum_out[10][15][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][15][14] = (sum_out[11][15][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][15][14] = (sum_out[12][15][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][15][14] = (sum_out[13][15][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][15][14] = (sum_out[14][15][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][15][14] = (sum_out[15][15][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][15][14] = (sum_out[16][15][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][15][14] = (sum_out[17][15][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][15][14] = (sum_out[18][15][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][15][14] = (sum_out[19][15][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][15][15] = (sum_out[0][15][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][15][15] = (sum_out[1][15][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][15][15] = (sum_out[2][15][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][15][15] = (sum_out[3][15][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][15][15] = (sum_out[4][15][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][15][15] = (sum_out[5][15][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][15][15] = (sum_out[6][15][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][15][15] = (sum_out[7][15][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][15][15] = (sum_out[8][15][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][15][15] = (sum_out[9][15][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][15][15] = (sum_out[10][15][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][15][15] = (sum_out[11][15][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][15][15] = (sum_out[12][15][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][15][15] = (sum_out[13][15][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][15][15] = (sum_out[14][15][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][15][15] = (sum_out[15][15][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][15][15] = (sum_out[16][15][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][15][15] = (sum_out[17][15][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][15][15] = (sum_out[18][15][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][15][15] = (sum_out[19][15][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][15][16] = (sum_out[0][15][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][15][16] = (sum_out[1][15][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][15][16] = (sum_out[2][15][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][15][16] = (sum_out[3][15][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][15][16] = (sum_out[4][15][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][15][16] = (sum_out[5][15][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][15][16] = (sum_out[6][15][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][15][16] = (sum_out[7][15][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][15][16] = (sum_out[8][15][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][15][16] = (sum_out[9][15][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][15][16] = (sum_out[10][15][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][15][16] = (sum_out[11][15][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][15][16] = (sum_out[12][15][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][15][16] = (sum_out[13][15][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][15][16] = (sum_out[14][15][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][15][16] = (sum_out[15][15][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][15][16] = (sum_out[16][15][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][15][16] = (sum_out[17][15][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][15][16] = (sum_out[18][15][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][15][16] = (sum_out[19][15][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][15][17] = (sum_out[0][15][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][15][17] = (sum_out[1][15][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][15][17] = (sum_out[2][15][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][15][17] = (sum_out[3][15][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][15][17] = (sum_out[4][15][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][15][17] = (sum_out[5][15][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][15][17] = (sum_out[6][15][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][15][17] = (sum_out[7][15][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][15][17] = (sum_out[8][15][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][15][17] = (sum_out[9][15][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][15][17] = (sum_out[10][15][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][15][17] = (sum_out[11][15][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][15][17] = (sum_out[12][15][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][15][17] = (sum_out[13][15][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][15][17] = (sum_out[14][15][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][15][17] = (sum_out[15][15][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][15][17] = (sum_out[16][15][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][15][17] = (sum_out[17][15][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][15][17] = (sum_out[18][15][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][15][17] = (sum_out[19][15][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][15][18] = (sum_out[0][15][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][15][18] = (sum_out[1][15][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][15][18] = (sum_out[2][15][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][15][18] = (sum_out[3][15][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][15][18] = (sum_out[4][15][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][15][18] = (sum_out[5][15][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][15][18] = (sum_out[6][15][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][15][18] = (sum_out[7][15][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][15][18] = (sum_out[8][15][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][15][18] = (sum_out[9][15][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][15][18] = (sum_out[10][15][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][15][18] = (sum_out[11][15][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][15][18] = (sum_out[12][15][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][15][18] = (sum_out[13][15][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][15][18] = (sum_out[14][15][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][15][18] = (sum_out[15][15][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][15][18] = (sum_out[16][15][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][15][18] = (sum_out[17][15][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][15][18] = (sum_out[18][15][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][15][18] = (sum_out[19][15][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][15][19] = (sum_out[0][15][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][15][19] = (sum_out[1][15][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][15][19] = (sum_out[2][15][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][15][19] = (sum_out[3][15][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][15][19] = (sum_out[4][15][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][15][19] = (sum_out[5][15][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][15][19] = (sum_out[6][15][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][15][19] = (sum_out[7][15][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][15][19] = (sum_out[8][15][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][15][19] = (sum_out[9][15][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][15][19] = (sum_out[10][15][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][15][19] = (sum_out[11][15][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][15][19] = (sum_out[12][15][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][15][19] = (sum_out[13][15][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][15][19] = (sum_out[14][15][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][15][19] = (sum_out[15][15][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][15][19] = (sum_out[16][15][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][15][19] = (sum_out[17][15][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][15][19] = (sum_out[18][15][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][15][19] = (sum_out[19][15][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][15][20] = (sum_out[0][15][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][15][20] = (sum_out[1][15][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][15][20] = (sum_out[2][15][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][15][20] = (sum_out[3][15][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][15][20] = (sum_out[4][15][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][15][20] = (sum_out[5][15][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][15][20] = (sum_out[6][15][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][15][20] = (sum_out[7][15][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][15][20] = (sum_out[8][15][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][15][20] = (sum_out[9][15][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][15][20] = (sum_out[10][15][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][15][20] = (sum_out[11][15][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][15][20] = (sum_out[12][15][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][15][20] = (sum_out[13][15][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][15][20] = (sum_out[14][15][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][15][20] = (sum_out[15][15][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][15][20] = (sum_out[16][15][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][15][20] = (sum_out[17][15][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][15][20] = (sum_out[18][15][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][15][20] = (sum_out[19][15][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][15][21] = (sum_out[0][15][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][15][21] = (sum_out[1][15][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][15][21] = (sum_out[2][15][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][15][21] = (sum_out[3][15][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][15][21] = (sum_out[4][15][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][15][21] = (sum_out[5][15][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][15][21] = (sum_out[6][15][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][15][21] = (sum_out[7][15][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][15][21] = (sum_out[8][15][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][15][21] = (sum_out[9][15][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][15][21] = (sum_out[10][15][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][15][21] = (sum_out[11][15][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][15][21] = (sum_out[12][15][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][15][21] = (sum_out[13][15][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][15][21] = (sum_out[14][15][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][15][21] = (sum_out[15][15][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][15][21] = (sum_out[16][15][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][15][21] = (sum_out[17][15][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][15][21] = (sum_out[18][15][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][15][21] = (sum_out[19][15][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][15][22] = (sum_out[0][15][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][15][22] = (sum_out[1][15][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][15][22] = (sum_out[2][15][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][15][22] = (sum_out[3][15][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][15][22] = (sum_out[4][15][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][15][22] = (sum_out[5][15][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][15][22] = (sum_out[6][15][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][15][22] = (sum_out[7][15][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][15][22] = (sum_out[8][15][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][15][22] = (sum_out[9][15][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][15][22] = (sum_out[10][15][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][15][22] = (sum_out[11][15][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][15][22] = (sum_out[12][15][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][15][22] = (sum_out[13][15][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][15][22] = (sum_out[14][15][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][15][22] = (sum_out[15][15][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][15][22] = (sum_out[16][15][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][15][22] = (sum_out[17][15][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][15][22] = (sum_out[18][15][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][15][22] = (sum_out[19][15][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][15][23] = (sum_out[0][15][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][15][23] = (sum_out[1][15][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][15][23] = (sum_out[2][15][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][15][23] = (sum_out[3][15][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][15][23] = (sum_out[4][15][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][15][23] = (sum_out[5][15][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][15][23] = (sum_out[6][15][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][15][23] = (sum_out[7][15][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][15][23] = (sum_out[8][15][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][15][23] = (sum_out[9][15][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][15][23] = (sum_out[10][15][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][15][23] = (sum_out[11][15][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][15][23] = (sum_out[12][15][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][15][23] = (sum_out[13][15][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][15][23] = (sum_out[14][15][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][15][23] = (sum_out[15][15][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][15][23] = (sum_out[16][15][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][15][23] = (sum_out[17][15][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][15][23] = (sum_out[18][15][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][15][23] = (sum_out[19][15][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][16][0] = (sum_out[0][16][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][16][0] = (sum_out[1][16][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][16][0] = (sum_out[2][16][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][16][0] = (sum_out[3][16][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][16][0] = (sum_out[4][16][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][16][0] = (sum_out[5][16][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][16][0] = (sum_out[6][16][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][16][0] = (sum_out[7][16][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][16][0] = (sum_out[8][16][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][16][0] = (sum_out[9][16][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][16][0] = (sum_out[10][16][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][16][0] = (sum_out[11][16][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][16][0] = (sum_out[12][16][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][16][0] = (sum_out[13][16][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][16][0] = (sum_out[14][16][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][16][0] = (sum_out[15][16][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][16][0] = (sum_out[16][16][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][16][0] = (sum_out[17][16][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][16][0] = (sum_out[18][16][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][16][0] = (sum_out[19][16][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][16][1] = (sum_out[0][16][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][16][1] = (sum_out[1][16][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][16][1] = (sum_out[2][16][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][16][1] = (sum_out[3][16][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][16][1] = (sum_out[4][16][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][16][1] = (sum_out[5][16][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][16][1] = (sum_out[6][16][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][16][1] = (sum_out[7][16][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][16][1] = (sum_out[8][16][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][16][1] = (sum_out[9][16][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][16][1] = (sum_out[10][16][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][16][1] = (sum_out[11][16][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][16][1] = (sum_out[12][16][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][16][1] = (sum_out[13][16][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][16][1] = (sum_out[14][16][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][16][1] = (sum_out[15][16][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][16][1] = (sum_out[16][16][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][16][1] = (sum_out[17][16][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][16][1] = (sum_out[18][16][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][16][1] = (sum_out[19][16][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][16][2] = (sum_out[0][16][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][16][2] = (sum_out[1][16][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][16][2] = (sum_out[2][16][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][16][2] = (sum_out[3][16][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][16][2] = (sum_out[4][16][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][16][2] = (sum_out[5][16][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][16][2] = (sum_out[6][16][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][16][2] = (sum_out[7][16][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][16][2] = (sum_out[8][16][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][16][2] = (sum_out[9][16][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][16][2] = (sum_out[10][16][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][16][2] = (sum_out[11][16][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][16][2] = (sum_out[12][16][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][16][2] = (sum_out[13][16][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][16][2] = (sum_out[14][16][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][16][2] = (sum_out[15][16][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][16][2] = (sum_out[16][16][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][16][2] = (sum_out[17][16][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][16][2] = (sum_out[18][16][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][16][2] = (sum_out[19][16][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][16][3] = (sum_out[0][16][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][16][3] = (sum_out[1][16][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][16][3] = (sum_out[2][16][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][16][3] = (sum_out[3][16][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][16][3] = (sum_out[4][16][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][16][3] = (sum_out[5][16][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][16][3] = (sum_out[6][16][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][16][3] = (sum_out[7][16][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][16][3] = (sum_out[8][16][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][16][3] = (sum_out[9][16][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][16][3] = (sum_out[10][16][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][16][3] = (sum_out[11][16][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][16][3] = (sum_out[12][16][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][16][3] = (sum_out[13][16][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][16][3] = (sum_out[14][16][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][16][3] = (sum_out[15][16][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][16][3] = (sum_out[16][16][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][16][3] = (sum_out[17][16][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][16][3] = (sum_out[18][16][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][16][3] = (sum_out[19][16][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][16][4] = (sum_out[0][16][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][16][4] = (sum_out[1][16][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][16][4] = (sum_out[2][16][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][16][4] = (sum_out[3][16][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][16][4] = (sum_out[4][16][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][16][4] = (sum_out[5][16][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][16][4] = (sum_out[6][16][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][16][4] = (sum_out[7][16][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][16][4] = (sum_out[8][16][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][16][4] = (sum_out[9][16][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][16][4] = (sum_out[10][16][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][16][4] = (sum_out[11][16][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][16][4] = (sum_out[12][16][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][16][4] = (sum_out[13][16][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][16][4] = (sum_out[14][16][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][16][4] = (sum_out[15][16][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][16][4] = (sum_out[16][16][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][16][4] = (sum_out[17][16][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][16][4] = (sum_out[18][16][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][16][4] = (sum_out[19][16][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][16][5] = (sum_out[0][16][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][16][5] = (sum_out[1][16][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][16][5] = (sum_out[2][16][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][16][5] = (sum_out[3][16][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][16][5] = (sum_out[4][16][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][16][5] = (sum_out[5][16][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][16][5] = (sum_out[6][16][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][16][5] = (sum_out[7][16][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][16][5] = (sum_out[8][16][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][16][5] = (sum_out[9][16][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][16][5] = (sum_out[10][16][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][16][5] = (sum_out[11][16][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][16][5] = (sum_out[12][16][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][16][5] = (sum_out[13][16][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][16][5] = (sum_out[14][16][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][16][5] = (sum_out[15][16][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][16][5] = (sum_out[16][16][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][16][5] = (sum_out[17][16][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][16][5] = (sum_out[18][16][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][16][5] = (sum_out[19][16][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][16][6] = (sum_out[0][16][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][16][6] = (sum_out[1][16][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][16][6] = (sum_out[2][16][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][16][6] = (sum_out[3][16][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][16][6] = (sum_out[4][16][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][16][6] = (sum_out[5][16][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][16][6] = (sum_out[6][16][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][16][6] = (sum_out[7][16][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][16][6] = (sum_out[8][16][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][16][6] = (sum_out[9][16][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][16][6] = (sum_out[10][16][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][16][6] = (sum_out[11][16][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][16][6] = (sum_out[12][16][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][16][6] = (sum_out[13][16][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][16][6] = (sum_out[14][16][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][16][6] = (sum_out[15][16][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][16][6] = (sum_out[16][16][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][16][6] = (sum_out[17][16][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][16][6] = (sum_out[18][16][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][16][6] = (sum_out[19][16][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][16][7] = (sum_out[0][16][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][16][7] = (sum_out[1][16][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][16][7] = (sum_out[2][16][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][16][7] = (sum_out[3][16][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][16][7] = (sum_out[4][16][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][16][7] = (sum_out[5][16][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][16][7] = (sum_out[6][16][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][16][7] = (sum_out[7][16][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][16][7] = (sum_out[8][16][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][16][7] = (sum_out[9][16][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][16][7] = (sum_out[10][16][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][16][7] = (sum_out[11][16][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][16][7] = (sum_out[12][16][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][16][7] = (sum_out[13][16][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][16][7] = (sum_out[14][16][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][16][7] = (sum_out[15][16][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][16][7] = (sum_out[16][16][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][16][7] = (sum_out[17][16][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][16][7] = (sum_out[18][16][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][16][7] = (sum_out[19][16][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][16][8] = (sum_out[0][16][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][16][8] = (sum_out[1][16][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][16][8] = (sum_out[2][16][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][16][8] = (sum_out[3][16][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][16][8] = (sum_out[4][16][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][16][8] = (sum_out[5][16][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][16][8] = (sum_out[6][16][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][16][8] = (sum_out[7][16][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][16][8] = (sum_out[8][16][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][16][8] = (sum_out[9][16][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][16][8] = (sum_out[10][16][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][16][8] = (sum_out[11][16][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][16][8] = (sum_out[12][16][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][16][8] = (sum_out[13][16][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][16][8] = (sum_out[14][16][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][16][8] = (sum_out[15][16][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][16][8] = (sum_out[16][16][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][16][8] = (sum_out[17][16][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][16][8] = (sum_out[18][16][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][16][8] = (sum_out[19][16][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][16][9] = (sum_out[0][16][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][16][9] = (sum_out[1][16][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][16][9] = (sum_out[2][16][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][16][9] = (sum_out[3][16][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][16][9] = (sum_out[4][16][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][16][9] = (sum_out[5][16][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][16][9] = (sum_out[6][16][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][16][9] = (sum_out[7][16][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][16][9] = (sum_out[8][16][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][16][9] = (sum_out[9][16][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][16][9] = (sum_out[10][16][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][16][9] = (sum_out[11][16][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][16][9] = (sum_out[12][16][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][16][9] = (sum_out[13][16][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][16][9] = (sum_out[14][16][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][16][9] = (sum_out[15][16][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][16][9] = (sum_out[16][16][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][16][9] = (sum_out[17][16][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][16][9] = (sum_out[18][16][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][16][9] = (sum_out[19][16][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][16][10] = (sum_out[0][16][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][16][10] = (sum_out[1][16][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][16][10] = (sum_out[2][16][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][16][10] = (sum_out[3][16][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][16][10] = (sum_out[4][16][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][16][10] = (sum_out[5][16][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][16][10] = (sum_out[6][16][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][16][10] = (sum_out[7][16][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][16][10] = (sum_out[8][16][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][16][10] = (sum_out[9][16][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][16][10] = (sum_out[10][16][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][16][10] = (sum_out[11][16][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][16][10] = (sum_out[12][16][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][16][10] = (sum_out[13][16][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][16][10] = (sum_out[14][16][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][16][10] = (sum_out[15][16][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][16][10] = (sum_out[16][16][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][16][10] = (sum_out[17][16][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][16][10] = (sum_out[18][16][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][16][10] = (sum_out[19][16][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][16][11] = (sum_out[0][16][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][16][11] = (sum_out[1][16][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][16][11] = (sum_out[2][16][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][16][11] = (sum_out[3][16][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][16][11] = (sum_out[4][16][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][16][11] = (sum_out[5][16][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][16][11] = (sum_out[6][16][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][16][11] = (sum_out[7][16][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][16][11] = (sum_out[8][16][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][16][11] = (sum_out[9][16][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][16][11] = (sum_out[10][16][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][16][11] = (sum_out[11][16][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][16][11] = (sum_out[12][16][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][16][11] = (sum_out[13][16][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][16][11] = (sum_out[14][16][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][16][11] = (sum_out[15][16][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][16][11] = (sum_out[16][16][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][16][11] = (sum_out[17][16][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][16][11] = (sum_out[18][16][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][16][11] = (sum_out[19][16][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][16][12] = (sum_out[0][16][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][16][12] = (sum_out[1][16][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][16][12] = (sum_out[2][16][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][16][12] = (sum_out[3][16][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][16][12] = (sum_out[4][16][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][16][12] = (sum_out[5][16][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][16][12] = (sum_out[6][16][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][16][12] = (sum_out[7][16][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][16][12] = (sum_out[8][16][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][16][12] = (sum_out[9][16][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][16][12] = (sum_out[10][16][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][16][12] = (sum_out[11][16][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][16][12] = (sum_out[12][16][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][16][12] = (sum_out[13][16][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][16][12] = (sum_out[14][16][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][16][12] = (sum_out[15][16][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][16][12] = (sum_out[16][16][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][16][12] = (sum_out[17][16][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][16][12] = (sum_out[18][16][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][16][12] = (sum_out[19][16][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][16][13] = (sum_out[0][16][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][16][13] = (sum_out[1][16][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][16][13] = (sum_out[2][16][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][16][13] = (sum_out[3][16][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][16][13] = (sum_out[4][16][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][16][13] = (sum_out[5][16][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][16][13] = (sum_out[6][16][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][16][13] = (sum_out[7][16][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][16][13] = (sum_out[8][16][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][16][13] = (sum_out[9][16][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][16][13] = (sum_out[10][16][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][16][13] = (sum_out[11][16][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][16][13] = (sum_out[12][16][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][16][13] = (sum_out[13][16][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][16][13] = (sum_out[14][16][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][16][13] = (sum_out[15][16][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][16][13] = (sum_out[16][16][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][16][13] = (sum_out[17][16][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][16][13] = (sum_out[18][16][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][16][13] = (sum_out[19][16][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][16][14] = (sum_out[0][16][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][16][14] = (sum_out[1][16][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][16][14] = (sum_out[2][16][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][16][14] = (sum_out[3][16][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][16][14] = (sum_out[4][16][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][16][14] = (sum_out[5][16][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][16][14] = (sum_out[6][16][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][16][14] = (sum_out[7][16][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][16][14] = (sum_out[8][16][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][16][14] = (sum_out[9][16][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][16][14] = (sum_out[10][16][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][16][14] = (sum_out[11][16][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][16][14] = (sum_out[12][16][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][16][14] = (sum_out[13][16][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][16][14] = (sum_out[14][16][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][16][14] = (sum_out[15][16][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][16][14] = (sum_out[16][16][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][16][14] = (sum_out[17][16][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][16][14] = (sum_out[18][16][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][16][14] = (sum_out[19][16][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][16][15] = (sum_out[0][16][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][16][15] = (sum_out[1][16][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][16][15] = (sum_out[2][16][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][16][15] = (sum_out[3][16][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][16][15] = (sum_out[4][16][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][16][15] = (sum_out[5][16][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][16][15] = (sum_out[6][16][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][16][15] = (sum_out[7][16][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][16][15] = (sum_out[8][16][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][16][15] = (sum_out[9][16][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][16][15] = (sum_out[10][16][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][16][15] = (sum_out[11][16][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][16][15] = (sum_out[12][16][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][16][15] = (sum_out[13][16][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][16][15] = (sum_out[14][16][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][16][15] = (sum_out[15][16][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][16][15] = (sum_out[16][16][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][16][15] = (sum_out[17][16][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][16][15] = (sum_out[18][16][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][16][15] = (sum_out[19][16][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][16][16] = (sum_out[0][16][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][16][16] = (sum_out[1][16][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][16][16] = (sum_out[2][16][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][16][16] = (sum_out[3][16][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][16][16] = (sum_out[4][16][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][16][16] = (sum_out[5][16][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][16][16] = (sum_out[6][16][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][16][16] = (sum_out[7][16][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][16][16] = (sum_out[8][16][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][16][16] = (sum_out[9][16][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][16][16] = (sum_out[10][16][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][16][16] = (sum_out[11][16][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][16][16] = (sum_out[12][16][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][16][16] = (sum_out[13][16][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][16][16] = (sum_out[14][16][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][16][16] = (sum_out[15][16][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][16][16] = (sum_out[16][16][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][16][16] = (sum_out[17][16][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][16][16] = (sum_out[18][16][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][16][16] = (sum_out[19][16][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][16][17] = (sum_out[0][16][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][16][17] = (sum_out[1][16][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][16][17] = (sum_out[2][16][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][16][17] = (sum_out[3][16][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][16][17] = (sum_out[4][16][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][16][17] = (sum_out[5][16][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][16][17] = (sum_out[6][16][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][16][17] = (sum_out[7][16][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][16][17] = (sum_out[8][16][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][16][17] = (sum_out[9][16][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][16][17] = (sum_out[10][16][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][16][17] = (sum_out[11][16][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][16][17] = (sum_out[12][16][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][16][17] = (sum_out[13][16][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][16][17] = (sum_out[14][16][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][16][17] = (sum_out[15][16][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][16][17] = (sum_out[16][16][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][16][17] = (sum_out[17][16][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][16][17] = (sum_out[18][16][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][16][17] = (sum_out[19][16][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][16][18] = (sum_out[0][16][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][16][18] = (sum_out[1][16][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][16][18] = (sum_out[2][16][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][16][18] = (sum_out[3][16][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][16][18] = (sum_out[4][16][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][16][18] = (sum_out[5][16][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][16][18] = (sum_out[6][16][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][16][18] = (sum_out[7][16][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][16][18] = (sum_out[8][16][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][16][18] = (sum_out[9][16][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][16][18] = (sum_out[10][16][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][16][18] = (sum_out[11][16][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][16][18] = (sum_out[12][16][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][16][18] = (sum_out[13][16][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][16][18] = (sum_out[14][16][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][16][18] = (sum_out[15][16][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][16][18] = (sum_out[16][16][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][16][18] = (sum_out[17][16][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][16][18] = (sum_out[18][16][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][16][18] = (sum_out[19][16][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][16][19] = (sum_out[0][16][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][16][19] = (sum_out[1][16][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][16][19] = (sum_out[2][16][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][16][19] = (sum_out[3][16][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][16][19] = (sum_out[4][16][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][16][19] = (sum_out[5][16][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][16][19] = (sum_out[6][16][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][16][19] = (sum_out[7][16][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][16][19] = (sum_out[8][16][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][16][19] = (sum_out[9][16][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][16][19] = (sum_out[10][16][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][16][19] = (sum_out[11][16][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][16][19] = (sum_out[12][16][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][16][19] = (sum_out[13][16][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][16][19] = (sum_out[14][16][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][16][19] = (sum_out[15][16][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][16][19] = (sum_out[16][16][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][16][19] = (sum_out[17][16][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][16][19] = (sum_out[18][16][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][16][19] = (sum_out[19][16][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][16][20] = (sum_out[0][16][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][16][20] = (sum_out[1][16][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][16][20] = (sum_out[2][16][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][16][20] = (sum_out[3][16][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][16][20] = (sum_out[4][16][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][16][20] = (sum_out[5][16][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][16][20] = (sum_out[6][16][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][16][20] = (sum_out[7][16][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][16][20] = (sum_out[8][16][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][16][20] = (sum_out[9][16][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][16][20] = (sum_out[10][16][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][16][20] = (sum_out[11][16][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][16][20] = (sum_out[12][16][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][16][20] = (sum_out[13][16][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][16][20] = (sum_out[14][16][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][16][20] = (sum_out[15][16][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][16][20] = (sum_out[16][16][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][16][20] = (sum_out[17][16][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][16][20] = (sum_out[18][16][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][16][20] = (sum_out[19][16][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][16][21] = (sum_out[0][16][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][16][21] = (sum_out[1][16][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][16][21] = (sum_out[2][16][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][16][21] = (sum_out[3][16][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][16][21] = (sum_out[4][16][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][16][21] = (sum_out[5][16][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][16][21] = (sum_out[6][16][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][16][21] = (sum_out[7][16][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][16][21] = (sum_out[8][16][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][16][21] = (sum_out[9][16][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][16][21] = (sum_out[10][16][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][16][21] = (sum_out[11][16][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][16][21] = (sum_out[12][16][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][16][21] = (sum_out[13][16][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][16][21] = (sum_out[14][16][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][16][21] = (sum_out[15][16][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][16][21] = (sum_out[16][16][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][16][21] = (sum_out[17][16][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][16][21] = (sum_out[18][16][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][16][21] = (sum_out[19][16][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][16][22] = (sum_out[0][16][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][16][22] = (sum_out[1][16][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][16][22] = (sum_out[2][16][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][16][22] = (sum_out[3][16][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][16][22] = (sum_out[4][16][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][16][22] = (sum_out[5][16][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][16][22] = (sum_out[6][16][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][16][22] = (sum_out[7][16][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][16][22] = (sum_out[8][16][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][16][22] = (sum_out[9][16][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][16][22] = (sum_out[10][16][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][16][22] = (sum_out[11][16][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][16][22] = (sum_out[12][16][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][16][22] = (sum_out[13][16][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][16][22] = (sum_out[14][16][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][16][22] = (sum_out[15][16][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][16][22] = (sum_out[16][16][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][16][22] = (sum_out[17][16][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][16][22] = (sum_out[18][16][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][16][22] = (sum_out[19][16][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][16][23] = (sum_out[0][16][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][16][23] = (sum_out[1][16][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][16][23] = (sum_out[2][16][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][16][23] = (sum_out[3][16][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][16][23] = (sum_out[4][16][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][16][23] = (sum_out[5][16][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][16][23] = (sum_out[6][16][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][16][23] = (sum_out[7][16][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][16][23] = (sum_out[8][16][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][16][23] = (sum_out[9][16][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][16][23] = (sum_out[10][16][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][16][23] = (sum_out[11][16][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][16][23] = (sum_out[12][16][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][16][23] = (sum_out[13][16][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][16][23] = (sum_out[14][16][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][16][23] = (sum_out[15][16][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][16][23] = (sum_out[16][16][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][16][23] = (sum_out[17][16][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][16][23] = (sum_out[18][16][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][16][23] = (sum_out[19][16][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][17][0] = (sum_out[0][17][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][17][0] = (sum_out[1][17][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][17][0] = (sum_out[2][17][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][17][0] = (sum_out[3][17][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][17][0] = (sum_out[4][17][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][17][0] = (sum_out[5][17][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][17][0] = (sum_out[6][17][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][17][0] = (sum_out[7][17][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][17][0] = (sum_out[8][17][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][17][0] = (sum_out[9][17][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][17][0] = (sum_out[10][17][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][17][0] = (sum_out[11][17][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][17][0] = (sum_out[12][17][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][17][0] = (sum_out[13][17][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][17][0] = (sum_out[14][17][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][17][0] = (sum_out[15][17][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][17][0] = (sum_out[16][17][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][17][0] = (sum_out[17][17][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][17][0] = (sum_out[18][17][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][17][0] = (sum_out[19][17][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][17][1] = (sum_out[0][17][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][17][1] = (sum_out[1][17][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][17][1] = (sum_out[2][17][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][17][1] = (sum_out[3][17][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][17][1] = (sum_out[4][17][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][17][1] = (sum_out[5][17][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][17][1] = (sum_out[6][17][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][17][1] = (sum_out[7][17][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][17][1] = (sum_out[8][17][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][17][1] = (sum_out[9][17][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][17][1] = (sum_out[10][17][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][17][1] = (sum_out[11][17][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][17][1] = (sum_out[12][17][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][17][1] = (sum_out[13][17][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][17][1] = (sum_out[14][17][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][17][1] = (sum_out[15][17][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][17][1] = (sum_out[16][17][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][17][1] = (sum_out[17][17][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][17][1] = (sum_out[18][17][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][17][1] = (sum_out[19][17][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][17][2] = (sum_out[0][17][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][17][2] = (sum_out[1][17][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][17][2] = (sum_out[2][17][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][17][2] = (sum_out[3][17][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][17][2] = (sum_out[4][17][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][17][2] = (sum_out[5][17][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][17][2] = (sum_out[6][17][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][17][2] = (sum_out[7][17][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][17][2] = (sum_out[8][17][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][17][2] = (sum_out[9][17][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][17][2] = (sum_out[10][17][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][17][2] = (sum_out[11][17][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][17][2] = (sum_out[12][17][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][17][2] = (sum_out[13][17][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][17][2] = (sum_out[14][17][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][17][2] = (sum_out[15][17][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][17][2] = (sum_out[16][17][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][17][2] = (sum_out[17][17][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][17][2] = (sum_out[18][17][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][17][2] = (sum_out[19][17][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][17][3] = (sum_out[0][17][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][17][3] = (sum_out[1][17][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][17][3] = (sum_out[2][17][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][17][3] = (sum_out[3][17][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][17][3] = (sum_out[4][17][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][17][3] = (sum_out[5][17][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][17][3] = (sum_out[6][17][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][17][3] = (sum_out[7][17][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][17][3] = (sum_out[8][17][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][17][3] = (sum_out[9][17][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][17][3] = (sum_out[10][17][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][17][3] = (sum_out[11][17][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][17][3] = (sum_out[12][17][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][17][3] = (sum_out[13][17][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][17][3] = (sum_out[14][17][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][17][3] = (sum_out[15][17][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][17][3] = (sum_out[16][17][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][17][3] = (sum_out[17][17][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][17][3] = (sum_out[18][17][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][17][3] = (sum_out[19][17][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][17][4] = (sum_out[0][17][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][17][4] = (sum_out[1][17][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][17][4] = (sum_out[2][17][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][17][4] = (sum_out[3][17][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][17][4] = (sum_out[4][17][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][17][4] = (sum_out[5][17][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][17][4] = (sum_out[6][17][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][17][4] = (sum_out[7][17][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][17][4] = (sum_out[8][17][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][17][4] = (sum_out[9][17][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][17][4] = (sum_out[10][17][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][17][4] = (sum_out[11][17][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][17][4] = (sum_out[12][17][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][17][4] = (sum_out[13][17][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][17][4] = (sum_out[14][17][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][17][4] = (sum_out[15][17][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][17][4] = (sum_out[16][17][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][17][4] = (sum_out[17][17][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][17][4] = (sum_out[18][17][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][17][4] = (sum_out[19][17][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][17][5] = (sum_out[0][17][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][17][5] = (sum_out[1][17][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][17][5] = (sum_out[2][17][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][17][5] = (sum_out[3][17][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][17][5] = (sum_out[4][17][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][17][5] = (sum_out[5][17][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][17][5] = (sum_out[6][17][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][17][5] = (sum_out[7][17][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][17][5] = (sum_out[8][17][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][17][5] = (sum_out[9][17][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][17][5] = (sum_out[10][17][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][17][5] = (sum_out[11][17][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][17][5] = (sum_out[12][17][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][17][5] = (sum_out[13][17][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][17][5] = (sum_out[14][17][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][17][5] = (sum_out[15][17][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][17][5] = (sum_out[16][17][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][17][5] = (sum_out[17][17][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][17][5] = (sum_out[18][17][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][17][5] = (sum_out[19][17][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][17][6] = (sum_out[0][17][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][17][6] = (sum_out[1][17][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][17][6] = (sum_out[2][17][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][17][6] = (sum_out[3][17][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][17][6] = (sum_out[4][17][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][17][6] = (sum_out[5][17][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][17][6] = (sum_out[6][17][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][17][6] = (sum_out[7][17][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][17][6] = (sum_out[8][17][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][17][6] = (sum_out[9][17][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][17][6] = (sum_out[10][17][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][17][6] = (sum_out[11][17][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][17][6] = (sum_out[12][17][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][17][6] = (sum_out[13][17][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][17][6] = (sum_out[14][17][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][17][6] = (sum_out[15][17][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][17][6] = (sum_out[16][17][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][17][6] = (sum_out[17][17][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][17][6] = (sum_out[18][17][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][17][6] = (sum_out[19][17][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][17][7] = (sum_out[0][17][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][17][7] = (sum_out[1][17][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][17][7] = (sum_out[2][17][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][17][7] = (sum_out[3][17][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][17][7] = (sum_out[4][17][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][17][7] = (sum_out[5][17][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][17][7] = (sum_out[6][17][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][17][7] = (sum_out[7][17][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][17][7] = (sum_out[8][17][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][17][7] = (sum_out[9][17][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][17][7] = (sum_out[10][17][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][17][7] = (sum_out[11][17][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][17][7] = (sum_out[12][17][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][17][7] = (sum_out[13][17][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][17][7] = (sum_out[14][17][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][17][7] = (sum_out[15][17][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][17][7] = (sum_out[16][17][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][17][7] = (sum_out[17][17][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][17][7] = (sum_out[18][17][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][17][7] = (sum_out[19][17][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][17][8] = (sum_out[0][17][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][17][8] = (sum_out[1][17][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][17][8] = (sum_out[2][17][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][17][8] = (sum_out[3][17][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][17][8] = (sum_out[4][17][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][17][8] = (sum_out[5][17][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][17][8] = (sum_out[6][17][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][17][8] = (sum_out[7][17][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][17][8] = (sum_out[8][17][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][17][8] = (sum_out[9][17][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][17][8] = (sum_out[10][17][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][17][8] = (sum_out[11][17][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][17][8] = (sum_out[12][17][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][17][8] = (sum_out[13][17][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][17][8] = (sum_out[14][17][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][17][8] = (sum_out[15][17][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][17][8] = (sum_out[16][17][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][17][8] = (sum_out[17][17][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][17][8] = (sum_out[18][17][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][17][8] = (sum_out[19][17][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][17][9] = (sum_out[0][17][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][17][9] = (sum_out[1][17][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][17][9] = (sum_out[2][17][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][17][9] = (sum_out[3][17][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][17][9] = (sum_out[4][17][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][17][9] = (sum_out[5][17][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][17][9] = (sum_out[6][17][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][17][9] = (sum_out[7][17][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][17][9] = (sum_out[8][17][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][17][9] = (sum_out[9][17][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][17][9] = (sum_out[10][17][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][17][9] = (sum_out[11][17][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][17][9] = (sum_out[12][17][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][17][9] = (sum_out[13][17][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][17][9] = (sum_out[14][17][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][17][9] = (sum_out[15][17][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][17][9] = (sum_out[16][17][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][17][9] = (sum_out[17][17][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][17][9] = (sum_out[18][17][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][17][9] = (sum_out[19][17][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][17][10] = (sum_out[0][17][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][17][10] = (sum_out[1][17][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][17][10] = (sum_out[2][17][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][17][10] = (sum_out[3][17][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][17][10] = (sum_out[4][17][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][17][10] = (sum_out[5][17][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][17][10] = (sum_out[6][17][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][17][10] = (sum_out[7][17][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][17][10] = (sum_out[8][17][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][17][10] = (sum_out[9][17][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][17][10] = (sum_out[10][17][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][17][10] = (sum_out[11][17][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][17][10] = (sum_out[12][17][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][17][10] = (sum_out[13][17][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][17][10] = (sum_out[14][17][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][17][10] = (sum_out[15][17][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][17][10] = (sum_out[16][17][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][17][10] = (sum_out[17][17][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][17][10] = (sum_out[18][17][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][17][10] = (sum_out[19][17][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][17][11] = (sum_out[0][17][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][17][11] = (sum_out[1][17][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][17][11] = (sum_out[2][17][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][17][11] = (sum_out[3][17][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][17][11] = (sum_out[4][17][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][17][11] = (sum_out[5][17][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][17][11] = (sum_out[6][17][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][17][11] = (sum_out[7][17][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][17][11] = (sum_out[8][17][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][17][11] = (sum_out[9][17][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][17][11] = (sum_out[10][17][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][17][11] = (sum_out[11][17][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][17][11] = (sum_out[12][17][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][17][11] = (sum_out[13][17][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][17][11] = (sum_out[14][17][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][17][11] = (sum_out[15][17][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][17][11] = (sum_out[16][17][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][17][11] = (sum_out[17][17][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][17][11] = (sum_out[18][17][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][17][11] = (sum_out[19][17][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][17][12] = (sum_out[0][17][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][17][12] = (sum_out[1][17][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][17][12] = (sum_out[2][17][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][17][12] = (sum_out[3][17][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][17][12] = (sum_out[4][17][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][17][12] = (sum_out[5][17][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][17][12] = (sum_out[6][17][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][17][12] = (sum_out[7][17][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][17][12] = (sum_out[8][17][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][17][12] = (sum_out[9][17][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][17][12] = (sum_out[10][17][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][17][12] = (sum_out[11][17][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][17][12] = (sum_out[12][17][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][17][12] = (sum_out[13][17][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][17][12] = (sum_out[14][17][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][17][12] = (sum_out[15][17][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][17][12] = (sum_out[16][17][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][17][12] = (sum_out[17][17][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][17][12] = (sum_out[18][17][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][17][12] = (sum_out[19][17][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][17][13] = (sum_out[0][17][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][17][13] = (sum_out[1][17][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][17][13] = (sum_out[2][17][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][17][13] = (sum_out[3][17][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][17][13] = (sum_out[4][17][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][17][13] = (sum_out[5][17][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][17][13] = (sum_out[6][17][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][17][13] = (sum_out[7][17][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][17][13] = (sum_out[8][17][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][17][13] = (sum_out[9][17][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][17][13] = (sum_out[10][17][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][17][13] = (sum_out[11][17][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][17][13] = (sum_out[12][17][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][17][13] = (sum_out[13][17][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][17][13] = (sum_out[14][17][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][17][13] = (sum_out[15][17][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][17][13] = (sum_out[16][17][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][17][13] = (sum_out[17][17][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][17][13] = (sum_out[18][17][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][17][13] = (sum_out[19][17][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][17][14] = (sum_out[0][17][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][17][14] = (sum_out[1][17][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][17][14] = (sum_out[2][17][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][17][14] = (sum_out[3][17][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][17][14] = (sum_out[4][17][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][17][14] = (sum_out[5][17][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][17][14] = (sum_out[6][17][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][17][14] = (sum_out[7][17][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][17][14] = (sum_out[8][17][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][17][14] = (sum_out[9][17][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][17][14] = (sum_out[10][17][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][17][14] = (sum_out[11][17][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][17][14] = (sum_out[12][17][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][17][14] = (sum_out[13][17][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][17][14] = (sum_out[14][17][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][17][14] = (sum_out[15][17][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][17][14] = (sum_out[16][17][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][17][14] = (sum_out[17][17][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][17][14] = (sum_out[18][17][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][17][14] = (sum_out[19][17][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][17][15] = (sum_out[0][17][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][17][15] = (sum_out[1][17][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][17][15] = (sum_out[2][17][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][17][15] = (sum_out[3][17][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][17][15] = (sum_out[4][17][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][17][15] = (sum_out[5][17][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][17][15] = (sum_out[6][17][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][17][15] = (sum_out[7][17][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][17][15] = (sum_out[8][17][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][17][15] = (sum_out[9][17][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][17][15] = (sum_out[10][17][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][17][15] = (sum_out[11][17][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][17][15] = (sum_out[12][17][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][17][15] = (sum_out[13][17][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][17][15] = (sum_out[14][17][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][17][15] = (sum_out[15][17][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][17][15] = (sum_out[16][17][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][17][15] = (sum_out[17][17][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][17][15] = (sum_out[18][17][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][17][15] = (sum_out[19][17][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][17][16] = (sum_out[0][17][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][17][16] = (sum_out[1][17][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][17][16] = (sum_out[2][17][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][17][16] = (sum_out[3][17][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][17][16] = (sum_out[4][17][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][17][16] = (sum_out[5][17][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][17][16] = (sum_out[6][17][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][17][16] = (sum_out[7][17][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][17][16] = (sum_out[8][17][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][17][16] = (sum_out[9][17][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][17][16] = (sum_out[10][17][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][17][16] = (sum_out[11][17][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][17][16] = (sum_out[12][17][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][17][16] = (sum_out[13][17][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][17][16] = (sum_out[14][17][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][17][16] = (sum_out[15][17][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][17][16] = (sum_out[16][17][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][17][16] = (sum_out[17][17][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][17][16] = (sum_out[18][17][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][17][16] = (sum_out[19][17][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][17][17] = (sum_out[0][17][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][17][17] = (sum_out[1][17][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][17][17] = (sum_out[2][17][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][17][17] = (sum_out[3][17][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][17][17] = (sum_out[4][17][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][17][17] = (sum_out[5][17][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][17][17] = (sum_out[6][17][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][17][17] = (sum_out[7][17][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][17][17] = (sum_out[8][17][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][17][17] = (sum_out[9][17][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][17][17] = (sum_out[10][17][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][17][17] = (sum_out[11][17][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][17][17] = (sum_out[12][17][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][17][17] = (sum_out[13][17][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][17][17] = (sum_out[14][17][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][17][17] = (sum_out[15][17][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][17][17] = (sum_out[16][17][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][17][17] = (sum_out[17][17][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][17][17] = (sum_out[18][17][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][17][17] = (sum_out[19][17][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][17][18] = (sum_out[0][17][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][17][18] = (sum_out[1][17][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][17][18] = (sum_out[2][17][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][17][18] = (sum_out[3][17][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][17][18] = (sum_out[4][17][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][17][18] = (sum_out[5][17][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][17][18] = (sum_out[6][17][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][17][18] = (sum_out[7][17][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][17][18] = (sum_out[8][17][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][17][18] = (sum_out[9][17][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][17][18] = (sum_out[10][17][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][17][18] = (sum_out[11][17][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][17][18] = (sum_out[12][17][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][17][18] = (sum_out[13][17][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][17][18] = (sum_out[14][17][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][17][18] = (sum_out[15][17][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][17][18] = (sum_out[16][17][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][17][18] = (sum_out[17][17][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][17][18] = (sum_out[18][17][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][17][18] = (sum_out[19][17][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][17][19] = (sum_out[0][17][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][17][19] = (sum_out[1][17][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][17][19] = (sum_out[2][17][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][17][19] = (sum_out[3][17][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][17][19] = (sum_out[4][17][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][17][19] = (sum_out[5][17][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][17][19] = (sum_out[6][17][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][17][19] = (sum_out[7][17][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][17][19] = (sum_out[8][17][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][17][19] = (sum_out[9][17][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][17][19] = (sum_out[10][17][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][17][19] = (sum_out[11][17][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][17][19] = (sum_out[12][17][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][17][19] = (sum_out[13][17][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][17][19] = (sum_out[14][17][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][17][19] = (sum_out[15][17][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][17][19] = (sum_out[16][17][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][17][19] = (sum_out[17][17][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][17][19] = (sum_out[18][17][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][17][19] = (sum_out[19][17][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][17][20] = (sum_out[0][17][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][17][20] = (sum_out[1][17][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][17][20] = (sum_out[2][17][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][17][20] = (sum_out[3][17][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][17][20] = (sum_out[4][17][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][17][20] = (sum_out[5][17][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][17][20] = (sum_out[6][17][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][17][20] = (sum_out[7][17][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][17][20] = (sum_out[8][17][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][17][20] = (sum_out[9][17][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][17][20] = (sum_out[10][17][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][17][20] = (sum_out[11][17][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][17][20] = (sum_out[12][17][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][17][20] = (sum_out[13][17][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][17][20] = (sum_out[14][17][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][17][20] = (sum_out[15][17][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][17][20] = (sum_out[16][17][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][17][20] = (sum_out[17][17][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][17][20] = (sum_out[18][17][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][17][20] = (sum_out[19][17][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][17][21] = (sum_out[0][17][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][17][21] = (sum_out[1][17][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][17][21] = (sum_out[2][17][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][17][21] = (sum_out[3][17][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][17][21] = (sum_out[4][17][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][17][21] = (sum_out[5][17][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][17][21] = (sum_out[6][17][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][17][21] = (sum_out[7][17][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][17][21] = (sum_out[8][17][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][17][21] = (sum_out[9][17][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][17][21] = (sum_out[10][17][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][17][21] = (sum_out[11][17][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][17][21] = (sum_out[12][17][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][17][21] = (sum_out[13][17][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][17][21] = (sum_out[14][17][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][17][21] = (sum_out[15][17][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][17][21] = (sum_out[16][17][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][17][21] = (sum_out[17][17][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][17][21] = (sum_out[18][17][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][17][21] = (sum_out[19][17][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][17][22] = (sum_out[0][17][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][17][22] = (sum_out[1][17][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][17][22] = (sum_out[2][17][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][17][22] = (sum_out[3][17][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][17][22] = (sum_out[4][17][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][17][22] = (sum_out[5][17][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][17][22] = (sum_out[6][17][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][17][22] = (sum_out[7][17][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][17][22] = (sum_out[8][17][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][17][22] = (sum_out[9][17][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][17][22] = (sum_out[10][17][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][17][22] = (sum_out[11][17][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][17][22] = (sum_out[12][17][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][17][22] = (sum_out[13][17][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][17][22] = (sum_out[14][17][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][17][22] = (sum_out[15][17][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][17][22] = (sum_out[16][17][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][17][22] = (sum_out[17][17][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][17][22] = (sum_out[18][17][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][17][22] = (sum_out[19][17][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][17][23] = (sum_out[0][17][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][17][23] = (sum_out[1][17][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][17][23] = (sum_out[2][17][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][17][23] = (sum_out[3][17][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][17][23] = (sum_out[4][17][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][17][23] = (sum_out[5][17][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][17][23] = (sum_out[6][17][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][17][23] = (sum_out[7][17][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][17][23] = (sum_out[8][17][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][17][23] = (sum_out[9][17][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][17][23] = (sum_out[10][17][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][17][23] = (sum_out[11][17][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][17][23] = (sum_out[12][17][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][17][23] = (sum_out[13][17][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][17][23] = (sum_out[14][17][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][17][23] = (sum_out[15][17][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][17][23] = (sum_out[16][17][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][17][23] = (sum_out[17][17][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][17][23] = (sum_out[18][17][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][17][23] = (sum_out[19][17][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][18][0] = (sum_out[0][18][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][18][0] = (sum_out[1][18][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][18][0] = (sum_out[2][18][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][18][0] = (sum_out[3][18][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][18][0] = (sum_out[4][18][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][18][0] = (sum_out[5][18][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][18][0] = (sum_out[6][18][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][18][0] = (sum_out[7][18][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][18][0] = (sum_out[8][18][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][18][0] = (sum_out[9][18][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][18][0] = (sum_out[10][18][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][18][0] = (sum_out[11][18][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][18][0] = (sum_out[12][18][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][18][0] = (sum_out[13][18][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][18][0] = (sum_out[14][18][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][18][0] = (sum_out[15][18][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][18][0] = (sum_out[16][18][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][18][0] = (sum_out[17][18][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][18][0] = (sum_out[18][18][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][18][0] = (sum_out[19][18][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][18][1] = (sum_out[0][18][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][18][1] = (sum_out[1][18][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][18][1] = (sum_out[2][18][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][18][1] = (sum_out[3][18][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][18][1] = (sum_out[4][18][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][18][1] = (sum_out[5][18][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][18][1] = (sum_out[6][18][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][18][1] = (sum_out[7][18][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][18][1] = (sum_out[8][18][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][18][1] = (sum_out[9][18][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][18][1] = (sum_out[10][18][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][18][1] = (sum_out[11][18][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][18][1] = (sum_out[12][18][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][18][1] = (sum_out[13][18][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][18][1] = (sum_out[14][18][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][18][1] = (sum_out[15][18][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][18][1] = (sum_out[16][18][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][18][1] = (sum_out[17][18][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][18][1] = (sum_out[18][18][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][18][1] = (sum_out[19][18][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][18][2] = (sum_out[0][18][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][18][2] = (sum_out[1][18][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][18][2] = (sum_out[2][18][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][18][2] = (sum_out[3][18][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][18][2] = (sum_out[4][18][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][18][2] = (sum_out[5][18][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][18][2] = (sum_out[6][18][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][18][2] = (sum_out[7][18][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][18][2] = (sum_out[8][18][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][18][2] = (sum_out[9][18][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][18][2] = (sum_out[10][18][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][18][2] = (sum_out[11][18][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][18][2] = (sum_out[12][18][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][18][2] = (sum_out[13][18][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][18][2] = (sum_out[14][18][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][18][2] = (sum_out[15][18][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][18][2] = (sum_out[16][18][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][18][2] = (sum_out[17][18][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][18][2] = (sum_out[18][18][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][18][2] = (sum_out[19][18][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][18][3] = (sum_out[0][18][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][18][3] = (sum_out[1][18][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][18][3] = (sum_out[2][18][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][18][3] = (sum_out[3][18][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][18][3] = (sum_out[4][18][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][18][3] = (sum_out[5][18][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][18][3] = (sum_out[6][18][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][18][3] = (sum_out[7][18][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][18][3] = (sum_out[8][18][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][18][3] = (sum_out[9][18][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][18][3] = (sum_out[10][18][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][18][3] = (sum_out[11][18][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][18][3] = (sum_out[12][18][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][18][3] = (sum_out[13][18][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][18][3] = (sum_out[14][18][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][18][3] = (sum_out[15][18][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][18][3] = (sum_out[16][18][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][18][3] = (sum_out[17][18][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][18][3] = (sum_out[18][18][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][18][3] = (sum_out[19][18][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][18][4] = (sum_out[0][18][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][18][4] = (sum_out[1][18][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][18][4] = (sum_out[2][18][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][18][4] = (sum_out[3][18][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][18][4] = (sum_out[4][18][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][18][4] = (sum_out[5][18][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][18][4] = (sum_out[6][18][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][18][4] = (sum_out[7][18][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][18][4] = (sum_out[8][18][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][18][4] = (sum_out[9][18][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][18][4] = (sum_out[10][18][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][18][4] = (sum_out[11][18][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][18][4] = (sum_out[12][18][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][18][4] = (sum_out[13][18][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][18][4] = (sum_out[14][18][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][18][4] = (sum_out[15][18][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][18][4] = (sum_out[16][18][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][18][4] = (sum_out[17][18][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][18][4] = (sum_out[18][18][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][18][4] = (sum_out[19][18][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][18][5] = (sum_out[0][18][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][18][5] = (sum_out[1][18][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][18][5] = (sum_out[2][18][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][18][5] = (sum_out[3][18][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][18][5] = (sum_out[4][18][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][18][5] = (sum_out[5][18][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][18][5] = (sum_out[6][18][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][18][5] = (sum_out[7][18][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][18][5] = (sum_out[8][18][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][18][5] = (sum_out[9][18][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][18][5] = (sum_out[10][18][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][18][5] = (sum_out[11][18][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][18][5] = (sum_out[12][18][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][18][5] = (sum_out[13][18][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][18][5] = (sum_out[14][18][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][18][5] = (sum_out[15][18][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][18][5] = (sum_out[16][18][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][18][5] = (sum_out[17][18][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][18][5] = (sum_out[18][18][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][18][5] = (sum_out[19][18][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][18][6] = (sum_out[0][18][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][18][6] = (sum_out[1][18][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][18][6] = (sum_out[2][18][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][18][6] = (sum_out[3][18][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][18][6] = (sum_out[4][18][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][18][6] = (sum_out[5][18][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][18][6] = (sum_out[6][18][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][18][6] = (sum_out[7][18][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][18][6] = (sum_out[8][18][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][18][6] = (sum_out[9][18][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][18][6] = (sum_out[10][18][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][18][6] = (sum_out[11][18][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][18][6] = (sum_out[12][18][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][18][6] = (sum_out[13][18][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][18][6] = (sum_out[14][18][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][18][6] = (sum_out[15][18][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][18][6] = (sum_out[16][18][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][18][6] = (sum_out[17][18][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][18][6] = (sum_out[18][18][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][18][6] = (sum_out[19][18][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][18][7] = (sum_out[0][18][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][18][7] = (sum_out[1][18][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][18][7] = (sum_out[2][18][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][18][7] = (sum_out[3][18][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][18][7] = (sum_out[4][18][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][18][7] = (sum_out[5][18][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][18][7] = (sum_out[6][18][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][18][7] = (sum_out[7][18][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][18][7] = (sum_out[8][18][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][18][7] = (sum_out[9][18][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][18][7] = (sum_out[10][18][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][18][7] = (sum_out[11][18][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][18][7] = (sum_out[12][18][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][18][7] = (sum_out[13][18][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][18][7] = (sum_out[14][18][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][18][7] = (sum_out[15][18][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][18][7] = (sum_out[16][18][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][18][7] = (sum_out[17][18][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][18][7] = (sum_out[18][18][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][18][7] = (sum_out[19][18][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][18][8] = (sum_out[0][18][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][18][8] = (sum_out[1][18][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][18][8] = (sum_out[2][18][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][18][8] = (sum_out[3][18][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][18][8] = (sum_out[4][18][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][18][8] = (sum_out[5][18][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][18][8] = (sum_out[6][18][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][18][8] = (sum_out[7][18][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][18][8] = (sum_out[8][18][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][18][8] = (sum_out[9][18][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][18][8] = (sum_out[10][18][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][18][8] = (sum_out[11][18][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][18][8] = (sum_out[12][18][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][18][8] = (sum_out[13][18][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][18][8] = (sum_out[14][18][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][18][8] = (sum_out[15][18][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][18][8] = (sum_out[16][18][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][18][8] = (sum_out[17][18][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][18][8] = (sum_out[18][18][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][18][8] = (sum_out[19][18][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][18][9] = (sum_out[0][18][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][18][9] = (sum_out[1][18][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][18][9] = (sum_out[2][18][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][18][9] = (sum_out[3][18][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][18][9] = (sum_out[4][18][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][18][9] = (sum_out[5][18][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][18][9] = (sum_out[6][18][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][18][9] = (sum_out[7][18][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][18][9] = (sum_out[8][18][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][18][9] = (sum_out[9][18][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][18][9] = (sum_out[10][18][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][18][9] = (sum_out[11][18][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][18][9] = (sum_out[12][18][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][18][9] = (sum_out[13][18][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][18][9] = (sum_out[14][18][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][18][9] = (sum_out[15][18][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][18][9] = (sum_out[16][18][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][18][9] = (sum_out[17][18][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][18][9] = (sum_out[18][18][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][18][9] = (sum_out[19][18][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][18][10] = (sum_out[0][18][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][18][10] = (sum_out[1][18][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][18][10] = (sum_out[2][18][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][18][10] = (sum_out[3][18][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][18][10] = (sum_out[4][18][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][18][10] = (sum_out[5][18][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][18][10] = (sum_out[6][18][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][18][10] = (sum_out[7][18][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][18][10] = (sum_out[8][18][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][18][10] = (sum_out[9][18][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][18][10] = (sum_out[10][18][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][18][10] = (sum_out[11][18][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][18][10] = (sum_out[12][18][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][18][10] = (sum_out[13][18][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][18][10] = (sum_out[14][18][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][18][10] = (sum_out[15][18][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][18][10] = (sum_out[16][18][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][18][10] = (sum_out[17][18][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][18][10] = (sum_out[18][18][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][18][10] = (sum_out[19][18][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][18][11] = (sum_out[0][18][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][18][11] = (sum_out[1][18][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][18][11] = (sum_out[2][18][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][18][11] = (sum_out[3][18][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][18][11] = (sum_out[4][18][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][18][11] = (sum_out[5][18][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][18][11] = (sum_out[6][18][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][18][11] = (sum_out[7][18][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][18][11] = (sum_out[8][18][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][18][11] = (sum_out[9][18][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][18][11] = (sum_out[10][18][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][18][11] = (sum_out[11][18][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][18][11] = (sum_out[12][18][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][18][11] = (sum_out[13][18][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][18][11] = (sum_out[14][18][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][18][11] = (sum_out[15][18][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][18][11] = (sum_out[16][18][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][18][11] = (sum_out[17][18][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][18][11] = (sum_out[18][18][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][18][11] = (sum_out[19][18][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][18][12] = (sum_out[0][18][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][18][12] = (sum_out[1][18][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][18][12] = (sum_out[2][18][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][18][12] = (sum_out[3][18][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][18][12] = (sum_out[4][18][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][18][12] = (sum_out[5][18][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][18][12] = (sum_out[6][18][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][18][12] = (sum_out[7][18][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][18][12] = (sum_out[8][18][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][18][12] = (sum_out[9][18][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][18][12] = (sum_out[10][18][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][18][12] = (sum_out[11][18][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][18][12] = (sum_out[12][18][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][18][12] = (sum_out[13][18][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][18][12] = (sum_out[14][18][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][18][12] = (sum_out[15][18][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][18][12] = (sum_out[16][18][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][18][12] = (sum_out[17][18][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][18][12] = (sum_out[18][18][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][18][12] = (sum_out[19][18][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][18][13] = (sum_out[0][18][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][18][13] = (sum_out[1][18][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][18][13] = (sum_out[2][18][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][18][13] = (sum_out[3][18][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][18][13] = (sum_out[4][18][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][18][13] = (sum_out[5][18][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][18][13] = (sum_out[6][18][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][18][13] = (sum_out[7][18][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][18][13] = (sum_out[8][18][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][18][13] = (sum_out[9][18][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][18][13] = (sum_out[10][18][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][18][13] = (sum_out[11][18][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][18][13] = (sum_out[12][18][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][18][13] = (sum_out[13][18][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][18][13] = (sum_out[14][18][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][18][13] = (sum_out[15][18][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][18][13] = (sum_out[16][18][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][18][13] = (sum_out[17][18][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][18][13] = (sum_out[18][18][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][18][13] = (sum_out[19][18][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][18][14] = (sum_out[0][18][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][18][14] = (sum_out[1][18][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][18][14] = (sum_out[2][18][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][18][14] = (sum_out[3][18][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][18][14] = (sum_out[4][18][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][18][14] = (sum_out[5][18][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][18][14] = (sum_out[6][18][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][18][14] = (sum_out[7][18][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][18][14] = (sum_out[8][18][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][18][14] = (sum_out[9][18][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][18][14] = (sum_out[10][18][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][18][14] = (sum_out[11][18][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][18][14] = (sum_out[12][18][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][18][14] = (sum_out[13][18][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][18][14] = (sum_out[14][18][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][18][14] = (sum_out[15][18][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][18][14] = (sum_out[16][18][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][18][14] = (sum_out[17][18][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][18][14] = (sum_out[18][18][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][18][14] = (sum_out[19][18][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][18][15] = (sum_out[0][18][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][18][15] = (sum_out[1][18][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][18][15] = (sum_out[2][18][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][18][15] = (sum_out[3][18][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][18][15] = (sum_out[4][18][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][18][15] = (sum_out[5][18][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][18][15] = (sum_out[6][18][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][18][15] = (sum_out[7][18][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][18][15] = (sum_out[8][18][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][18][15] = (sum_out[9][18][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][18][15] = (sum_out[10][18][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][18][15] = (sum_out[11][18][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][18][15] = (sum_out[12][18][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][18][15] = (sum_out[13][18][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][18][15] = (sum_out[14][18][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][18][15] = (sum_out[15][18][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][18][15] = (sum_out[16][18][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][18][15] = (sum_out[17][18][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][18][15] = (sum_out[18][18][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][18][15] = (sum_out[19][18][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][18][16] = (sum_out[0][18][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][18][16] = (sum_out[1][18][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][18][16] = (sum_out[2][18][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][18][16] = (sum_out[3][18][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][18][16] = (sum_out[4][18][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][18][16] = (sum_out[5][18][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][18][16] = (sum_out[6][18][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][18][16] = (sum_out[7][18][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][18][16] = (sum_out[8][18][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][18][16] = (sum_out[9][18][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][18][16] = (sum_out[10][18][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][18][16] = (sum_out[11][18][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][18][16] = (sum_out[12][18][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][18][16] = (sum_out[13][18][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][18][16] = (sum_out[14][18][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][18][16] = (sum_out[15][18][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][18][16] = (sum_out[16][18][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][18][16] = (sum_out[17][18][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][18][16] = (sum_out[18][18][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][18][16] = (sum_out[19][18][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][18][17] = (sum_out[0][18][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][18][17] = (sum_out[1][18][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][18][17] = (sum_out[2][18][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][18][17] = (sum_out[3][18][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][18][17] = (sum_out[4][18][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][18][17] = (sum_out[5][18][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][18][17] = (sum_out[6][18][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][18][17] = (sum_out[7][18][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][18][17] = (sum_out[8][18][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][18][17] = (sum_out[9][18][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][18][17] = (sum_out[10][18][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][18][17] = (sum_out[11][18][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][18][17] = (sum_out[12][18][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][18][17] = (sum_out[13][18][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][18][17] = (sum_out[14][18][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][18][17] = (sum_out[15][18][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][18][17] = (sum_out[16][18][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][18][17] = (sum_out[17][18][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][18][17] = (sum_out[18][18][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][18][17] = (sum_out[19][18][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][18][18] = (sum_out[0][18][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][18][18] = (sum_out[1][18][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][18][18] = (sum_out[2][18][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][18][18] = (sum_out[3][18][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][18][18] = (sum_out[4][18][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][18][18] = (sum_out[5][18][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][18][18] = (sum_out[6][18][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][18][18] = (sum_out[7][18][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][18][18] = (sum_out[8][18][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][18][18] = (sum_out[9][18][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][18][18] = (sum_out[10][18][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][18][18] = (sum_out[11][18][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][18][18] = (sum_out[12][18][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][18][18] = (sum_out[13][18][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][18][18] = (sum_out[14][18][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][18][18] = (sum_out[15][18][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][18][18] = (sum_out[16][18][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][18][18] = (sum_out[17][18][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][18][18] = (sum_out[18][18][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][18][18] = (sum_out[19][18][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][18][19] = (sum_out[0][18][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][18][19] = (sum_out[1][18][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][18][19] = (sum_out[2][18][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][18][19] = (sum_out[3][18][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][18][19] = (sum_out[4][18][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][18][19] = (sum_out[5][18][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][18][19] = (sum_out[6][18][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][18][19] = (sum_out[7][18][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][18][19] = (sum_out[8][18][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][18][19] = (sum_out[9][18][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][18][19] = (sum_out[10][18][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][18][19] = (sum_out[11][18][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][18][19] = (sum_out[12][18][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][18][19] = (sum_out[13][18][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][18][19] = (sum_out[14][18][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][18][19] = (sum_out[15][18][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][18][19] = (sum_out[16][18][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][18][19] = (sum_out[17][18][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][18][19] = (sum_out[18][18][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][18][19] = (sum_out[19][18][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][18][20] = (sum_out[0][18][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][18][20] = (sum_out[1][18][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][18][20] = (sum_out[2][18][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][18][20] = (sum_out[3][18][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][18][20] = (sum_out[4][18][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][18][20] = (sum_out[5][18][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][18][20] = (sum_out[6][18][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][18][20] = (sum_out[7][18][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][18][20] = (sum_out[8][18][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][18][20] = (sum_out[9][18][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][18][20] = (sum_out[10][18][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][18][20] = (sum_out[11][18][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][18][20] = (sum_out[12][18][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][18][20] = (sum_out[13][18][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][18][20] = (sum_out[14][18][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][18][20] = (sum_out[15][18][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][18][20] = (sum_out[16][18][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][18][20] = (sum_out[17][18][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][18][20] = (sum_out[18][18][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][18][20] = (sum_out[19][18][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][18][21] = (sum_out[0][18][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][18][21] = (sum_out[1][18][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][18][21] = (sum_out[2][18][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][18][21] = (sum_out[3][18][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][18][21] = (sum_out[4][18][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][18][21] = (sum_out[5][18][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][18][21] = (sum_out[6][18][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][18][21] = (sum_out[7][18][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][18][21] = (sum_out[8][18][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][18][21] = (sum_out[9][18][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][18][21] = (sum_out[10][18][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][18][21] = (sum_out[11][18][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][18][21] = (sum_out[12][18][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][18][21] = (sum_out[13][18][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][18][21] = (sum_out[14][18][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][18][21] = (sum_out[15][18][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][18][21] = (sum_out[16][18][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][18][21] = (sum_out[17][18][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][18][21] = (sum_out[18][18][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][18][21] = (sum_out[19][18][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][18][22] = (sum_out[0][18][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][18][22] = (sum_out[1][18][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][18][22] = (sum_out[2][18][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][18][22] = (sum_out[3][18][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][18][22] = (sum_out[4][18][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][18][22] = (sum_out[5][18][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][18][22] = (sum_out[6][18][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][18][22] = (sum_out[7][18][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][18][22] = (sum_out[8][18][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][18][22] = (sum_out[9][18][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][18][22] = (sum_out[10][18][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][18][22] = (sum_out[11][18][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][18][22] = (sum_out[12][18][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][18][22] = (sum_out[13][18][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][18][22] = (sum_out[14][18][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][18][22] = (sum_out[15][18][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][18][22] = (sum_out[16][18][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][18][22] = (sum_out[17][18][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][18][22] = (sum_out[18][18][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][18][22] = (sum_out[19][18][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][18][23] = (sum_out[0][18][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][18][23] = (sum_out[1][18][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][18][23] = (sum_out[2][18][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][18][23] = (sum_out[3][18][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][18][23] = (sum_out[4][18][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][18][23] = (sum_out[5][18][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][18][23] = (sum_out[6][18][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][18][23] = (sum_out[7][18][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][18][23] = (sum_out[8][18][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][18][23] = (sum_out[9][18][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][18][23] = (sum_out[10][18][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][18][23] = (sum_out[11][18][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][18][23] = (sum_out[12][18][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][18][23] = (sum_out[13][18][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][18][23] = (sum_out[14][18][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][18][23] = (sum_out[15][18][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][18][23] = (sum_out[16][18][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][18][23] = (sum_out[17][18][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][18][23] = (sum_out[18][18][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][18][23] = (sum_out[19][18][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][19][0] = (sum_out[0][19][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][19][0] = (sum_out[1][19][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][19][0] = (sum_out[2][19][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][19][0] = (sum_out[3][19][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][19][0] = (sum_out[4][19][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][19][0] = (sum_out[5][19][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][19][0] = (sum_out[6][19][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][19][0] = (sum_out[7][19][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][19][0] = (sum_out[8][19][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][19][0] = (sum_out[9][19][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][19][0] = (sum_out[10][19][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][19][0] = (sum_out[11][19][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][19][0] = (sum_out[12][19][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][19][0] = (sum_out[13][19][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][19][0] = (sum_out[14][19][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][19][0] = (sum_out[15][19][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][19][0] = (sum_out[16][19][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][19][0] = (sum_out[17][19][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][19][0] = (sum_out[18][19][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][19][0] = (sum_out[19][19][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][19][1] = (sum_out[0][19][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][19][1] = (sum_out[1][19][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][19][1] = (sum_out[2][19][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][19][1] = (sum_out[3][19][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][19][1] = (sum_out[4][19][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][19][1] = (sum_out[5][19][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][19][1] = (sum_out[6][19][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][19][1] = (sum_out[7][19][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][19][1] = (sum_out[8][19][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][19][1] = (sum_out[9][19][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][19][1] = (sum_out[10][19][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][19][1] = (sum_out[11][19][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][19][1] = (sum_out[12][19][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][19][1] = (sum_out[13][19][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][19][1] = (sum_out[14][19][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][19][1] = (sum_out[15][19][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][19][1] = (sum_out[16][19][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][19][1] = (sum_out[17][19][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][19][1] = (sum_out[18][19][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][19][1] = (sum_out[19][19][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][19][2] = (sum_out[0][19][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][19][2] = (sum_out[1][19][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][19][2] = (sum_out[2][19][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][19][2] = (sum_out[3][19][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][19][2] = (sum_out[4][19][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][19][2] = (sum_out[5][19][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][19][2] = (sum_out[6][19][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][19][2] = (sum_out[7][19][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][19][2] = (sum_out[8][19][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][19][2] = (sum_out[9][19][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][19][2] = (sum_out[10][19][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][19][2] = (sum_out[11][19][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][19][2] = (sum_out[12][19][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][19][2] = (sum_out[13][19][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][19][2] = (sum_out[14][19][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][19][2] = (sum_out[15][19][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][19][2] = (sum_out[16][19][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][19][2] = (sum_out[17][19][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][19][2] = (sum_out[18][19][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][19][2] = (sum_out[19][19][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][19][3] = (sum_out[0][19][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][19][3] = (sum_out[1][19][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][19][3] = (sum_out[2][19][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][19][3] = (sum_out[3][19][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][19][3] = (sum_out[4][19][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][19][3] = (sum_out[5][19][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][19][3] = (sum_out[6][19][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][19][3] = (sum_out[7][19][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][19][3] = (sum_out[8][19][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][19][3] = (sum_out[9][19][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][19][3] = (sum_out[10][19][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][19][3] = (sum_out[11][19][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][19][3] = (sum_out[12][19][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][19][3] = (sum_out[13][19][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][19][3] = (sum_out[14][19][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][19][3] = (sum_out[15][19][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][19][3] = (sum_out[16][19][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][19][3] = (sum_out[17][19][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][19][3] = (sum_out[18][19][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][19][3] = (sum_out[19][19][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][19][4] = (sum_out[0][19][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][19][4] = (sum_out[1][19][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][19][4] = (sum_out[2][19][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][19][4] = (sum_out[3][19][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][19][4] = (sum_out[4][19][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][19][4] = (sum_out[5][19][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][19][4] = (sum_out[6][19][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][19][4] = (sum_out[7][19][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][19][4] = (sum_out[8][19][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][19][4] = (sum_out[9][19][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][19][4] = (sum_out[10][19][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][19][4] = (sum_out[11][19][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][19][4] = (sum_out[12][19][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][19][4] = (sum_out[13][19][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][19][4] = (sum_out[14][19][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][19][4] = (sum_out[15][19][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][19][4] = (sum_out[16][19][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][19][4] = (sum_out[17][19][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][19][4] = (sum_out[18][19][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][19][4] = (sum_out[19][19][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][19][5] = (sum_out[0][19][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][19][5] = (sum_out[1][19][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][19][5] = (sum_out[2][19][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][19][5] = (sum_out[3][19][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][19][5] = (sum_out[4][19][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][19][5] = (sum_out[5][19][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][19][5] = (sum_out[6][19][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][19][5] = (sum_out[7][19][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][19][5] = (sum_out[8][19][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][19][5] = (sum_out[9][19][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][19][5] = (sum_out[10][19][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][19][5] = (sum_out[11][19][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][19][5] = (sum_out[12][19][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][19][5] = (sum_out[13][19][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][19][5] = (sum_out[14][19][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][19][5] = (sum_out[15][19][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][19][5] = (sum_out[16][19][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][19][5] = (sum_out[17][19][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][19][5] = (sum_out[18][19][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][19][5] = (sum_out[19][19][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][19][6] = (sum_out[0][19][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][19][6] = (sum_out[1][19][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][19][6] = (sum_out[2][19][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][19][6] = (sum_out[3][19][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][19][6] = (sum_out[4][19][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][19][6] = (sum_out[5][19][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][19][6] = (sum_out[6][19][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][19][6] = (sum_out[7][19][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][19][6] = (sum_out[8][19][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][19][6] = (sum_out[9][19][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][19][6] = (sum_out[10][19][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][19][6] = (sum_out[11][19][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][19][6] = (sum_out[12][19][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][19][6] = (sum_out[13][19][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][19][6] = (sum_out[14][19][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][19][6] = (sum_out[15][19][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][19][6] = (sum_out[16][19][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][19][6] = (sum_out[17][19][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][19][6] = (sum_out[18][19][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][19][6] = (sum_out[19][19][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][19][7] = (sum_out[0][19][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][19][7] = (sum_out[1][19][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][19][7] = (sum_out[2][19][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][19][7] = (sum_out[3][19][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][19][7] = (sum_out[4][19][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][19][7] = (sum_out[5][19][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][19][7] = (sum_out[6][19][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][19][7] = (sum_out[7][19][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][19][7] = (sum_out[8][19][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][19][7] = (sum_out[9][19][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][19][7] = (sum_out[10][19][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][19][7] = (sum_out[11][19][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][19][7] = (sum_out[12][19][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][19][7] = (sum_out[13][19][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][19][7] = (sum_out[14][19][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][19][7] = (sum_out[15][19][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][19][7] = (sum_out[16][19][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][19][7] = (sum_out[17][19][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][19][7] = (sum_out[18][19][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][19][7] = (sum_out[19][19][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][19][8] = (sum_out[0][19][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][19][8] = (sum_out[1][19][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][19][8] = (sum_out[2][19][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][19][8] = (sum_out[3][19][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][19][8] = (sum_out[4][19][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][19][8] = (sum_out[5][19][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][19][8] = (sum_out[6][19][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][19][8] = (sum_out[7][19][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][19][8] = (sum_out[8][19][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][19][8] = (sum_out[9][19][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][19][8] = (sum_out[10][19][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][19][8] = (sum_out[11][19][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][19][8] = (sum_out[12][19][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][19][8] = (sum_out[13][19][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][19][8] = (sum_out[14][19][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][19][8] = (sum_out[15][19][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][19][8] = (sum_out[16][19][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][19][8] = (sum_out[17][19][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][19][8] = (sum_out[18][19][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][19][8] = (sum_out[19][19][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][19][9] = (sum_out[0][19][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][19][9] = (sum_out[1][19][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][19][9] = (sum_out[2][19][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][19][9] = (sum_out[3][19][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][19][9] = (sum_out[4][19][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][19][9] = (sum_out[5][19][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][19][9] = (sum_out[6][19][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][19][9] = (sum_out[7][19][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][19][9] = (sum_out[8][19][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][19][9] = (sum_out[9][19][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][19][9] = (sum_out[10][19][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][19][9] = (sum_out[11][19][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][19][9] = (sum_out[12][19][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][19][9] = (sum_out[13][19][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][19][9] = (sum_out[14][19][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][19][9] = (sum_out[15][19][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][19][9] = (sum_out[16][19][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][19][9] = (sum_out[17][19][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][19][9] = (sum_out[18][19][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][19][9] = (sum_out[19][19][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][19][10] = (sum_out[0][19][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][19][10] = (sum_out[1][19][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][19][10] = (sum_out[2][19][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][19][10] = (sum_out[3][19][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][19][10] = (sum_out[4][19][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][19][10] = (sum_out[5][19][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][19][10] = (sum_out[6][19][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][19][10] = (sum_out[7][19][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][19][10] = (sum_out[8][19][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][19][10] = (sum_out[9][19][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][19][10] = (sum_out[10][19][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][19][10] = (sum_out[11][19][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][19][10] = (sum_out[12][19][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][19][10] = (sum_out[13][19][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][19][10] = (sum_out[14][19][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][19][10] = (sum_out[15][19][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][19][10] = (sum_out[16][19][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][19][10] = (sum_out[17][19][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][19][10] = (sum_out[18][19][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][19][10] = (sum_out[19][19][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][19][11] = (sum_out[0][19][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][19][11] = (sum_out[1][19][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][19][11] = (sum_out[2][19][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][19][11] = (sum_out[3][19][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][19][11] = (sum_out[4][19][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][19][11] = (sum_out[5][19][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][19][11] = (sum_out[6][19][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][19][11] = (sum_out[7][19][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][19][11] = (sum_out[8][19][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][19][11] = (sum_out[9][19][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][19][11] = (sum_out[10][19][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][19][11] = (sum_out[11][19][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][19][11] = (sum_out[12][19][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][19][11] = (sum_out[13][19][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][19][11] = (sum_out[14][19][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][19][11] = (sum_out[15][19][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][19][11] = (sum_out[16][19][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][19][11] = (sum_out[17][19][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][19][11] = (sum_out[18][19][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][19][11] = (sum_out[19][19][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][19][12] = (sum_out[0][19][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][19][12] = (sum_out[1][19][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][19][12] = (sum_out[2][19][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][19][12] = (sum_out[3][19][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][19][12] = (sum_out[4][19][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][19][12] = (sum_out[5][19][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][19][12] = (sum_out[6][19][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][19][12] = (sum_out[7][19][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][19][12] = (sum_out[8][19][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][19][12] = (sum_out[9][19][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][19][12] = (sum_out[10][19][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][19][12] = (sum_out[11][19][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][19][12] = (sum_out[12][19][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][19][12] = (sum_out[13][19][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][19][12] = (sum_out[14][19][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][19][12] = (sum_out[15][19][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][19][12] = (sum_out[16][19][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][19][12] = (sum_out[17][19][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][19][12] = (sum_out[18][19][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][19][12] = (sum_out[19][19][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][19][13] = (sum_out[0][19][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][19][13] = (sum_out[1][19][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][19][13] = (sum_out[2][19][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][19][13] = (sum_out[3][19][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][19][13] = (sum_out[4][19][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][19][13] = (sum_out[5][19][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][19][13] = (sum_out[6][19][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][19][13] = (sum_out[7][19][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][19][13] = (sum_out[8][19][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][19][13] = (sum_out[9][19][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][19][13] = (sum_out[10][19][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][19][13] = (sum_out[11][19][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][19][13] = (sum_out[12][19][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][19][13] = (sum_out[13][19][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][19][13] = (sum_out[14][19][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][19][13] = (sum_out[15][19][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][19][13] = (sum_out[16][19][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][19][13] = (sum_out[17][19][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][19][13] = (sum_out[18][19][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][19][13] = (sum_out[19][19][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][19][14] = (sum_out[0][19][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][19][14] = (sum_out[1][19][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][19][14] = (sum_out[2][19][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][19][14] = (sum_out[3][19][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][19][14] = (sum_out[4][19][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][19][14] = (sum_out[5][19][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][19][14] = (sum_out[6][19][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][19][14] = (sum_out[7][19][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][19][14] = (sum_out[8][19][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][19][14] = (sum_out[9][19][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][19][14] = (sum_out[10][19][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][19][14] = (sum_out[11][19][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][19][14] = (sum_out[12][19][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][19][14] = (sum_out[13][19][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][19][14] = (sum_out[14][19][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][19][14] = (sum_out[15][19][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][19][14] = (sum_out[16][19][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][19][14] = (sum_out[17][19][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][19][14] = (sum_out[18][19][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][19][14] = (sum_out[19][19][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][19][15] = (sum_out[0][19][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][19][15] = (sum_out[1][19][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][19][15] = (sum_out[2][19][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][19][15] = (sum_out[3][19][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][19][15] = (sum_out[4][19][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][19][15] = (sum_out[5][19][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][19][15] = (sum_out[6][19][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][19][15] = (sum_out[7][19][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][19][15] = (sum_out[8][19][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][19][15] = (sum_out[9][19][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][19][15] = (sum_out[10][19][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][19][15] = (sum_out[11][19][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][19][15] = (sum_out[12][19][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][19][15] = (sum_out[13][19][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][19][15] = (sum_out[14][19][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][19][15] = (sum_out[15][19][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][19][15] = (sum_out[16][19][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][19][15] = (sum_out[17][19][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][19][15] = (sum_out[18][19][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][19][15] = (sum_out[19][19][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][19][16] = (sum_out[0][19][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][19][16] = (sum_out[1][19][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][19][16] = (sum_out[2][19][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][19][16] = (sum_out[3][19][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][19][16] = (sum_out[4][19][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][19][16] = (sum_out[5][19][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][19][16] = (sum_out[6][19][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][19][16] = (sum_out[7][19][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][19][16] = (sum_out[8][19][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][19][16] = (sum_out[9][19][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][19][16] = (sum_out[10][19][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][19][16] = (sum_out[11][19][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][19][16] = (sum_out[12][19][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][19][16] = (sum_out[13][19][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][19][16] = (sum_out[14][19][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][19][16] = (sum_out[15][19][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][19][16] = (sum_out[16][19][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][19][16] = (sum_out[17][19][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][19][16] = (sum_out[18][19][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][19][16] = (sum_out[19][19][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][19][17] = (sum_out[0][19][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][19][17] = (sum_out[1][19][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][19][17] = (sum_out[2][19][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][19][17] = (sum_out[3][19][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][19][17] = (sum_out[4][19][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][19][17] = (sum_out[5][19][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][19][17] = (sum_out[6][19][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][19][17] = (sum_out[7][19][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][19][17] = (sum_out[8][19][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][19][17] = (sum_out[9][19][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][19][17] = (sum_out[10][19][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][19][17] = (sum_out[11][19][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][19][17] = (sum_out[12][19][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][19][17] = (sum_out[13][19][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][19][17] = (sum_out[14][19][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][19][17] = (sum_out[15][19][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][19][17] = (sum_out[16][19][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][19][17] = (sum_out[17][19][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][19][17] = (sum_out[18][19][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][19][17] = (sum_out[19][19][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][19][18] = (sum_out[0][19][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][19][18] = (sum_out[1][19][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][19][18] = (sum_out[2][19][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][19][18] = (sum_out[3][19][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][19][18] = (sum_out[4][19][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][19][18] = (sum_out[5][19][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][19][18] = (sum_out[6][19][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][19][18] = (sum_out[7][19][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][19][18] = (sum_out[8][19][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][19][18] = (sum_out[9][19][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][19][18] = (sum_out[10][19][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][19][18] = (sum_out[11][19][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][19][18] = (sum_out[12][19][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][19][18] = (sum_out[13][19][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][19][18] = (sum_out[14][19][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][19][18] = (sum_out[15][19][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][19][18] = (sum_out[16][19][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][19][18] = (sum_out[17][19][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][19][18] = (sum_out[18][19][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][19][18] = (sum_out[19][19][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][19][19] = (sum_out[0][19][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][19][19] = (sum_out[1][19][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][19][19] = (sum_out[2][19][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][19][19] = (sum_out[3][19][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][19][19] = (sum_out[4][19][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][19][19] = (sum_out[5][19][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][19][19] = (sum_out[6][19][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][19][19] = (sum_out[7][19][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][19][19] = (sum_out[8][19][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][19][19] = (sum_out[9][19][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][19][19] = (sum_out[10][19][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][19][19] = (sum_out[11][19][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][19][19] = (sum_out[12][19][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][19][19] = (sum_out[13][19][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][19][19] = (sum_out[14][19][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][19][19] = (sum_out[15][19][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][19][19] = (sum_out[16][19][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][19][19] = (sum_out[17][19][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][19][19] = (sum_out[18][19][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][19][19] = (sum_out[19][19][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][19][20] = (sum_out[0][19][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][19][20] = (sum_out[1][19][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][19][20] = (sum_out[2][19][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][19][20] = (sum_out[3][19][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][19][20] = (sum_out[4][19][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][19][20] = (sum_out[5][19][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][19][20] = (sum_out[6][19][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][19][20] = (sum_out[7][19][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][19][20] = (sum_out[8][19][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][19][20] = (sum_out[9][19][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][19][20] = (sum_out[10][19][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][19][20] = (sum_out[11][19][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][19][20] = (sum_out[12][19][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][19][20] = (sum_out[13][19][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][19][20] = (sum_out[14][19][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][19][20] = (sum_out[15][19][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][19][20] = (sum_out[16][19][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][19][20] = (sum_out[17][19][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][19][20] = (sum_out[18][19][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][19][20] = (sum_out[19][19][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][19][21] = (sum_out[0][19][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][19][21] = (sum_out[1][19][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][19][21] = (sum_out[2][19][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][19][21] = (sum_out[3][19][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][19][21] = (sum_out[4][19][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][19][21] = (sum_out[5][19][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][19][21] = (sum_out[6][19][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][19][21] = (sum_out[7][19][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][19][21] = (sum_out[8][19][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][19][21] = (sum_out[9][19][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][19][21] = (sum_out[10][19][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][19][21] = (sum_out[11][19][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][19][21] = (sum_out[12][19][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][19][21] = (sum_out[13][19][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][19][21] = (sum_out[14][19][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][19][21] = (sum_out[15][19][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][19][21] = (sum_out[16][19][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][19][21] = (sum_out[17][19][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][19][21] = (sum_out[18][19][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][19][21] = (sum_out[19][19][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][19][22] = (sum_out[0][19][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][19][22] = (sum_out[1][19][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][19][22] = (sum_out[2][19][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][19][22] = (sum_out[3][19][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][19][22] = (sum_out[4][19][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][19][22] = (sum_out[5][19][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][19][22] = (sum_out[6][19][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][19][22] = (sum_out[7][19][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][19][22] = (sum_out[8][19][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][19][22] = (sum_out[9][19][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][19][22] = (sum_out[10][19][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][19][22] = (sum_out[11][19][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][19][22] = (sum_out[12][19][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][19][22] = (sum_out[13][19][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][19][22] = (sum_out[14][19][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][19][22] = (sum_out[15][19][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][19][22] = (sum_out[16][19][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][19][22] = (sum_out[17][19][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][19][22] = (sum_out[18][19][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][19][22] = (sum_out[19][19][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][19][23] = (sum_out[0][19][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][19][23] = (sum_out[1][19][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][19][23] = (sum_out[2][19][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][19][23] = (sum_out[3][19][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][19][23] = (sum_out[4][19][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][19][23] = (sum_out[5][19][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][19][23] = (sum_out[6][19][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][19][23] = (sum_out[7][19][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][19][23] = (sum_out[8][19][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][19][23] = (sum_out[9][19][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][19][23] = (sum_out[10][19][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][19][23] = (sum_out[11][19][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][19][23] = (sum_out[12][19][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][19][23] = (sum_out[13][19][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][19][23] = (sum_out[14][19][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][19][23] = (sum_out[15][19][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][19][23] = (sum_out[16][19][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][19][23] = (sum_out[17][19][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][19][23] = (sum_out[18][19][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][19][23] = (sum_out[19][19][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][20][0] = (sum_out[0][20][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][20][0] = (sum_out[1][20][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][20][0] = (sum_out[2][20][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][20][0] = (sum_out[3][20][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][20][0] = (sum_out[4][20][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][20][0] = (sum_out[5][20][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][20][0] = (sum_out[6][20][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][20][0] = (sum_out[7][20][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][20][0] = (sum_out[8][20][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][20][0] = (sum_out[9][20][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][20][0] = (sum_out[10][20][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][20][0] = (sum_out[11][20][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][20][0] = (sum_out[12][20][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][20][0] = (sum_out[13][20][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][20][0] = (sum_out[14][20][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][20][0] = (sum_out[15][20][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][20][0] = (sum_out[16][20][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][20][0] = (sum_out[17][20][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][20][0] = (sum_out[18][20][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][20][0] = (sum_out[19][20][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][20][1] = (sum_out[0][20][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][20][1] = (sum_out[1][20][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][20][1] = (sum_out[2][20][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][20][1] = (sum_out[3][20][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][20][1] = (sum_out[4][20][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][20][1] = (sum_out[5][20][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][20][1] = (sum_out[6][20][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][20][1] = (sum_out[7][20][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][20][1] = (sum_out[8][20][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][20][1] = (sum_out[9][20][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][20][1] = (sum_out[10][20][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][20][1] = (sum_out[11][20][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][20][1] = (sum_out[12][20][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][20][1] = (sum_out[13][20][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][20][1] = (sum_out[14][20][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][20][1] = (sum_out[15][20][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][20][1] = (sum_out[16][20][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][20][1] = (sum_out[17][20][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][20][1] = (sum_out[18][20][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][20][1] = (sum_out[19][20][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][20][2] = (sum_out[0][20][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][20][2] = (sum_out[1][20][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][20][2] = (sum_out[2][20][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][20][2] = (sum_out[3][20][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][20][2] = (sum_out[4][20][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][20][2] = (sum_out[5][20][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][20][2] = (sum_out[6][20][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][20][2] = (sum_out[7][20][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][20][2] = (sum_out[8][20][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][20][2] = (sum_out[9][20][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][20][2] = (sum_out[10][20][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][20][2] = (sum_out[11][20][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][20][2] = (sum_out[12][20][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][20][2] = (sum_out[13][20][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][20][2] = (sum_out[14][20][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][20][2] = (sum_out[15][20][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][20][2] = (sum_out[16][20][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][20][2] = (sum_out[17][20][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][20][2] = (sum_out[18][20][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][20][2] = (sum_out[19][20][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][20][3] = (sum_out[0][20][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][20][3] = (sum_out[1][20][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][20][3] = (sum_out[2][20][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][20][3] = (sum_out[3][20][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][20][3] = (sum_out[4][20][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][20][3] = (sum_out[5][20][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][20][3] = (sum_out[6][20][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][20][3] = (sum_out[7][20][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][20][3] = (sum_out[8][20][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][20][3] = (sum_out[9][20][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][20][3] = (sum_out[10][20][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][20][3] = (sum_out[11][20][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][20][3] = (sum_out[12][20][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][20][3] = (sum_out[13][20][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][20][3] = (sum_out[14][20][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][20][3] = (sum_out[15][20][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][20][3] = (sum_out[16][20][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][20][3] = (sum_out[17][20][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][20][3] = (sum_out[18][20][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][20][3] = (sum_out[19][20][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][20][4] = (sum_out[0][20][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][20][4] = (sum_out[1][20][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][20][4] = (sum_out[2][20][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][20][4] = (sum_out[3][20][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][20][4] = (sum_out[4][20][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][20][4] = (sum_out[5][20][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][20][4] = (sum_out[6][20][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][20][4] = (sum_out[7][20][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][20][4] = (sum_out[8][20][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][20][4] = (sum_out[9][20][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][20][4] = (sum_out[10][20][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][20][4] = (sum_out[11][20][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][20][4] = (sum_out[12][20][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][20][4] = (sum_out[13][20][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][20][4] = (sum_out[14][20][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][20][4] = (sum_out[15][20][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][20][4] = (sum_out[16][20][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][20][4] = (sum_out[17][20][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][20][4] = (sum_out[18][20][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][20][4] = (sum_out[19][20][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][20][5] = (sum_out[0][20][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][20][5] = (sum_out[1][20][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][20][5] = (sum_out[2][20][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][20][5] = (sum_out[3][20][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][20][5] = (sum_out[4][20][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][20][5] = (sum_out[5][20][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][20][5] = (sum_out[6][20][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][20][5] = (sum_out[7][20][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][20][5] = (sum_out[8][20][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][20][5] = (sum_out[9][20][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][20][5] = (sum_out[10][20][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][20][5] = (sum_out[11][20][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][20][5] = (sum_out[12][20][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][20][5] = (sum_out[13][20][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][20][5] = (sum_out[14][20][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][20][5] = (sum_out[15][20][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][20][5] = (sum_out[16][20][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][20][5] = (sum_out[17][20][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][20][5] = (sum_out[18][20][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][20][5] = (sum_out[19][20][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][20][6] = (sum_out[0][20][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][20][6] = (sum_out[1][20][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][20][6] = (sum_out[2][20][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][20][6] = (sum_out[3][20][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][20][6] = (sum_out[4][20][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][20][6] = (sum_out[5][20][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][20][6] = (sum_out[6][20][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][20][6] = (sum_out[7][20][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][20][6] = (sum_out[8][20][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][20][6] = (sum_out[9][20][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][20][6] = (sum_out[10][20][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][20][6] = (sum_out[11][20][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][20][6] = (sum_out[12][20][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][20][6] = (sum_out[13][20][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][20][6] = (sum_out[14][20][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][20][6] = (sum_out[15][20][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][20][6] = (sum_out[16][20][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][20][6] = (sum_out[17][20][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][20][6] = (sum_out[18][20][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][20][6] = (sum_out[19][20][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][20][7] = (sum_out[0][20][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][20][7] = (sum_out[1][20][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][20][7] = (sum_out[2][20][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][20][7] = (sum_out[3][20][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][20][7] = (sum_out[4][20][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][20][7] = (sum_out[5][20][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][20][7] = (sum_out[6][20][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][20][7] = (sum_out[7][20][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][20][7] = (sum_out[8][20][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][20][7] = (sum_out[9][20][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][20][7] = (sum_out[10][20][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][20][7] = (sum_out[11][20][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][20][7] = (sum_out[12][20][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][20][7] = (sum_out[13][20][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][20][7] = (sum_out[14][20][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][20][7] = (sum_out[15][20][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][20][7] = (sum_out[16][20][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][20][7] = (sum_out[17][20][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][20][7] = (sum_out[18][20][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][20][7] = (sum_out[19][20][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][20][8] = (sum_out[0][20][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][20][8] = (sum_out[1][20][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][20][8] = (sum_out[2][20][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][20][8] = (sum_out[3][20][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][20][8] = (sum_out[4][20][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][20][8] = (sum_out[5][20][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][20][8] = (sum_out[6][20][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][20][8] = (sum_out[7][20][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][20][8] = (sum_out[8][20][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][20][8] = (sum_out[9][20][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][20][8] = (sum_out[10][20][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][20][8] = (sum_out[11][20][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][20][8] = (sum_out[12][20][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][20][8] = (sum_out[13][20][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][20][8] = (sum_out[14][20][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][20][8] = (sum_out[15][20][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][20][8] = (sum_out[16][20][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][20][8] = (sum_out[17][20][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][20][8] = (sum_out[18][20][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][20][8] = (sum_out[19][20][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][20][9] = (sum_out[0][20][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][20][9] = (sum_out[1][20][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][20][9] = (sum_out[2][20][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][20][9] = (sum_out[3][20][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][20][9] = (sum_out[4][20][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][20][9] = (sum_out[5][20][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][20][9] = (sum_out[6][20][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][20][9] = (sum_out[7][20][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][20][9] = (sum_out[8][20][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][20][9] = (sum_out[9][20][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][20][9] = (sum_out[10][20][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][20][9] = (sum_out[11][20][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][20][9] = (sum_out[12][20][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][20][9] = (sum_out[13][20][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][20][9] = (sum_out[14][20][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][20][9] = (sum_out[15][20][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][20][9] = (sum_out[16][20][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][20][9] = (sum_out[17][20][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][20][9] = (sum_out[18][20][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][20][9] = (sum_out[19][20][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][20][10] = (sum_out[0][20][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][20][10] = (sum_out[1][20][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][20][10] = (sum_out[2][20][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][20][10] = (sum_out[3][20][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][20][10] = (sum_out[4][20][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][20][10] = (sum_out[5][20][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][20][10] = (sum_out[6][20][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][20][10] = (sum_out[7][20][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][20][10] = (sum_out[8][20][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][20][10] = (sum_out[9][20][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][20][10] = (sum_out[10][20][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][20][10] = (sum_out[11][20][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][20][10] = (sum_out[12][20][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][20][10] = (sum_out[13][20][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][20][10] = (sum_out[14][20][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][20][10] = (sum_out[15][20][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][20][10] = (sum_out[16][20][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][20][10] = (sum_out[17][20][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][20][10] = (sum_out[18][20][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][20][10] = (sum_out[19][20][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][20][11] = (sum_out[0][20][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][20][11] = (sum_out[1][20][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][20][11] = (sum_out[2][20][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][20][11] = (sum_out[3][20][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][20][11] = (sum_out[4][20][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][20][11] = (sum_out[5][20][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][20][11] = (sum_out[6][20][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][20][11] = (sum_out[7][20][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][20][11] = (sum_out[8][20][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][20][11] = (sum_out[9][20][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][20][11] = (sum_out[10][20][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][20][11] = (sum_out[11][20][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][20][11] = (sum_out[12][20][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][20][11] = (sum_out[13][20][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][20][11] = (sum_out[14][20][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][20][11] = (sum_out[15][20][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][20][11] = (sum_out[16][20][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][20][11] = (sum_out[17][20][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][20][11] = (sum_out[18][20][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][20][11] = (sum_out[19][20][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][20][12] = (sum_out[0][20][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][20][12] = (sum_out[1][20][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][20][12] = (sum_out[2][20][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][20][12] = (sum_out[3][20][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][20][12] = (sum_out[4][20][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][20][12] = (sum_out[5][20][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][20][12] = (sum_out[6][20][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][20][12] = (sum_out[7][20][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][20][12] = (sum_out[8][20][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][20][12] = (sum_out[9][20][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][20][12] = (sum_out[10][20][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][20][12] = (sum_out[11][20][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][20][12] = (sum_out[12][20][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][20][12] = (sum_out[13][20][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][20][12] = (sum_out[14][20][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][20][12] = (sum_out[15][20][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][20][12] = (sum_out[16][20][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][20][12] = (sum_out[17][20][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][20][12] = (sum_out[18][20][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][20][12] = (sum_out[19][20][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][20][13] = (sum_out[0][20][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][20][13] = (sum_out[1][20][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][20][13] = (sum_out[2][20][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][20][13] = (sum_out[3][20][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][20][13] = (sum_out[4][20][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][20][13] = (sum_out[5][20][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][20][13] = (sum_out[6][20][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][20][13] = (sum_out[7][20][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][20][13] = (sum_out[8][20][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][20][13] = (sum_out[9][20][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][20][13] = (sum_out[10][20][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][20][13] = (sum_out[11][20][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][20][13] = (sum_out[12][20][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][20][13] = (sum_out[13][20][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][20][13] = (sum_out[14][20][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][20][13] = (sum_out[15][20][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][20][13] = (sum_out[16][20][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][20][13] = (sum_out[17][20][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][20][13] = (sum_out[18][20][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][20][13] = (sum_out[19][20][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][20][14] = (sum_out[0][20][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][20][14] = (sum_out[1][20][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][20][14] = (sum_out[2][20][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][20][14] = (sum_out[3][20][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][20][14] = (sum_out[4][20][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][20][14] = (sum_out[5][20][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][20][14] = (sum_out[6][20][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][20][14] = (sum_out[7][20][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][20][14] = (sum_out[8][20][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][20][14] = (sum_out[9][20][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][20][14] = (sum_out[10][20][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][20][14] = (sum_out[11][20][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][20][14] = (sum_out[12][20][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][20][14] = (sum_out[13][20][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][20][14] = (sum_out[14][20][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][20][14] = (sum_out[15][20][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][20][14] = (sum_out[16][20][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][20][14] = (sum_out[17][20][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][20][14] = (sum_out[18][20][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][20][14] = (sum_out[19][20][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][20][15] = (sum_out[0][20][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][20][15] = (sum_out[1][20][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][20][15] = (sum_out[2][20][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][20][15] = (sum_out[3][20][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][20][15] = (sum_out[4][20][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][20][15] = (sum_out[5][20][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][20][15] = (sum_out[6][20][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][20][15] = (sum_out[7][20][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][20][15] = (sum_out[8][20][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][20][15] = (sum_out[9][20][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][20][15] = (sum_out[10][20][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][20][15] = (sum_out[11][20][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][20][15] = (sum_out[12][20][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][20][15] = (sum_out[13][20][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][20][15] = (sum_out[14][20][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][20][15] = (sum_out[15][20][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][20][15] = (sum_out[16][20][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][20][15] = (sum_out[17][20][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][20][15] = (sum_out[18][20][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][20][15] = (sum_out[19][20][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][20][16] = (sum_out[0][20][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][20][16] = (sum_out[1][20][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][20][16] = (sum_out[2][20][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][20][16] = (sum_out[3][20][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][20][16] = (sum_out[4][20][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][20][16] = (sum_out[5][20][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][20][16] = (sum_out[6][20][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][20][16] = (sum_out[7][20][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][20][16] = (sum_out[8][20][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][20][16] = (sum_out[9][20][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][20][16] = (sum_out[10][20][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][20][16] = (sum_out[11][20][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][20][16] = (sum_out[12][20][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][20][16] = (sum_out[13][20][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][20][16] = (sum_out[14][20][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][20][16] = (sum_out[15][20][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][20][16] = (sum_out[16][20][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][20][16] = (sum_out[17][20][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][20][16] = (sum_out[18][20][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][20][16] = (sum_out[19][20][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][20][17] = (sum_out[0][20][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][20][17] = (sum_out[1][20][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][20][17] = (sum_out[2][20][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][20][17] = (sum_out[3][20][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][20][17] = (sum_out[4][20][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][20][17] = (sum_out[5][20][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][20][17] = (sum_out[6][20][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][20][17] = (sum_out[7][20][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][20][17] = (sum_out[8][20][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][20][17] = (sum_out[9][20][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][20][17] = (sum_out[10][20][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][20][17] = (sum_out[11][20][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][20][17] = (sum_out[12][20][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][20][17] = (sum_out[13][20][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][20][17] = (sum_out[14][20][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][20][17] = (sum_out[15][20][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][20][17] = (sum_out[16][20][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][20][17] = (sum_out[17][20][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][20][17] = (sum_out[18][20][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][20][17] = (sum_out[19][20][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][20][18] = (sum_out[0][20][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][20][18] = (sum_out[1][20][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][20][18] = (sum_out[2][20][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][20][18] = (sum_out[3][20][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][20][18] = (sum_out[4][20][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][20][18] = (sum_out[5][20][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][20][18] = (sum_out[6][20][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][20][18] = (sum_out[7][20][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][20][18] = (sum_out[8][20][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][20][18] = (sum_out[9][20][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][20][18] = (sum_out[10][20][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][20][18] = (sum_out[11][20][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][20][18] = (sum_out[12][20][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][20][18] = (sum_out[13][20][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][20][18] = (sum_out[14][20][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][20][18] = (sum_out[15][20][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][20][18] = (sum_out[16][20][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][20][18] = (sum_out[17][20][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][20][18] = (sum_out[18][20][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][20][18] = (sum_out[19][20][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][20][19] = (sum_out[0][20][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][20][19] = (sum_out[1][20][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][20][19] = (sum_out[2][20][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][20][19] = (sum_out[3][20][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][20][19] = (sum_out[4][20][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][20][19] = (sum_out[5][20][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][20][19] = (sum_out[6][20][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][20][19] = (sum_out[7][20][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][20][19] = (sum_out[8][20][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][20][19] = (sum_out[9][20][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][20][19] = (sum_out[10][20][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][20][19] = (sum_out[11][20][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][20][19] = (sum_out[12][20][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][20][19] = (sum_out[13][20][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][20][19] = (sum_out[14][20][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][20][19] = (sum_out[15][20][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][20][19] = (sum_out[16][20][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][20][19] = (sum_out[17][20][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][20][19] = (sum_out[18][20][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][20][19] = (sum_out[19][20][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][20][20] = (sum_out[0][20][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][20][20] = (sum_out[1][20][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][20][20] = (sum_out[2][20][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][20][20] = (sum_out[3][20][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][20][20] = (sum_out[4][20][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][20][20] = (sum_out[5][20][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][20][20] = (sum_out[6][20][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][20][20] = (sum_out[7][20][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][20][20] = (sum_out[8][20][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][20][20] = (sum_out[9][20][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][20][20] = (sum_out[10][20][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][20][20] = (sum_out[11][20][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][20][20] = (sum_out[12][20][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][20][20] = (sum_out[13][20][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][20][20] = (sum_out[14][20][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][20][20] = (sum_out[15][20][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][20][20] = (sum_out[16][20][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][20][20] = (sum_out[17][20][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][20][20] = (sum_out[18][20][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][20][20] = (sum_out[19][20][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][20][21] = (sum_out[0][20][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][20][21] = (sum_out[1][20][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][20][21] = (sum_out[2][20][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][20][21] = (sum_out[3][20][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][20][21] = (sum_out[4][20][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][20][21] = (sum_out[5][20][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][20][21] = (sum_out[6][20][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][20][21] = (sum_out[7][20][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][20][21] = (sum_out[8][20][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][20][21] = (sum_out[9][20][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][20][21] = (sum_out[10][20][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][20][21] = (sum_out[11][20][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][20][21] = (sum_out[12][20][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][20][21] = (sum_out[13][20][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][20][21] = (sum_out[14][20][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][20][21] = (sum_out[15][20][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][20][21] = (sum_out[16][20][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][20][21] = (sum_out[17][20][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][20][21] = (sum_out[18][20][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][20][21] = (sum_out[19][20][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][20][22] = (sum_out[0][20][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][20][22] = (sum_out[1][20][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][20][22] = (sum_out[2][20][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][20][22] = (sum_out[3][20][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][20][22] = (sum_out[4][20][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][20][22] = (sum_out[5][20][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][20][22] = (sum_out[6][20][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][20][22] = (sum_out[7][20][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][20][22] = (sum_out[8][20][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][20][22] = (sum_out[9][20][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][20][22] = (sum_out[10][20][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][20][22] = (sum_out[11][20][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][20][22] = (sum_out[12][20][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][20][22] = (sum_out[13][20][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][20][22] = (sum_out[14][20][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][20][22] = (sum_out[15][20][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][20][22] = (sum_out[16][20][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][20][22] = (sum_out[17][20][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][20][22] = (sum_out[18][20][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][20][22] = (sum_out[19][20][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][20][23] = (sum_out[0][20][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][20][23] = (sum_out[1][20][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][20][23] = (sum_out[2][20][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][20][23] = (sum_out[3][20][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][20][23] = (sum_out[4][20][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][20][23] = (sum_out[5][20][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][20][23] = (sum_out[6][20][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][20][23] = (sum_out[7][20][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][20][23] = (sum_out[8][20][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][20][23] = (sum_out[9][20][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][20][23] = (sum_out[10][20][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][20][23] = (sum_out[11][20][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][20][23] = (sum_out[12][20][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][20][23] = (sum_out[13][20][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][20][23] = (sum_out[14][20][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][20][23] = (sum_out[15][20][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][20][23] = (sum_out[16][20][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][20][23] = (sum_out[17][20][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][20][23] = (sum_out[18][20][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][20][23] = (sum_out[19][20][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][21][0] = (sum_out[0][21][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][21][0] = (sum_out[1][21][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][21][0] = (sum_out[2][21][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][21][0] = (sum_out[3][21][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][21][0] = (sum_out[4][21][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][21][0] = (sum_out[5][21][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][21][0] = (sum_out[6][21][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][21][0] = (sum_out[7][21][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][21][0] = (sum_out[8][21][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][21][0] = (sum_out[9][21][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][21][0] = (sum_out[10][21][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][21][0] = (sum_out[11][21][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][21][0] = (sum_out[12][21][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][21][0] = (sum_out[13][21][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][21][0] = (sum_out[14][21][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][21][0] = (sum_out[15][21][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][21][0] = (sum_out[16][21][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][21][0] = (sum_out[17][21][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][21][0] = (sum_out[18][21][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][21][0] = (sum_out[19][21][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][21][1] = (sum_out[0][21][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][21][1] = (sum_out[1][21][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][21][1] = (sum_out[2][21][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][21][1] = (sum_out[3][21][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][21][1] = (sum_out[4][21][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][21][1] = (sum_out[5][21][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][21][1] = (sum_out[6][21][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][21][1] = (sum_out[7][21][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][21][1] = (sum_out[8][21][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][21][1] = (sum_out[9][21][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][21][1] = (sum_out[10][21][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][21][1] = (sum_out[11][21][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][21][1] = (sum_out[12][21][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][21][1] = (sum_out[13][21][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][21][1] = (sum_out[14][21][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][21][1] = (sum_out[15][21][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][21][1] = (sum_out[16][21][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][21][1] = (sum_out[17][21][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][21][1] = (sum_out[18][21][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][21][1] = (sum_out[19][21][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][21][2] = (sum_out[0][21][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][21][2] = (sum_out[1][21][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][21][2] = (sum_out[2][21][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][21][2] = (sum_out[3][21][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][21][2] = (sum_out[4][21][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][21][2] = (sum_out[5][21][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][21][2] = (sum_out[6][21][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][21][2] = (sum_out[7][21][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][21][2] = (sum_out[8][21][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][21][2] = (sum_out[9][21][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][21][2] = (sum_out[10][21][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][21][2] = (sum_out[11][21][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][21][2] = (sum_out[12][21][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][21][2] = (sum_out[13][21][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][21][2] = (sum_out[14][21][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][21][2] = (sum_out[15][21][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][21][2] = (sum_out[16][21][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][21][2] = (sum_out[17][21][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][21][2] = (sum_out[18][21][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][21][2] = (sum_out[19][21][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][21][3] = (sum_out[0][21][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][21][3] = (sum_out[1][21][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][21][3] = (sum_out[2][21][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][21][3] = (sum_out[3][21][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][21][3] = (sum_out[4][21][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][21][3] = (sum_out[5][21][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][21][3] = (sum_out[6][21][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][21][3] = (sum_out[7][21][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][21][3] = (sum_out[8][21][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][21][3] = (sum_out[9][21][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][21][3] = (sum_out[10][21][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][21][3] = (sum_out[11][21][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][21][3] = (sum_out[12][21][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][21][3] = (sum_out[13][21][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][21][3] = (sum_out[14][21][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][21][3] = (sum_out[15][21][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][21][3] = (sum_out[16][21][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][21][3] = (sum_out[17][21][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][21][3] = (sum_out[18][21][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][21][3] = (sum_out[19][21][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][21][4] = (sum_out[0][21][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][21][4] = (sum_out[1][21][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][21][4] = (sum_out[2][21][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][21][4] = (sum_out[3][21][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][21][4] = (sum_out[4][21][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][21][4] = (sum_out[5][21][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][21][4] = (sum_out[6][21][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][21][4] = (sum_out[7][21][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][21][4] = (sum_out[8][21][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][21][4] = (sum_out[9][21][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][21][4] = (sum_out[10][21][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][21][4] = (sum_out[11][21][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][21][4] = (sum_out[12][21][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][21][4] = (sum_out[13][21][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][21][4] = (sum_out[14][21][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][21][4] = (sum_out[15][21][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][21][4] = (sum_out[16][21][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][21][4] = (sum_out[17][21][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][21][4] = (sum_out[18][21][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][21][4] = (sum_out[19][21][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][21][5] = (sum_out[0][21][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][21][5] = (sum_out[1][21][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][21][5] = (sum_out[2][21][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][21][5] = (sum_out[3][21][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][21][5] = (sum_out[4][21][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][21][5] = (sum_out[5][21][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][21][5] = (sum_out[6][21][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][21][5] = (sum_out[7][21][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][21][5] = (sum_out[8][21][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][21][5] = (sum_out[9][21][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][21][5] = (sum_out[10][21][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][21][5] = (sum_out[11][21][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][21][5] = (sum_out[12][21][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][21][5] = (sum_out[13][21][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][21][5] = (sum_out[14][21][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][21][5] = (sum_out[15][21][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][21][5] = (sum_out[16][21][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][21][5] = (sum_out[17][21][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][21][5] = (sum_out[18][21][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][21][5] = (sum_out[19][21][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][21][6] = (sum_out[0][21][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][21][6] = (sum_out[1][21][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][21][6] = (sum_out[2][21][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][21][6] = (sum_out[3][21][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][21][6] = (sum_out[4][21][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][21][6] = (sum_out[5][21][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][21][6] = (sum_out[6][21][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][21][6] = (sum_out[7][21][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][21][6] = (sum_out[8][21][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][21][6] = (sum_out[9][21][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][21][6] = (sum_out[10][21][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][21][6] = (sum_out[11][21][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][21][6] = (sum_out[12][21][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][21][6] = (sum_out[13][21][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][21][6] = (sum_out[14][21][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][21][6] = (sum_out[15][21][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][21][6] = (sum_out[16][21][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][21][6] = (sum_out[17][21][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][21][6] = (sum_out[18][21][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][21][6] = (sum_out[19][21][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][21][7] = (sum_out[0][21][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][21][7] = (sum_out[1][21][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][21][7] = (sum_out[2][21][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][21][7] = (sum_out[3][21][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][21][7] = (sum_out[4][21][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][21][7] = (sum_out[5][21][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][21][7] = (sum_out[6][21][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][21][7] = (sum_out[7][21][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][21][7] = (sum_out[8][21][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][21][7] = (sum_out[9][21][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][21][7] = (sum_out[10][21][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][21][7] = (sum_out[11][21][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][21][7] = (sum_out[12][21][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][21][7] = (sum_out[13][21][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][21][7] = (sum_out[14][21][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][21][7] = (sum_out[15][21][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][21][7] = (sum_out[16][21][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][21][7] = (sum_out[17][21][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][21][7] = (sum_out[18][21][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][21][7] = (sum_out[19][21][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][21][8] = (sum_out[0][21][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][21][8] = (sum_out[1][21][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][21][8] = (sum_out[2][21][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][21][8] = (sum_out[3][21][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][21][8] = (sum_out[4][21][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][21][8] = (sum_out[5][21][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][21][8] = (sum_out[6][21][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][21][8] = (sum_out[7][21][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][21][8] = (sum_out[8][21][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][21][8] = (sum_out[9][21][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][21][8] = (sum_out[10][21][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][21][8] = (sum_out[11][21][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][21][8] = (sum_out[12][21][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][21][8] = (sum_out[13][21][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][21][8] = (sum_out[14][21][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][21][8] = (sum_out[15][21][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][21][8] = (sum_out[16][21][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][21][8] = (sum_out[17][21][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][21][8] = (sum_out[18][21][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][21][8] = (sum_out[19][21][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][21][9] = (sum_out[0][21][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][21][9] = (sum_out[1][21][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][21][9] = (sum_out[2][21][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][21][9] = (sum_out[3][21][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][21][9] = (sum_out[4][21][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][21][9] = (sum_out[5][21][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][21][9] = (sum_out[6][21][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][21][9] = (sum_out[7][21][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][21][9] = (sum_out[8][21][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][21][9] = (sum_out[9][21][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][21][9] = (sum_out[10][21][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][21][9] = (sum_out[11][21][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][21][9] = (sum_out[12][21][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][21][9] = (sum_out[13][21][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][21][9] = (sum_out[14][21][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][21][9] = (sum_out[15][21][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][21][9] = (sum_out[16][21][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][21][9] = (sum_out[17][21][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][21][9] = (sum_out[18][21][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][21][9] = (sum_out[19][21][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][21][10] = (sum_out[0][21][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][21][10] = (sum_out[1][21][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][21][10] = (sum_out[2][21][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][21][10] = (sum_out[3][21][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][21][10] = (sum_out[4][21][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][21][10] = (sum_out[5][21][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][21][10] = (sum_out[6][21][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][21][10] = (sum_out[7][21][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][21][10] = (sum_out[8][21][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][21][10] = (sum_out[9][21][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][21][10] = (sum_out[10][21][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][21][10] = (sum_out[11][21][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][21][10] = (sum_out[12][21][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][21][10] = (sum_out[13][21][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][21][10] = (sum_out[14][21][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][21][10] = (sum_out[15][21][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][21][10] = (sum_out[16][21][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][21][10] = (sum_out[17][21][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][21][10] = (sum_out[18][21][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][21][10] = (sum_out[19][21][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][21][11] = (sum_out[0][21][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][21][11] = (sum_out[1][21][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][21][11] = (sum_out[2][21][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][21][11] = (sum_out[3][21][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][21][11] = (sum_out[4][21][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][21][11] = (sum_out[5][21][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][21][11] = (sum_out[6][21][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][21][11] = (sum_out[7][21][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][21][11] = (sum_out[8][21][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][21][11] = (sum_out[9][21][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][21][11] = (sum_out[10][21][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][21][11] = (sum_out[11][21][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][21][11] = (sum_out[12][21][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][21][11] = (sum_out[13][21][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][21][11] = (sum_out[14][21][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][21][11] = (sum_out[15][21][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][21][11] = (sum_out[16][21][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][21][11] = (sum_out[17][21][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][21][11] = (sum_out[18][21][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][21][11] = (sum_out[19][21][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][21][12] = (sum_out[0][21][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][21][12] = (sum_out[1][21][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][21][12] = (sum_out[2][21][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][21][12] = (sum_out[3][21][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][21][12] = (sum_out[4][21][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][21][12] = (sum_out[5][21][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][21][12] = (sum_out[6][21][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][21][12] = (sum_out[7][21][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][21][12] = (sum_out[8][21][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][21][12] = (sum_out[9][21][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][21][12] = (sum_out[10][21][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][21][12] = (sum_out[11][21][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][21][12] = (sum_out[12][21][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][21][12] = (sum_out[13][21][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][21][12] = (sum_out[14][21][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][21][12] = (sum_out[15][21][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][21][12] = (sum_out[16][21][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][21][12] = (sum_out[17][21][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][21][12] = (sum_out[18][21][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][21][12] = (sum_out[19][21][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][21][13] = (sum_out[0][21][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][21][13] = (sum_out[1][21][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][21][13] = (sum_out[2][21][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][21][13] = (sum_out[3][21][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][21][13] = (sum_out[4][21][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][21][13] = (sum_out[5][21][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][21][13] = (sum_out[6][21][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][21][13] = (sum_out[7][21][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][21][13] = (sum_out[8][21][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][21][13] = (sum_out[9][21][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][21][13] = (sum_out[10][21][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][21][13] = (sum_out[11][21][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][21][13] = (sum_out[12][21][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][21][13] = (sum_out[13][21][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][21][13] = (sum_out[14][21][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][21][13] = (sum_out[15][21][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][21][13] = (sum_out[16][21][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][21][13] = (sum_out[17][21][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][21][13] = (sum_out[18][21][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][21][13] = (sum_out[19][21][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][21][14] = (sum_out[0][21][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][21][14] = (sum_out[1][21][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][21][14] = (sum_out[2][21][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][21][14] = (sum_out[3][21][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][21][14] = (sum_out[4][21][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][21][14] = (sum_out[5][21][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][21][14] = (sum_out[6][21][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][21][14] = (sum_out[7][21][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][21][14] = (sum_out[8][21][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][21][14] = (sum_out[9][21][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][21][14] = (sum_out[10][21][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][21][14] = (sum_out[11][21][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][21][14] = (sum_out[12][21][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][21][14] = (sum_out[13][21][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][21][14] = (sum_out[14][21][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][21][14] = (sum_out[15][21][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][21][14] = (sum_out[16][21][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][21][14] = (sum_out[17][21][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][21][14] = (sum_out[18][21][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][21][14] = (sum_out[19][21][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][21][15] = (sum_out[0][21][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][21][15] = (sum_out[1][21][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][21][15] = (sum_out[2][21][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][21][15] = (sum_out[3][21][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][21][15] = (sum_out[4][21][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][21][15] = (sum_out[5][21][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][21][15] = (sum_out[6][21][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][21][15] = (sum_out[7][21][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][21][15] = (sum_out[8][21][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][21][15] = (sum_out[9][21][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][21][15] = (sum_out[10][21][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][21][15] = (sum_out[11][21][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][21][15] = (sum_out[12][21][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][21][15] = (sum_out[13][21][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][21][15] = (sum_out[14][21][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][21][15] = (sum_out[15][21][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][21][15] = (sum_out[16][21][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][21][15] = (sum_out[17][21][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][21][15] = (sum_out[18][21][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][21][15] = (sum_out[19][21][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][21][16] = (sum_out[0][21][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][21][16] = (sum_out[1][21][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][21][16] = (sum_out[2][21][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][21][16] = (sum_out[3][21][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][21][16] = (sum_out[4][21][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][21][16] = (sum_out[5][21][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][21][16] = (sum_out[6][21][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][21][16] = (sum_out[7][21][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][21][16] = (sum_out[8][21][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][21][16] = (sum_out[9][21][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][21][16] = (sum_out[10][21][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][21][16] = (sum_out[11][21][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][21][16] = (sum_out[12][21][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][21][16] = (sum_out[13][21][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][21][16] = (sum_out[14][21][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][21][16] = (sum_out[15][21][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][21][16] = (sum_out[16][21][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][21][16] = (sum_out[17][21][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][21][16] = (sum_out[18][21][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][21][16] = (sum_out[19][21][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][21][17] = (sum_out[0][21][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][21][17] = (sum_out[1][21][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][21][17] = (sum_out[2][21][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][21][17] = (sum_out[3][21][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][21][17] = (sum_out[4][21][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][21][17] = (sum_out[5][21][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][21][17] = (sum_out[6][21][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][21][17] = (sum_out[7][21][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][21][17] = (sum_out[8][21][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][21][17] = (sum_out[9][21][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][21][17] = (sum_out[10][21][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][21][17] = (sum_out[11][21][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][21][17] = (sum_out[12][21][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][21][17] = (sum_out[13][21][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][21][17] = (sum_out[14][21][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][21][17] = (sum_out[15][21][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][21][17] = (sum_out[16][21][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][21][17] = (sum_out[17][21][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][21][17] = (sum_out[18][21][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][21][17] = (sum_out[19][21][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][21][18] = (sum_out[0][21][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][21][18] = (sum_out[1][21][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][21][18] = (sum_out[2][21][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][21][18] = (sum_out[3][21][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][21][18] = (sum_out[4][21][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][21][18] = (sum_out[5][21][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][21][18] = (sum_out[6][21][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][21][18] = (sum_out[7][21][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][21][18] = (sum_out[8][21][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][21][18] = (sum_out[9][21][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][21][18] = (sum_out[10][21][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][21][18] = (sum_out[11][21][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][21][18] = (sum_out[12][21][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][21][18] = (sum_out[13][21][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][21][18] = (sum_out[14][21][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][21][18] = (sum_out[15][21][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][21][18] = (sum_out[16][21][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][21][18] = (sum_out[17][21][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][21][18] = (sum_out[18][21][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][21][18] = (sum_out[19][21][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][21][19] = (sum_out[0][21][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][21][19] = (sum_out[1][21][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][21][19] = (sum_out[2][21][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][21][19] = (sum_out[3][21][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][21][19] = (sum_out[4][21][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][21][19] = (sum_out[5][21][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][21][19] = (sum_out[6][21][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][21][19] = (sum_out[7][21][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][21][19] = (sum_out[8][21][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][21][19] = (sum_out[9][21][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][21][19] = (sum_out[10][21][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][21][19] = (sum_out[11][21][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][21][19] = (sum_out[12][21][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][21][19] = (sum_out[13][21][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][21][19] = (sum_out[14][21][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][21][19] = (sum_out[15][21][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][21][19] = (sum_out[16][21][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][21][19] = (sum_out[17][21][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][21][19] = (sum_out[18][21][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][21][19] = (sum_out[19][21][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][21][20] = (sum_out[0][21][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][21][20] = (sum_out[1][21][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][21][20] = (sum_out[2][21][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][21][20] = (sum_out[3][21][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][21][20] = (sum_out[4][21][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][21][20] = (sum_out[5][21][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][21][20] = (sum_out[6][21][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][21][20] = (sum_out[7][21][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][21][20] = (sum_out[8][21][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][21][20] = (sum_out[9][21][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][21][20] = (sum_out[10][21][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][21][20] = (sum_out[11][21][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][21][20] = (sum_out[12][21][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][21][20] = (sum_out[13][21][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][21][20] = (sum_out[14][21][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][21][20] = (sum_out[15][21][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][21][20] = (sum_out[16][21][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][21][20] = (sum_out[17][21][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][21][20] = (sum_out[18][21][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][21][20] = (sum_out[19][21][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][21][21] = (sum_out[0][21][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][21][21] = (sum_out[1][21][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][21][21] = (sum_out[2][21][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][21][21] = (sum_out[3][21][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][21][21] = (sum_out[4][21][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][21][21] = (sum_out[5][21][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][21][21] = (sum_out[6][21][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][21][21] = (sum_out[7][21][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][21][21] = (sum_out[8][21][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][21][21] = (sum_out[9][21][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][21][21] = (sum_out[10][21][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][21][21] = (sum_out[11][21][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][21][21] = (sum_out[12][21][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][21][21] = (sum_out[13][21][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][21][21] = (sum_out[14][21][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][21][21] = (sum_out[15][21][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][21][21] = (sum_out[16][21][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][21][21] = (sum_out[17][21][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][21][21] = (sum_out[18][21][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][21][21] = (sum_out[19][21][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][21][22] = (sum_out[0][21][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][21][22] = (sum_out[1][21][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][21][22] = (sum_out[2][21][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][21][22] = (sum_out[3][21][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][21][22] = (sum_out[4][21][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][21][22] = (sum_out[5][21][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][21][22] = (sum_out[6][21][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][21][22] = (sum_out[7][21][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][21][22] = (sum_out[8][21][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][21][22] = (sum_out[9][21][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][21][22] = (sum_out[10][21][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][21][22] = (sum_out[11][21][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][21][22] = (sum_out[12][21][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][21][22] = (sum_out[13][21][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][21][22] = (sum_out[14][21][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][21][22] = (sum_out[15][21][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][21][22] = (sum_out[16][21][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][21][22] = (sum_out[17][21][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][21][22] = (sum_out[18][21][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][21][22] = (sum_out[19][21][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][21][23] = (sum_out[0][21][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][21][23] = (sum_out[1][21][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][21][23] = (sum_out[2][21][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][21][23] = (sum_out[3][21][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][21][23] = (sum_out[4][21][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][21][23] = (sum_out[5][21][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][21][23] = (sum_out[6][21][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][21][23] = (sum_out[7][21][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][21][23] = (sum_out[8][21][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][21][23] = (sum_out[9][21][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][21][23] = (sum_out[10][21][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][21][23] = (sum_out[11][21][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][21][23] = (sum_out[12][21][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][21][23] = (sum_out[13][21][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][21][23] = (sum_out[14][21][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][21][23] = (sum_out[15][21][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][21][23] = (sum_out[16][21][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][21][23] = (sum_out[17][21][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][21][23] = (sum_out[18][21][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][21][23] = (sum_out[19][21][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][22][0] = (sum_out[0][22][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][22][0] = (sum_out[1][22][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][22][0] = (sum_out[2][22][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][22][0] = (sum_out[3][22][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][22][0] = (sum_out[4][22][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][22][0] = (sum_out[5][22][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][22][0] = (sum_out[6][22][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][22][0] = (sum_out[7][22][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][22][0] = (sum_out[8][22][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][22][0] = (sum_out[9][22][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][22][0] = (sum_out[10][22][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][22][0] = (sum_out[11][22][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][22][0] = (sum_out[12][22][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][22][0] = (sum_out[13][22][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][22][0] = (sum_out[14][22][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][22][0] = (sum_out[15][22][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][22][0] = (sum_out[16][22][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][22][0] = (sum_out[17][22][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][22][0] = (sum_out[18][22][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][22][0] = (sum_out[19][22][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][22][1] = (sum_out[0][22][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][22][1] = (sum_out[1][22][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][22][1] = (sum_out[2][22][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][22][1] = (sum_out[3][22][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][22][1] = (sum_out[4][22][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][22][1] = (sum_out[5][22][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][22][1] = (sum_out[6][22][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][22][1] = (sum_out[7][22][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][22][1] = (sum_out[8][22][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][22][1] = (sum_out[9][22][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][22][1] = (sum_out[10][22][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][22][1] = (sum_out[11][22][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][22][1] = (sum_out[12][22][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][22][1] = (sum_out[13][22][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][22][1] = (sum_out[14][22][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][22][1] = (sum_out[15][22][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][22][1] = (sum_out[16][22][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][22][1] = (sum_out[17][22][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][22][1] = (sum_out[18][22][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][22][1] = (sum_out[19][22][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][22][2] = (sum_out[0][22][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][22][2] = (sum_out[1][22][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][22][2] = (sum_out[2][22][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][22][2] = (sum_out[3][22][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][22][2] = (sum_out[4][22][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][22][2] = (sum_out[5][22][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][22][2] = (sum_out[6][22][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][22][2] = (sum_out[7][22][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][22][2] = (sum_out[8][22][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][22][2] = (sum_out[9][22][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][22][2] = (sum_out[10][22][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][22][2] = (sum_out[11][22][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][22][2] = (sum_out[12][22][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][22][2] = (sum_out[13][22][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][22][2] = (sum_out[14][22][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][22][2] = (sum_out[15][22][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][22][2] = (sum_out[16][22][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][22][2] = (sum_out[17][22][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][22][2] = (sum_out[18][22][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][22][2] = (sum_out[19][22][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][22][3] = (sum_out[0][22][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][22][3] = (sum_out[1][22][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][22][3] = (sum_out[2][22][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][22][3] = (sum_out[3][22][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][22][3] = (sum_out[4][22][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][22][3] = (sum_out[5][22][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][22][3] = (sum_out[6][22][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][22][3] = (sum_out[7][22][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][22][3] = (sum_out[8][22][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][22][3] = (sum_out[9][22][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][22][3] = (sum_out[10][22][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][22][3] = (sum_out[11][22][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][22][3] = (sum_out[12][22][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][22][3] = (sum_out[13][22][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][22][3] = (sum_out[14][22][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][22][3] = (sum_out[15][22][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][22][3] = (sum_out[16][22][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][22][3] = (sum_out[17][22][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][22][3] = (sum_out[18][22][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][22][3] = (sum_out[19][22][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][22][4] = (sum_out[0][22][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][22][4] = (sum_out[1][22][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][22][4] = (sum_out[2][22][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][22][4] = (sum_out[3][22][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][22][4] = (sum_out[4][22][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][22][4] = (sum_out[5][22][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][22][4] = (sum_out[6][22][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][22][4] = (sum_out[7][22][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][22][4] = (sum_out[8][22][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][22][4] = (sum_out[9][22][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][22][4] = (sum_out[10][22][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][22][4] = (sum_out[11][22][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][22][4] = (sum_out[12][22][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][22][4] = (sum_out[13][22][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][22][4] = (sum_out[14][22][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][22][4] = (sum_out[15][22][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][22][4] = (sum_out[16][22][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][22][4] = (sum_out[17][22][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][22][4] = (sum_out[18][22][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][22][4] = (sum_out[19][22][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][22][5] = (sum_out[0][22][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][22][5] = (sum_out[1][22][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][22][5] = (sum_out[2][22][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][22][5] = (sum_out[3][22][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][22][5] = (sum_out[4][22][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][22][5] = (sum_out[5][22][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][22][5] = (sum_out[6][22][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][22][5] = (sum_out[7][22][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][22][5] = (sum_out[8][22][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][22][5] = (sum_out[9][22][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][22][5] = (sum_out[10][22][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][22][5] = (sum_out[11][22][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][22][5] = (sum_out[12][22][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][22][5] = (sum_out[13][22][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][22][5] = (sum_out[14][22][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][22][5] = (sum_out[15][22][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][22][5] = (sum_out[16][22][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][22][5] = (sum_out[17][22][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][22][5] = (sum_out[18][22][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][22][5] = (sum_out[19][22][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][22][6] = (sum_out[0][22][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][22][6] = (sum_out[1][22][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][22][6] = (sum_out[2][22][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][22][6] = (sum_out[3][22][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][22][6] = (sum_out[4][22][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][22][6] = (sum_out[5][22][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][22][6] = (sum_out[6][22][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][22][6] = (sum_out[7][22][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][22][6] = (sum_out[8][22][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][22][6] = (sum_out[9][22][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][22][6] = (sum_out[10][22][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][22][6] = (sum_out[11][22][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][22][6] = (sum_out[12][22][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][22][6] = (sum_out[13][22][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][22][6] = (sum_out[14][22][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][22][6] = (sum_out[15][22][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][22][6] = (sum_out[16][22][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][22][6] = (sum_out[17][22][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][22][6] = (sum_out[18][22][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][22][6] = (sum_out[19][22][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][22][7] = (sum_out[0][22][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][22][7] = (sum_out[1][22][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][22][7] = (sum_out[2][22][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][22][7] = (sum_out[3][22][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][22][7] = (sum_out[4][22][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][22][7] = (sum_out[5][22][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][22][7] = (sum_out[6][22][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][22][7] = (sum_out[7][22][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][22][7] = (sum_out[8][22][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][22][7] = (sum_out[9][22][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][22][7] = (sum_out[10][22][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][22][7] = (sum_out[11][22][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][22][7] = (sum_out[12][22][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][22][7] = (sum_out[13][22][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][22][7] = (sum_out[14][22][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][22][7] = (sum_out[15][22][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][22][7] = (sum_out[16][22][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][22][7] = (sum_out[17][22][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][22][7] = (sum_out[18][22][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][22][7] = (sum_out[19][22][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][22][8] = (sum_out[0][22][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][22][8] = (sum_out[1][22][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][22][8] = (sum_out[2][22][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][22][8] = (sum_out[3][22][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][22][8] = (sum_out[4][22][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][22][8] = (sum_out[5][22][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][22][8] = (sum_out[6][22][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][22][8] = (sum_out[7][22][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][22][8] = (sum_out[8][22][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][22][8] = (sum_out[9][22][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][22][8] = (sum_out[10][22][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][22][8] = (sum_out[11][22][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][22][8] = (sum_out[12][22][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][22][8] = (sum_out[13][22][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][22][8] = (sum_out[14][22][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][22][8] = (sum_out[15][22][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][22][8] = (sum_out[16][22][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][22][8] = (sum_out[17][22][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][22][8] = (sum_out[18][22][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][22][8] = (sum_out[19][22][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][22][9] = (sum_out[0][22][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][22][9] = (sum_out[1][22][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][22][9] = (sum_out[2][22][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][22][9] = (sum_out[3][22][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][22][9] = (sum_out[4][22][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][22][9] = (sum_out[5][22][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][22][9] = (sum_out[6][22][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][22][9] = (sum_out[7][22][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][22][9] = (sum_out[8][22][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][22][9] = (sum_out[9][22][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][22][9] = (sum_out[10][22][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][22][9] = (sum_out[11][22][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][22][9] = (sum_out[12][22][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][22][9] = (sum_out[13][22][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][22][9] = (sum_out[14][22][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][22][9] = (sum_out[15][22][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][22][9] = (sum_out[16][22][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][22][9] = (sum_out[17][22][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][22][9] = (sum_out[18][22][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][22][9] = (sum_out[19][22][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][22][10] = (sum_out[0][22][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][22][10] = (sum_out[1][22][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][22][10] = (sum_out[2][22][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][22][10] = (sum_out[3][22][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][22][10] = (sum_out[4][22][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][22][10] = (sum_out[5][22][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][22][10] = (sum_out[6][22][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][22][10] = (sum_out[7][22][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][22][10] = (sum_out[8][22][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][22][10] = (sum_out[9][22][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][22][10] = (sum_out[10][22][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][22][10] = (sum_out[11][22][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][22][10] = (sum_out[12][22][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][22][10] = (sum_out[13][22][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][22][10] = (sum_out[14][22][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][22][10] = (sum_out[15][22][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][22][10] = (sum_out[16][22][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][22][10] = (sum_out[17][22][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][22][10] = (sum_out[18][22][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][22][10] = (sum_out[19][22][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][22][11] = (sum_out[0][22][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][22][11] = (sum_out[1][22][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][22][11] = (sum_out[2][22][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][22][11] = (sum_out[3][22][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][22][11] = (sum_out[4][22][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][22][11] = (sum_out[5][22][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][22][11] = (sum_out[6][22][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][22][11] = (sum_out[7][22][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][22][11] = (sum_out[8][22][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][22][11] = (sum_out[9][22][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][22][11] = (sum_out[10][22][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][22][11] = (sum_out[11][22][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][22][11] = (sum_out[12][22][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][22][11] = (sum_out[13][22][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][22][11] = (sum_out[14][22][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][22][11] = (sum_out[15][22][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][22][11] = (sum_out[16][22][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][22][11] = (sum_out[17][22][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][22][11] = (sum_out[18][22][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][22][11] = (sum_out[19][22][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][22][12] = (sum_out[0][22][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][22][12] = (sum_out[1][22][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][22][12] = (sum_out[2][22][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][22][12] = (sum_out[3][22][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][22][12] = (sum_out[4][22][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][22][12] = (sum_out[5][22][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][22][12] = (sum_out[6][22][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][22][12] = (sum_out[7][22][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][22][12] = (sum_out[8][22][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][22][12] = (sum_out[9][22][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][22][12] = (sum_out[10][22][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][22][12] = (sum_out[11][22][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][22][12] = (sum_out[12][22][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][22][12] = (sum_out[13][22][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][22][12] = (sum_out[14][22][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][22][12] = (sum_out[15][22][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][22][12] = (sum_out[16][22][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][22][12] = (sum_out[17][22][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][22][12] = (sum_out[18][22][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][22][12] = (sum_out[19][22][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][22][13] = (sum_out[0][22][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][22][13] = (sum_out[1][22][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][22][13] = (sum_out[2][22][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][22][13] = (sum_out[3][22][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][22][13] = (sum_out[4][22][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][22][13] = (sum_out[5][22][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][22][13] = (sum_out[6][22][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][22][13] = (sum_out[7][22][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][22][13] = (sum_out[8][22][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][22][13] = (sum_out[9][22][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][22][13] = (sum_out[10][22][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][22][13] = (sum_out[11][22][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][22][13] = (sum_out[12][22][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][22][13] = (sum_out[13][22][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][22][13] = (sum_out[14][22][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][22][13] = (sum_out[15][22][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][22][13] = (sum_out[16][22][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][22][13] = (sum_out[17][22][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][22][13] = (sum_out[18][22][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][22][13] = (sum_out[19][22][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][22][14] = (sum_out[0][22][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][22][14] = (sum_out[1][22][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][22][14] = (sum_out[2][22][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][22][14] = (sum_out[3][22][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][22][14] = (sum_out[4][22][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][22][14] = (sum_out[5][22][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][22][14] = (sum_out[6][22][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][22][14] = (sum_out[7][22][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][22][14] = (sum_out[8][22][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][22][14] = (sum_out[9][22][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][22][14] = (sum_out[10][22][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][22][14] = (sum_out[11][22][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][22][14] = (sum_out[12][22][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][22][14] = (sum_out[13][22][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][22][14] = (sum_out[14][22][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][22][14] = (sum_out[15][22][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][22][14] = (sum_out[16][22][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][22][14] = (sum_out[17][22][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][22][14] = (sum_out[18][22][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][22][14] = (sum_out[19][22][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][22][15] = (sum_out[0][22][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][22][15] = (sum_out[1][22][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][22][15] = (sum_out[2][22][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][22][15] = (sum_out[3][22][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][22][15] = (sum_out[4][22][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][22][15] = (sum_out[5][22][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][22][15] = (sum_out[6][22][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][22][15] = (sum_out[7][22][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][22][15] = (sum_out[8][22][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][22][15] = (sum_out[9][22][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][22][15] = (sum_out[10][22][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][22][15] = (sum_out[11][22][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][22][15] = (sum_out[12][22][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][22][15] = (sum_out[13][22][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][22][15] = (sum_out[14][22][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][22][15] = (sum_out[15][22][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][22][15] = (sum_out[16][22][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][22][15] = (sum_out[17][22][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][22][15] = (sum_out[18][22][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][22][15] = (sum_out[19][22][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][22][16] = (sum_out[0][22][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][22][16] = (sum_out[1][22][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][22][16] = (sum_out[2][22][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][22][16] = (sum_out[3][22][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][22][16] = (sum_out[4][22][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][22][16] = (sum_out[5][22][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][22][16] = (sum_out[6][22][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][22][16] = (sum_out[7][22][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][22][16] = (sum_out[8][22][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][22][16] = (sum_out[9][22][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][22][16] = (sum_out[10][22][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][22][16] = (sum_out[11][22][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][22][16] = (sum_out[12][22][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][22][16] = (sum_out[13][22][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][22][16] = (sum_out[14][22][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][22][16] = (sum_out[15][22][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][22][16] = (sum_out[16][22][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][22][16] = (sum_out[17][22][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][22][16] = (sum_out[18][22][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][22][16] = (sum_out[19][22][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][22][17] = (sum_out[0][22][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][22][17] = (sum_out[1][22][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][22][17] = (sum_out[2][22][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][22][17] = (sum_out[3][22][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][22][17] = (sum_out[4][22][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][22][17] = (sum_out[5][22][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][22][17] = (sum_out[6][22][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][22][17] = (sum_out[7][22][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][22][17] = (sum_out[8][22][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][22][17] = (sum_out[9][22][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][22][17] = (sum_out[10][22][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][22][17] = (sum_out[11][22][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][22][17] = (sum_out[12][22][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][22][17] = (sum_out[13][22][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][22][17] = (sum_out[14][22][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][22][17] = (sum_out[15][22][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][22][17] = (sum_out[16][22][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][22][17] = (sum_out[17][22][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][22][17] = (sum_out[18][22][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][22][17] = (sum_out[19][22][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][22][18] = (sum_out[0][22][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][22][18] = (sum_out[1][22][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][22][18] = (sum_out[2][22][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][22][18] = (sum_out[3][22][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][22][18] = (sum_out[4][22][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][22][18] = (sum_out[5][22][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][22][18] = (sum_out[6][22][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][22][18] = (sum_out[7][22][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][22][18] = (sum_out[8][22][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][22][18] = (sum_out[9][22][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][22][18] = (sum_out[10][22][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][22][18] = (sum_out[11][22][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][22][18] = (sum_out[12][22][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][22][18] = (sum_out[13][22][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][22][18] = (sum_out[14][22][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][22][18] = (sum_out[15][22][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][22][18] = (sum_out[16][22][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][22][18] = (sum_out[17][22][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][22][18] = (sum_out[18][22][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][22][18] = (sum_out[19][22][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][22][19] = (sum_out[0][22][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][22][19] = (sum_out[1][22][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][22][19] = (sum_out[2][22][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][22][19] = (sum_out[3][22][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][22][19] = (sum_out[4][22][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][22][19] = (sum_out[5][22][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][22][19] = (sum_out[6][22][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][22][19] = (sum_out[7][22][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][22][19] = (sum_out[8][22][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][22][19] = (sum_out[9][22][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][22][19] = (sum_out[10][22][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][22][19] = (sum_out[11][22][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][22][19] = (sum_out[12][22][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][22][19] = (sum_out[13][22][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][22][19] = (sum_out[14][22][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][22][19] = (sum_out[15][22][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][22][19] = (sum_out[16][22][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][22][19] = (sum_out[17][22][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][22][19] = (sum_out[18][22][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][22][19] = (sum_out[19][22][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][22][20] = (sum_out[0][22][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][22][20] = (sum_out[1][22][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][22][20] = (sum_out[2][22][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][22][20] = (sum_out[3][22][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][22][20] = (sum_out[4][22][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][22][20] = (sum_out[5][22][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][22][20] = (sum_out[6][22][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][22][20] = (sum_out[7][22][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][22][20] = (sum_out[8][22][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][22][20] = (sum_out[9][22][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][22][20] = (sum_out[10][22][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][22][20] = (sum_out[11][22][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][22][20] = (sum_out[12][22][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][22][20] = (sum_out[13][22][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][22][20] = (sum_out[14][22][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][22][20] = (sum_out[15][22][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][22][20] = (sum_out[16][22][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][22][20] = (sum_out[17][22][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][22][20] = (sum_out[18][22][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][22][20] = (sum_out[19][22][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][22][21] = (sum_out[0][22][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][22][21] = (sum_out[1][22][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][22][21] = (sum_out[2][22][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][22][21] = (sum_out[3][22][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][22][21] = (sum_out[4][22][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][22][21] = (sum_out[5][22][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][22][21] = (sum_out[6][22][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][22][21] = (sum_out[7][22][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][22][21] = (sum_out[8][22][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][22][21] = (sum_out[9][22][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][22][21] = (sum_out[10][22][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][22][21] = (sum_out[11][22][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][22][21] = (sum_out[12][22][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][22][21] = (sum_out[13][22][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][22][21] = (sum_out[14][22][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][22][21] = (sum_out[15][22][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][22][21] = (sum_out[16][22][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][22][21] = (sum_out[17][22][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][22][21] = (sum_out[18][22][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][22][21] = (sum_out[19][22][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][22][22] = (sum_out[0][22][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][22][22] = (sum_out[1][22][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][22][22] = (sum_out[2][22][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][22][22] = (sum_out[3][22][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][22][22] = (sum_out[4][22][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][22][22] = (sum_out[5][22][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][22][22] = (sum_out[6][22][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][22][22] = (sum_out[7][22][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][22][22] = (sum_out[8][22][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][22][22] = (sum_out[9][22][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][22][22] = (sum_out[10][22][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][22][22] = (sum_out[11][22][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][22][22] = (sum_out[12][22][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][22][22] = (sum_out[13][22][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][22][22] = (sum_out[14][22][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][22][22] = (sum_out[15][22][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][22][22] = (sum_out[16][22][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][22][22] = (sum_out[17][22][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][22][22] = (sum_out[18][22][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][22][22] = (sum_out[19][22][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][22][23] = (sum_out[0][22][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][22][23] = (sum_out[1][22][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][22][23] = (sum_out[2][22][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][22][23] = (sum_out[3][22][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][22][23] = (sum_out[4][22][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][22][23] = (sum_out[5][22][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][22][23] = (sum_out[6][22][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][22][23] = (sum_out[7][22][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][22][23] = (sum_out[8][22][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][22][23] = (sum_out[9][22][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][22][23] = (sum_out[10][22][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][22][23] = (sum_out[11][22][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][22][23] = (sum_out[12][22][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][22][23] = (sum_out[13][22][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][22][23] = (sum_out[14][22][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][22][23] = (sum_out[15][22][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][22][23] = (sum_out[16][22][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][22][23] = (sum_out[17][22][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][22][23] = (sum_out[18][22][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][22][23] = (sum_out[19][22][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][23][0] = (sum_out[0][23][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][23][0] = (sum_out[1][23][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][23][0] = (sum_out[2][23][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][23][0] = (sum_out[3][23][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][23][0] = (sum_out[4][23][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][23][0] = (sum_out[5][23][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][23][0] = (sum_out[6][23][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][23][0] = (sum_out[7][23][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][23][0] = (sum_out[8][23][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][23][0] = (sum_out[9][23][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][23][0] = (sum_out[10][23][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][23][0] = (sum_out[11][23][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][23][0] = (sum_out[12][23][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][23][0] = (sum_out[13][23][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][23][0] = (sum_out[14][23][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][23][0] = (sum_out[15][23][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][23][0] = (sum_out[16][23][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][23][0] = (sum_out[17][23][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][23][0] = (sum_out[18][23][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][23][0] = (sum_out[19][23][0] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][23][1] = (sum_out[0][23][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][23][1] = (sum_out[1][23][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][23][1] = (sum_out[2][23][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][23][1] = (sum_out[3][23][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][23][1] = (sum_out[4][23][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][23][1] = (sum_out[5][23][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][23][1] = (sum_out[6][23][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][23][1] = (sum_out[7][23][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][23][1] = (sum_out[8][23][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][23][1] = (sum_out[9][23][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][23][1] = (sum_out[10][23][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][23][1] = (sum_out[11][23][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][23][1] = (sum_out[12][23][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][23][1] = (sum_out[13][23][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][23][1] = (sum_out[14][23][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][23][1] = (sum_out[15][23][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][23][1] = (sum_out[16][23][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][23][1] = (sum_out[17][23][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][23][1] = (sum_out[18][23][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][23][1] = (sum_out[19][23][1] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][23][2] = (sum_out[0][23][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][23][2] = (sum_out[1][23][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][23][2] = (sum_out[2][23][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][23][2] = (sum_out[3][23][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][23][2] = (sum_out[4][23][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][23][2] = (sum_out[5][23][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][23][2] = (sum_out[6][23][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][23][2] = (sum_out[7][23][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][23][2] = (sum_out[8][23][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][23][2] = (sum_out[9][23][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][23][2] = (sum_out[10][23][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][23][2] = (sum_out[11][23][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][23][2] = (sum_out[12][23][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][23][2] = (sum_out[13][23][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][23][2] = (sum_out[14][23][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][23][2] = (sum_out[15][23][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][23][2] = (sum_out[16][23][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][23][2] = (sum_out[17][23][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][23][2] = (sum_out[18][23][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][23][2] = (sum_out[19][23][2] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][23][3] = (sum_out[0][23][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][23][3] = (sum_out[1][23][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][23][3] = (sum_out[2][23][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][23][3] = (sum_out[3][23][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][23][3] = (sum_out[4][23][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][23][3] = (sum_out[5][23][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][23][3] = (sum_out[6][23][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][23][3] = (sum_out[7][23][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][23][3] = (sum_out[8][23][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][23][3] = (sum_out[9][23][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][23][3] = (sum_out[10][23][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][23][3] = (sum_out[11][23][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][23][3] = (sum_out[12][23][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][23][3] = (sum_out[13][23][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][23][3] = (sum_out[14][23][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][23][3] = (sum_out[15][23][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][23][3] = (sum_out[16][23][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][23][3] = (sum_out[17][23][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][23][3] = (sum_out[18][23][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][23][3] = (sum_out[19][23][3] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][23][4] = (sum_out[0][23][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][23][4] = (sum_out[1][23][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][23][4] = (sum_out[2][23][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][23][4] = (sum_out[3][23][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][23][4] = (sum_out[4][23][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][23][4] = (sum_out[5][23][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][23][4] = (sum_out[6][23][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][23][4] = (sum_out[7][23][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][23][4] = (sum_out[8][23][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][23][4] = (sum_out[9][23][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][23][4] = (sum_out[10][23][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][23][4] = (sum_out[11][23][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][23][4] = (sum_out[12][23][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][23][4] = (sum_out[13][23][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][23][4] = (sum_out[14][23][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][23][4] = (sum_out[15][23][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][23][4] = (sum_out[16][23][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][23][4] = (sum_out[17][23][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][23][4] = (sum_out[18][23][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][23][4] = (sum_out[19][23][4] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][23][5] = (sum_out[0][23][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][23][5] = (sum_out[1][23][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][23][5] = (sum_out[2][23][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][23][5] = (sum_out[3][23][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][23][5] = (sum_out[4][23][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][23][5] = (sum_out[5][23][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][23][5] = (sum_out[6][23][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][23][5] = (sum_out[7][23][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][23][5] = (sum_out[8][23][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][23][5] = (sum_out[9][23][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][23][5] = (sum_out[10][23][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][23][5] = (sum_out[11][23][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][23][5] = (sum_out[12][23][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][23][5] = (sum_out[13][23][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][23][5] = (sum_out[14][23][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][23][5] = (sum_out[15][23][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][23][5] = (sum_out[16][23][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][23][5] = (sum_out[17][23][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][23][5] = (sum_out[18][23][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][23][5] = (sum_out[19][23][5] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][23][6] = (sum_out[0][23][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][23][6] = (sum_out[1][23][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][23][6] = (sum_out[2][23][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][23][6] = (sum_out[3][23][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][23][6] = (sum_out[4][23][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][23][6] = (sum_out[5][23][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][23][6] = (sum_out[6][23][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][23][6] = (sum_out[7][23][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][23][6] = (sum_out[8][23][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][23][6] = (sum_out[9][23][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][23][6] = (sum_out[10][23][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][23][6] = (sum_out[11][23][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][23][6] = (sum_out[12][23][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][23][6] = (sum_out[13][23][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][23][6] = (sum_out[14][23][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][23][6] = (sum_out[15][23][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][23][6] = (sum_out[16][23][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][23][6] = (sum_out[17][23][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][23][6] = (sum_out[18][23][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][23][6] = (sum_out[19][23][6] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][23][7] = (sum_out[0][23][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][23][7] = (sum_out[1][23][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][23][7] = (sum_out[2][23][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][23][7] = (sum_out[3][23][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][23][7] = (sum_out[4][23][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][23][7] = (sum_out[5][23][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][23][7] = (sum_out[6][23][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][23][7] = (sum_out[7][23][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][23][7] = (sum_out[8][23][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][23][7] = (sum_out[9][23][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][23][7] = (sum_out[10][23][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][23][7] = (sum_out[11][23][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][23][7] = (sum_out[12][23][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][23][7] = (sum_out[13][23][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][23][7] = (sum_out[14][23][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][23][7] = (sum_out[15][23][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][23][7] = (sum_out[16][23][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][23][7] = (sum_out[17][23][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][23][7] = (sum_out[18][23][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][23][7] = (sum_out[19][23][7] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][23][8] = (sum_out[0][23][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][23][8] = (sum_out[1][23][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][23][8] = (sum_out[2][23][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][23][8] = (sum_out[3][23][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][23][8] = (sum_out[4][23][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][23][8] = (sum_out[5][23][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][23][8] = (sum_out[6][23][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][23][8] = (sum_out[7][23][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][23][8] = (sum_out[8][23][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][23][8] = (sum_out[9][23][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][23][8] = (sum_out[10][23][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][23][8] = (sum_out[11][23][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][23][8] = (sum_out[12][23][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][23][8] = (sum_out[13][23][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][23][8] = (sum_out[14][23][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][23][8] = (sum_out[15][23][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][23][8] = (sum_out[16][23][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][23][8] = (sum_out[17][23][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][23][8] = (sum_out[18][23][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][23][8] = (sum_out[19][23][8] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][23][9] = (sum_out[0][23][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][23][9] = (sum_out[1][23][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][23][9] = (sum_out[2][23][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][23][9] = (sum_out[3][23][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][23][9] = (sum_out[4][23][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][23][9] = (sum_out[5][23][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][23][9] = (sum_out[6][23][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][23][9] = (sum_out[7][23][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][23][9] = (sum_out[8][23][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][23][9] = (sum_out[9][23][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][23][9] = (sum_out[10][23][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][23][9] = (sum_out[11][23][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][23][9] = (sum_out[12][23][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][23][9] = (sum_out[13][23][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][23][9] = (sum_out[14][23][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][23][9] = (sum_out[15][23][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][23][9] = (sum_out[16][23][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][23][9] = (sum_out[17][23][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][23][9] = (sum_out[18][23][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][23][9] = (sum_out[19][23][9] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][23][10] = (sum_out[0][23][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][23][10] = (sum_out[1][23][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][23][10] = (sum_out[2][23][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][23][10] = (sum_out[3][23][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][23][10] = (sum_out[4][23][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][23][10] = (sum_out[5][23][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][23][10] = (sum_out[6][23][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][23][10] = (sum_out[7][23][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][23][10] = (sum_out[8][23][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][23][10] = (sum_out[9][23][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][23][10] = (sum_out[10][23][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][23][10] = (sum_out[11][23][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][23][10] = (sum_out[12][23][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][23][10] = (sum_out[13][23][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][23][10] = (sum_out[14][23][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][23][10] = (sum_out[15][23][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][23][10] = (sum_out[16][23][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][23][10] = (sum_out[17][23][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][23][10] = (sum_out[18][23][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][23][10] = (sum_out[19][23][10] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][23][11] = (sum_out[0][23][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][23][11] = (sum_out[1][23][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][23][11] = (sum_out[2][23][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][23][11] = (sum_out[3][23][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][23][11] = (sum_out[4][23][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][23][11] = (sum_out[5][23][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][23][11] = (sum_out[6][23][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][23][11] = (sum_out[7][23][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][23][11] = (sum_out[8][23][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][23][11] = (sum_out[9][23][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][23][11] = (sum_out[10][23][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][23][11] = (sum_out[11][23][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][23][11] = (sum_out[12][23][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][23][11] = (sum_out[13][23][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][23][11] = (sum_out[14][23][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][23][11] = (sum_out[15][23][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][23][11] = (sum_out[16][23][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][23][11] = (sum_out[17][23][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][23][11] = (sum_out[18][23][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][23][11] = (sum_out[19][23][11] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][23][12] = (sum_out[0][23][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][23][12] = (sum_out[1][23][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][23][12] = (sum_out[2][23][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][23][12] = (sum_out[3][23][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][23][12] = (sum_out[4][23][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][23][12] = (sum_out[5][23][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][23][12] = (sum_out[6][23][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][23][12] = (sum_out[7][23][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][23][12] = (sum_out[8][23][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][23][12] = (sum_out[9][23][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][23][12] = (sum_out[10][23][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][23][12] = (sum_out[11][23][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][23][12] = (sum_out[12][23][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][23][12] = (sum_out[13][23][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][23][12] = (sum_out[14][23][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][23][12] = (sum_out[15][23][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][23][12] = (sum_out[16][23][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][23][12] = (sum_out[17][23][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][23][12] = (sum_out[18][23][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][23][12] = (sum_out[19][23][12] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][23][13] = (sum_out[0][23][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][23][13] = (sum_out[1][23][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][23][13] = (sum_out[2][23][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][23][13] = (sum_out[3][23][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][23][13] = (sum_out[4][23][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][23][13] = (sum_out[5][23][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][23][13] = (sum_out[6][23][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][23][13] = (sum_out[7][23][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][23][13] = (sum_out[8][23][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][23][13] = (sum_out[9][23][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][23][13] = (sum_out[10][23][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][23][13] = (sum_out[11][23][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][23][13] = (sum_out[12][23][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][23][13] = (sum_out[13][23][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][23][13] = (sum_out[14][23][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][23][13] = (sum_out[15][23][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][23][13] = (sum_out[16][23][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][23][13] = (sum_out[17][23][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][23][13] = (sum_out[18][23][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][23][13] = (sum_out[19][23][13] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][23][14] = (sum_out[0][23][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][23][14] = (sum_out[1][23][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][23][14] = (sum_out[2][23][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][23][14] = (sum_out[3][23][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][23][14] = (sum_out[4][23][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][23][14] = (sum_out[5][23][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][23][14] = (sum_out[6][23][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][23][14] = (sum_out[7][23][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][23][14] = (sum_out[8][23][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][23][14] = (sum_out[9][23][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][23][14] = (sum_out[10][23][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][23][14] = (sum_out[11][23][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][23][14] = (sum_out[12][23][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][23][14] = (sum_out[13][23][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][23][14] = (sum_out[14][23][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][23][14] = (sum_out[15][23][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][23][14] = (sum_out[16][23][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][23][14] = (sum_out[17][23][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][23][14] = (sum_out[18][23][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][23][14] = (sum_out[19][23][14] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][23][15] = (sum_out[0][23][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][23][15] = (sum_out[1][23][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][23][15] = (sum_out[2][23][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][23][15] = (sum_out[3][23][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][23][15] = (sum_out[4][23][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][23][15] = (sum_out[5][23][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][23][15] = (sum_out[6][23][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][23][15] = (sum_out[7][23][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][23][15] = (sum_out[8][23][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][23][15] = (sum_out[9][23][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][23][15] = (sum_out[10][23][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][23][15] = (sum_out[11][23][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][23][15] = (sum_out[12][23][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][23][15] = (sum_out[13][23][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][23][15] = (sum_out[14][23][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][23][15] = (sum_out[15][23][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][23][15] = (sum_out[16][23][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][23][15] = (sum_out[17][23][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][23][15] = (sum_out[18][23][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][23][15] = (sum_out[19][23][15] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][23][16] = (sum_out[0][23][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][23][16] = (sum_out[1][23][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][23][16] = (sum_out[2][23][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][23][16] = (sum_out[3][23][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][23][16] = (sum_out[4][23][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][23][16] = (sum_out[5][23][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][23][16] = (sum_out[6][23][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][23][16] = (sum_out[7][23][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][23][16] = (sum_out[8][23][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][23][16] = (sum_out[9][23][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][23][16] = (sum_out[10][23][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][23][16] = (sum_out[11][23][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][23][16] = (sum_out[12][23][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][23][16] = (sum_out[13][23][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][23][16] = (sum_out[14][23][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][23][16] = (sum_out[15][23][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][23][16] = (sum_out[16][23][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][23][16] = (sum_out[17][23][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][23][16] = (sum_out[18][23][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][23][16] = (sum_out[19][23][16] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][23][17] = (sum_out[0][23][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][23][17] = (sum_out[1][23][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][23][17] = (sum_out[2][23][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][23][17] = (sum_out[3][23][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][23][17] = (sum_out[4][23][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][23][17] = (sum_out[5][23][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][23][17] = (sum_out[6][23][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][23][17] = (sum_out[7][23][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][23][17] = (sum_out[8][23][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][23][17] = (sum_out[9][23][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][23][17] = (sum_out[10][23][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][23][17] = (sum_out[11][23][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][23][17] = (sum_out[12][23][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][23][17] = (sum_out[13][23][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][23][17] = (sum_out[14][23][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][23][17] = (sum_out[15][23][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][23][17] = (sum_out[16][23][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][23][17] = (sum_out[17][23][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][23][17] = (sum_out[18][23][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][23][17] = (sum_out[19][23][17] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][23][18] = (sum_out[0][23][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][23][18] = (sum_out[1][23][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][23][18] = (sum_out[2][23][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][23][18] = (sum_out[3][23][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][23][18] = (sum_out[4][23][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][23][18] = (sum_out[5][23][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][23][18] = (sum_out[6][23][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][23][18] = (sum_out[7][23][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][23][18] = (sum_out[8][23][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][23][18] = (sum_out[9][23][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][23][18] = (sum_out[10][23][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][23][18] = (sum_out[11][23][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][23][18] = (sum_out[12][23][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][23][18] = (sum_out[13][23][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][23][18] = (sum_out[14][23][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][23][18] = (sum_out[15][23][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][23][18] = (sum_out[16][23][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][23][18] = (sum_out[17][23][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][23][18] = (sum_out[18][23][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][23][18] = (sum_out[19][23][18] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][23][19] = (sum_out[0][23][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][23][19] = (sum_out[1][23][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][23][19] = (sum_out[2][23][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][23][19] = (sum_out[3][23][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][23][19] = (sum_out[4][23][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][23][19] = (sum_out[5][23][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][23][19] = (sum_out[6][23][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][23][19] = (sum_out[7][23][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][23][19] = (sum_out[8][23][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][23][19] = (sum_out[9][23][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][23][19] = (sum_out[10][23][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][23][19] = (sum_out[11][23][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][23][19] = (sum_out[12][23][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][23][19] = (sum_out[13][23][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][23][19] = (sum_out[14][23][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][23][19] = (sum_out[15][23][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][23][19] = (sum_out[16][23][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][23][19] = (sum_out[17][23][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][23][19] = (sum_out[18][23][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][23][19] = (sum_out[19][23][19] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][23][20] = (sum_out[0][23][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][23][20] = (sum_out[1][23][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][23][20] = (sum_out[2][23][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][23][20] = (sum_out[3][23][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][23][20] = (sum_out[4][23][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][23][20] = (sum_out[5][23][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][23][20] = (sum_out[6][23][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][23][20] = (sum_out[7][23][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][23][20] = (sum_out[8][23][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][23][20] = (sum_out[9][23][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][23][20] = (sum_out[10][23][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][23][20] = (sum_out[11][23][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][23][20] = (sum_out[12][23][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][23][20] = (sum_out[13][23][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][23][20] = (sum_out[14][23][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][23][20] = (sum_out[15][23][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][23][20] = (sum_out[16][23][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][23][20] = (sum_out[17][23][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][23][20] = (sum_out[18][23][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][23][20] = (sum_out[19][23][20] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][23][21] = (sum_out[0][23][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][23][21] = (sum_out[1][23][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][23][21] = (sum_out[2][23][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][23][21] = (sum_out[3][23][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][23][21] = (sum_out[4][23][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][23][21] = (sum_out[5][23][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][23][21] = (sum_out[6][23][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][23][21] = (sum_out[7][23][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][23][21] = (sum_out[8][23][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][23][21] = (sum_out[9][23][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][23][21] = (sum_out[10][23][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][23][21] = (sum_out[11][23][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][23][21] = (sum_out[12][23][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][23][21] = (sum_out[13][23][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][23][21] = (sum_out[14][23][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][23][21] = (sum_out[15][23][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][23][21] = (sum_out[16][23][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][23][21] = (sum_out[17][23][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][23][21] = (sum_out[18][23][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][23][21] = (sum_out[19][23][21] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][23][22] = (sum_out[0][23][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][23][22] = (sum_out[1][23][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][23][22] = (sum_out[2][23][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][23][22] = (sum_out[3][23][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][23][22] = (sum_out[4][23][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][23][22] = (sum_out[5][23][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][23][22] = (sum_out[6][23][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][23][22] = (sum_out[7][23][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][23][22] = (sum_out[8][23][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][23][22] = (sum_out[9][23][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][23][22] = (sum_out[10][23][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][23][22] = (sum_out[11][23][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][23][22] = (sum_out[12][23][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][23][22] = (sum_out[13][23][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][23][22] = (sum_out[14][23][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][23][22] = (sum_out[15][23][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][23][22] = (sum_out[16][23][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][23][22] = (sum_out[17][23][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][23][22] = (sum_out[18][23][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][23][22] = (sum_out[19][23][22] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[0][23][23] = (sum_out[0][23][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[1][23][23] = (sum_out[1][23][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[2][23][23] = (sum_out[2][23][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[3][23][23] = (sum_out[3][23][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[4][23][23] = (sum_out[4][23][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[5][23][23] = (sum_out[5][23][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[6][23][23] = (sum_out[6][23][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[7][23][23] = (sum_out[7][23][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[8][23][23] = (sum_out[8][23][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[9][23][23] = (sum_out[9][23][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[10][23][23] = (sum_out[10][23][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[11][23][23] = (sum_out[11][23][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[12][23][23] = (sum_out[12][23][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[13][23][23] = (sum_out[13][23][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[14][23][23] = (sum_out[14][23][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[15][23][23] = (sum_out[15][23][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[16][23][23] = (sum_out[16][23][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[17][23][23] = (sum_out[17][23][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[18][23][23] = (sum_out[18][23][23] >= 3'b011) ? 1'b1: 1'b0;
assign conv_one_out[19][23][23] = (sum_out[19][23][23] >= 3'b011) ? 1'b1: 1'b0;

endmodule