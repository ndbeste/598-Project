module fully_connected 
	#( parameter bW = 8,
	   parameter fI = 960, // Fan in
	   parameter sW = 10) // Sum width -> clog2(fI)
(
    input  logic clk,
    input  logic rst_n,
    input  logic fc_valid,
    output logic sum_valid,
    input  logic [fI-1   :0] fan_in,
    input  logic [bW-1   :0] weights        [0:9],
    input  logic [fI-1   :0] binary_weights [0:9],
    output logic [bW+sW-2:0] fan_out        [0:9]
);

    logic [fI-1:0] xnor_result              [0:9]; // will store 0/1 strings for all output nodes
    logic [sW-1:0] accumulation_result      [0:9]; // will store total # of 1's observed
    logic [sW-1:0] accumulation_after_bias  [0:9]; // will store total # of 1's - fI/2 -> which is like (x*2 - 960)/2 observed

    logic processing; // lazy way - shift register as we know it takes only 2 cycles
    always_ff @(posedge clk) begin
      if (~rst_n) begin
         processing <= 1'b0;
      end else begin
         processing <= fc_valid;
      end
    end

    always_ff @(posedge clk) begin
      if (~rst_n) begin
         sum_valid <= 1'b0;
      end else begin
         sum_valid <= processing;
      end
    end

assign xnor_result[0] = (binary_weights[0] ~^ fan_in);
assign xnor_result[1] = (binary_weights[1] ~^ fan_in);
assign xnor_result[2] = (binary_weights[2] ~^ fan_in);
assign xnor_result[3] = (binary_weights[3] ~^ fan_in);
assign xnor_result[4] = (binary_weights[4] ~^ fan_in);
assign xnor_result[5] = (binary_weights[5] ~^ fan_in);
assign xnor_result[6] = (binary_weights[6] ~^ fan_in);
assign xnor_result[7] = (binary_weights[7] ~^ fan_in);
assign xnor_result[8] = (binary_weights[8] ~^ fan_in);
assign xnor_result[9] = (binary_weights[9] ~^ fan_in);
assign accumulation_result[0] = xnor_result[0][0] + xnor_result[0][1] + xnor_result[0][2] + xnor_result[0][3] + xnor_result[0][4] + xnor_result[0][5] + xnor_result[0][6] + xnor_result[0][7] + xnor_result[0][8] + xnor_result[0][9] + xnor_result[0][10] + xnor_result[0][11] + xnor_result[0][12] + xnor_result[0][13] + xnor_result[0][14] + xnor_result[0][15] + xnor_result[0][16] + xnor_result[0][17] + xnor_result[0][18] + xnor_result[0][19] + xnor_result[0][20] + xnor_result[0][21] + xnor_result[0][22] + xnor_result[0][23] + xnor_result[0][24] + xnor_result[0][25] + xnor_result[0][26] + xnor_result[0][27] + xnor_result[0][28] + xnor_result[0][29] + xnor_result[0][30] + xnor_result[0][31] + xnor_result[0][32] + xnor_result[0][33] + xnor_result[0][34] + xnor_result[0][35] + xnor_result[0][36] + xnor_result[0][37] + xnor_result[0][38] + xnor_result[0][39] + xnor_result[0][40] + xnor_result[0][41] + xnor_result[0][42] + xnor_result[0][43] + xnor_result[0][44] + xnor_result[0][45] + xnor_result[0][46] + xnor_result[0][47] + xnor_result[0][48] + xnor_result[0][49] + xnor_result[0][50] + xnor_result[0][51] + xnor_result[0][52] + xnor_result[0][53] + xnor_result[0][54] + xnor_result[0][55] + xnor_result[0][56] + xnor_result[0][57] + xnor_result[0][58] + xnor_result[0][59] + xnor_result[0][60] + xnor_result[0][61] + xnor_result[0][62] + xnor_result[0][63] + xnor_result[0][64] + xnor_result[0][65] + xnor_result[0][66] + xnor_result[0][67] + xnor_result[0][68] + xnor_result[0][69] + xnor_result[0][70] + xnor_result[0][71] + xnor_result[0][72] + xnor_result[0][73] + xnor_result[0][74] + xnor_result[0][75] + xnor_result[0][76] + xnor_result[0][77] + xnor_result[0][78] + xnor_result[0][79] + xnor_result[0][80] + xnor_result[0][81] + xnor_result[0][82] + xnor_result[0][83] + xnor_result[0][84] + xnor_result[0][85] + xnor_result[0][86] + xnor_result[0][87] + xnor_result[0][88] + xnor_result[0][89] + xnor_result[0][90] + xnor_result[0][91] + xnor_result[0][92] + xnor_result[0][93] + xnor_result[0][94] + xnor_result[0][95] + xnor_result[0][96] + xnor_result[0][97] + xnor_result[0][98] + xnor_result[0][99] + xnor_result[0][100] + xnor_result[0][101] + xnor_result[0][102] + xnor_result[0][103] + xnor_result[0][104] + xnor_result[0][105] + xnor_result[0][106] + xnor_result[0][107] + xnor_result[0][108] + xnor_result[0][109] + xnor_result[0][110] + xnor_result[0][111] + xnor_result[0][112] + xnor_result[0][113] + xnor_result[0][114] + xnor_result[0][115] + xnor_result[0][116] + xnor_result[0][117] + xnor_result[0][118] + xnor_result[0][119] + xnor_result[0][120] + xnor_result[0][121] + xnor_result[0][122] + xnor_result[0][123] + xnor_result[0][124] + xnor_result[0][125] + xnor_result[0][126] + xnor_result[0][127] + xnor_result[0][128] + xnor_result[0][129] + xnor_result[0][130] + xnor_result[0][131] + xnor_result[0][132] + xnor_result[0][133] + xnor_result[0][134] + xnor_result[0][135] + xnor_result[0][136] + xnor_result[0][137] + xnor_result[0][138] + xnor_result[0][139] + xnor_result[0][140] + xnor_result[0][141] + xnor_result[0][142] + xnor_result[0][143] + xnor_result[0][144] + xnor_result[0][145] + xnor_result[0][146] + xnor_result[0][147] + xnor_result[0][148] + xnor_result[0][149] + xnor_result[0][150] + xnor_result[0][151] + xnor_result[0][152] + xnor_result[0][153] + xnor_result[0][154] + xnor_result[0][155] + xnor_result[0][156] + xnor_result[0][157] + xnor_result[0][158] + xnor_result[0][159] + xnor_result[0][160] + xnor_result[0][161] + xnor_result[0][162] + xnor_result[0][163] + xnor_result[0][164] + xnor_result[0][165] + xnor_result[0][166] + xnor_result[0][167] + xnor_result[0][168] + xnor_result[0][169] + xnor_result[0][170] + xnor_result[0][171] + xnor_result[0][172] + xnor_result[0][173] + xnor_result[0][174] + xnor_result[0][175] + xnor_result[0][176] + xnor_result[0][177] + xnor_result[0][178] + xnor_result[0][179] + xnor_result[0][180] + xnor_result[0][181] + xnor_result[0][182] + xnor_result[0][183] + xnor_result[0][184] + xnor_result[0][185] + xnor_result[0][186] + xnor_result[0][187] + xnor_result[0][188] + xnor_result[0][189] + xnor_result[0][190] + xnor_result[0][191] + xnor_result[0][192] + xnor_result[0][193] + xnor_result[0][194] + xnor_result[0][195] + xnor_result[0][196] + xnor_result[0][197] + xnor_result[0][198] + xnor_result[0][199] + xnor_result[0][200] + xnor_result[0][201] + xnor_result[0][202] + xnor_result[0][203] + xnor_result[0][204] + xnor_result[0][205] + xnor_result[0][206] + xnor_result[0][207] + xnor_result[0][208] + xnor_result[0][209] + xnor_result[0][210] + xnor_result[0][211] + xnor_result[0][212] + xnor_result[0][213] + xnor_result[0][214] + xnor_result[0][215] + xnor_result[0][216] + xnor_result[0][217] + xnor_result[0][218] + xnor_result[0][219] + xnor_result[0][220] + xnor_result[0][221] + xnor_result[0][222] + xnor_result[0][223] + xnor_result[0][224] + xnor_result[0][225] + xnor_result[0][226] + xnor_result[0][227] + xnor_result[0][228] + xnor_result[0][229] + xnor_result[0][230] + xnor_result[0][231] + xnor_result[0][232] + xnor_result[0][233] + xnor_result[0][234] + xnor_result[0][235] + xnor_result[0][236] + xnor_result[0][237] + xnor_result[0][238] + xnor_result[0][239] + xnor_result[0][240] + xnor_result[0][241] + xnor_result[0][242] + xnor_result[0][243] + xnor_result[0][244] + xnor_result[0][245] + xnor_result[0][246] + xnor_result[0][247] + xnor_result[0][248] + xnor_result[0][249] + xnor_result[0][250] + xnor_result[0][251] + xnor_result[0][252] + xnor_result[0][253] + xnor_result[0][254] + xnor_result[0][255] + xnor_result[0][256] + xnor_result[0][257] + xnor_result[0][258] + xnor_result[0][259] + xnor_result[0][260] + xnor_result[0][261] + xnor_result[0][262] + xnor_result[0][263] + xnor_result[0][264] + xnor_result[0][265] + xnor_result[0][266] + xnor_result[0][267] + xnor_result[0][268] + xnor_result[0][269] + xnor_result[0][270] + xnor_result[0][271] + xnor_result[0][272] + xnor_result[0][273] + xnor_result[0][274] + xnor_result[0][275] + xnor_result[0][276] + xnor_result[0][277] + xnor_result[0][278] + xnor_result[0][279] + xnor_result[0][280] + xnor_result[0][281] + xnor_result[0][282] + xnor_result[0][283] + xnor_result[0][284] + xnor_result[0][285] + xnor_result[0][286] + xnor_result[0][287] + xnor_result[0][288] + xnor_result[0][289] + xnor_result[0][290] + xnor_result[0][291] + xnor_result[0][292] + xnor_result[0][293] + xnor_result[0][294] + xnor_result[0][295] + xnor_result[0][296] + xnor_result[0][297] + xnor_result[0][298] + xnor_result[0][299] + xnor_result[0][300] + xnor_result[0][301] + xnor_result[0][302] + xnor_result[0][303] + xnor_result[0][304] + xnor_result[0][305] + xnor_result[0][306] + xnor_result[0][307] + xnor_result[0][308] + xnor_result[0][309] + xnor_result[0][310] + xnor_result[0][311] + xnor_result[0][312] + xnor_result[0][313] + xnor_result[0][314] + xnor_result[0][315] + xnor_result[0][316] + xnor_result[0][317] + xnor_result[0][318] + xnor_result[0][319] + xnor_result[0][320] + xnor_result[0][321] + xnor_result[0][322] + xnor_result[0][323] + xnor_result[0][324] + xnor_result[0][325] + xnor_result[0][326] + xnor_result[0][327] + xnor_result[0][328] + xnor_result[0][329] + xnor_result[0][330] + xnor_result[0][331] + xnor_result[0][332] + xnor_result[0][333] + xnor_result[0][334] + xnor_result[0][335] + xnor_result[0][336] + xnor_result[0][337] + xnor_result[0][338] + xnor_result[0][339] + xnor_result[0][340] + xnor_result[0][341] + xnor_result[0][342] + xnor_result[0][343] + xnor_result[0][344] + xnor_result[0][345] + xnor_result[0][346] + xnor_result[0][347] + xnor_result[0][348] + xnor_result[0][349] + xnor_result[0][350] + xnor_result[0][351] + xnor_result[0][352] + xnor_result[0][353] + xnor_result[0][354] + xnor_result[0][355] + xnor_result[0][356] + xnor_result[0][357] + xnor_result[0][358] + xnor_result[0][359] + xnor_result[0][360] + xnor_result[0][361] + xnor_result[0][362] + xnor_result[0][363] + xnor_result[0][364] + xnor_result[0][365] + xnor_result[0][366] + xnor_result[0][367] + xnor_result[0][368] + xnor_result[0][369] + xnor_result[0][370] + xnor_result[0][371] + xnor_result[0][372] + xnor_result[0][373] + xnor_result[0][374] + xnor_result[0][375] + xnor_result[0][376] + xnor_result[0][377] + xnor_result[0][378] + xnor_result[0][379] + xnor_result[0][380] + xnor_result[0][381] + xnor_result[0][382] + xnor_result[0][383] + xnor_result[0][384] + xnor_result[0][385] + xnor_result[0][386] + xnor_result[0][387] + xnor_result[0][388] + xnor_result[0][389] + xnor_result[0][390] + xnor_result[0][391] + xnor_result[0][392] + xnor_result[0][393] + xnor_result[0][394] + xnor_result[0][395] + xnor_result[0][396] + xnor_result[0][397] + xnor_result[0][398] + xnor_result[0][399] + xnor_result[0][400] + xnor_result[0][401] + xnor_result[0][402] + xnor_result[0][403] + xnor_result[0][404] + xnor_result[0][405] + xnor_result[0][406] + xnor_result[0][407] + xnor_result[0][408] + xnor_result[0][409] + xnor_result[0][410] + xnor_result[0][411] + xnor_result[0][412] + xnor_result[0][413] + xnor_result[0][414] + xnor_result[0][415] + xnor_result[0][416] + xnor_result[0][417] + xnor_result[0][418] + xnor_result[0][419] + xnor_result[0][420] + xnor_result[0][421] + xnor_result[0][422] + xnor_result[0][423] + xnor_result[0][424] + xnor_result[0][425] + xnor_result[0][426] + xnor_result[0][427] + xnor_result[0][428] + xnor_result[0][429] + xnor_result[0][430] + xnor_result[0][431] + xnor_result[0][432] + xnor_result[0][433] + xnor_result[0][434] + xnor_result[0][435] + xnor_result[0][436] + xnor_result[0][437] + xnor_result[0][438] + xnor_result[0][439] + xnor_result[0][440] + xnor_result[0][441] + xnor_result[0][442] + xnor_result[0][443] + xnor_result[0][444] + xnor_result[0][445] + xnor_result[0][446] + xnor_result[0][447] + xnor_result[0][448] + xnor_result[0][449] + xnor_result[0][450] + xnor_result[0][451] + xnor_result[0][452] + xnor_result[0][453] + xnor_result[0][454] + xnor_result[0][455] + xnor_result[0][456] + xnor_result[0][457] + xnor_result[0][458] + xnor_result[0][459] + xnor_result[0][460] + xnor_result[0][461] + xnor_result[0][462] + xnor_result[0][463] + xnor_result[0][464] + xnor_result[0][465] + xnor_result[0][466] + xnor_result[0][467] + xnor_result[0][468] + xnor_result[0][469] + xnor_result[0][470] + xnor_result[0][471] + xnor_result[0][472] + xnor_result[0][473] + xnor_result[0][474] + xnor_result[0][475] + xnor_result[0][476] + xnor_result[0][477] + xnor_result[0][478] + xnor_result[0][479] + xnor_result[0][480] + xnor_result[0][481] + xnor_result[0][482] + xnor_result[0][483] + xnor_result[0][484] + xnor_result[0][485] + xnor_result[0][486] + xnor_result[0][487] + xnor_result[0][488] + xnor_result[0][489] + xnor_result[0][490] + xnor_result[0][491] + xnor_result[0][492] + xnor_result[0][493] + xnor_result[0][494] + xnor_result[0][495] + xnor_result[0][496] + xnor_result[0][497] + xnor_result[0][498] + xnor_result[0][499] + xnor_result[0][500] + xnor_result[0][501] + xnor_result[0][502] + xnor_result[0][503] + xnor_result[0][504] + xnor_result[0][505] + xnor_result[0][506] + xnor_result[0][507] + xnor_result[0][508] + xnor_result[0][509] + xnor_result[0][510] + xnor_result[0][511] + xnor_result[0][512] + xnor_result[0][513] + xnor_result[0][514] + xnor_result[0][515] + xnor_result[0][516] + xnor_result[0][517] + xnor_result[0][518] + xnor_result[0][519] + xnor_result[0][520] + xnor_result[0][521] + xnor_result[0][522] + xnor_result[0][523] + xnor_result[0][524] + xnor_result[0][525] + xnor_result[0][526] + xnor_result[0][527] + xnor_result[0][528] + xnor_result[0][529] + xnor_result[0][530] + xnor_result[0][531] + xnor_result[0][532] + xnor_result[0][533] + xnor_result[0][534] + xnor_result[0][535] + xnor_result[0][536] + xnor_result[0][537] + xnor_result[0][538] + xnor_result[0][539] + xnor_result[0][540] + xnor_result[0][541] + xnor_result[0][542] + xnor_result[0][543] + xnor_result[0][544] + xnor_result[0][545] + xnor_result[0][546] + xnor_result[0][547] + xnor_result[0][548] + xnor_result[0][549] + xnor_result[0][550] + xnor_result[0][551] + xnor_result[0][552] + xnor_result[0][553] + xnor_result[0][554] + xnor_result[0][555] + xnor_result[0][556] + xnor_result[0][557] + xnor_result[0][558] + xnor_result[0][559] + xnor_result[0][560] + xnor_result[0][561] + xnor_result[0][562] + xnor_result[0][563] + xnor_result[0][564] + xnor_result[0][565] + xnor_result[0][566] + xnor_result[0][567] + xnor_result[0][568] + xnor_result[0][569] + xnor_result[0][570] + xnor_result[0][571] + xnor_result[0][572] + xnor_result[0][573] + xnor_result[0][574] + xnor_result[0][575] + xnor_result[0][576] + xnor_result[0][577] + xnor_result[0][578] + xnor_result[0][579] + xnor_result[0][580] + xnor_result[0][581] + xnor_result[0][582] + xnor_result[0][583] + xnor_result[0][584] + xnor_result[0][585] + xnor_result[0][586] + xnor_result[0][587] + xnor_result[0][588] + xnor_result[0][589] + xnor_result[0][590] + xnor_result[0][591] + xnor_result[0][592] + xnor_result[0][593] + xnor_result[0][594] + xnor_result[0][595] + xnor_result[0][596] + xnor_result[0][597] + xnor_result[0][598] + xnor_result[0][599] + xnor_result[0][600] + xnor_result[0][601] + xnor_result[0][602] + xnor_result[0][603] + xnor_result[0][604] + xnor_result[0][605] + xnor_result[0][606] + xnor_result[0][607] + xnor_result[0][608] + xnor_result[0][609] + xnor_result[0][610] + xnor_result[0][611] + xnor_result[0][612] + xnor_result[0][613] + xnor_result[0][614] + xnor_result[0][615] + xnor_result[0][616] + xnor_result[0][617] + xnor_result[0][618] + xnor_result[0][619] + xnor_result[0][620] + xnor_result[0][621] + xnor_result[0][622] + xnor_result[0][623] + xnor_result[0][624] + xnor_result[0][625] + xnor_result[0][626] + xnor_result[0][627] + xnor_result[0][628] + xnor_result[0][629] + xnor_result[0][630] + xnor_result[0][631] + xnor_result[0][632] + xnor_result[0][633] + xnor_result[0][634] + xnor_result[0][635] + xnor_result[0][636] + xnor_result[0][637] + xnor_result[0][638] + xnor_result[0][639] + xnor_result[0][640] + xnor_result[0][641] + xnor_result[0][642] + xnor_result[0][643] + xnor_result[0][644] + xnor_result[0][645] + xnor_result[0][646] + xnor_result[0][647] + xnor_result[0][648] + xnor_result[0][649] + xnor_result[0][650] + xnor_result[0][651] + xnor_result[0][652] + xnor_result[0][653] + xnor_result[0][654] + xnor_result[0][655] + xnor_result[0][656] + xnor_result[0][657] + xnor_result[0][658] + xnor_result[0][659] + xnor_result[0][660] + xnor_result[0][661] + xnor_result[0][662] + xnor_result[0][663] + xnor_result[0][664] + xnor_result[0][665] + xnor_result[0][666] + xnor_result[0][667] + xnor_result[0][668] + xnor_result[0][669] + xnor_result[0][670] + xnor_result[0][671] + xnor_result[0][672] + xnor_result[0][673] + xnor_result[0][674] + xnor_result[0][675] + xnor_result[0][676] + xnor_result[0][677] + xnor_result[0][678] + xnor_result[0][679] + xnor_result[0][680] + xnor_result[0][681] + xnor_result[0][682] + xnor_result[0][683] + xnor_result[0][684] + xnor_result[0][685] + xnor_result[0][686] + xnor_result[0][687] + xnor_result[0][688] + xnor_result[0][689] + xnor_result[0][690] + xnor_result[0][691] + xnor_result[0][692] + xnor_result[0][693] + xnor_result[0][694] + xnor_result[0][695] + xnor_result[0][696] + xnor_result[0][697] + xnor_result[0][698] + xnor_result[0][699] + xnor_result[0][700] + xnor_result[0][701] + xnor_result[0][702] + xnor_result[0][703] + xnor_result[0][704] + xnor_result[0][705] + xnor_result[0][706] + xnor_result[0][707] + xnor_result[0][708] + xnor_result[0][709] + xnor_result[0][710] + xnor_result[0][711] + xnor_result[0][712] + xnor_result[0][713] + xnor_result[0][714] + xnor_result[0][715] + xnor_result[0][716] + xnor_result[0][717] + xnor_result[0][718] + xnor_result[0][719] + xnor_result[0][720] + xnor_result[0][721] + xnor_result[0][722] + xnor_result[0][723] + xnor_result[0][724] + xnor_result[0][725] + xnor_result[0][726] + xnor_result[0][727] + xnor_result[0][728] + xnor_result[0][729] + xnor_result[0][730] + xnor_result[0][731] + xnor_result[0][732] + xnor_result[0][733] + xnor_result[0][734] + xnor_result[0][735] + xnor_result[0][736] + xnor_result[0][737] + xnor_result[0][738] + xnor_result[0][739] + xnor_result[0][740] + xnor_result[0][741] + xnor_result[0][742] + xnor_result[0][743] + xnor_result[0][744] + xnor_result[0][745] + xnor_result[0][746] + xnor_result[0][747] + xnor_result[0][748] + xnor_result[0][749] + xnor_result[0][750] + xnor_result[0][751] + xnor_result[0][752] + xnor_result[0][753] + xnor_result[0][754] + xnor_result[0][755] + xnor_result[0][756] + xnor_result[0][757] + xnor_result[0][758] + xnor_result[0][759] + xnor_result[0][760] + xnor_result[0][761] + xnor_result[0][762] + xnor_result[0][763] + xnor_result[0][764] + xnor_result[0][765] + xnor_result[0][766] + xnor_result[0][767] + xnor_result[0][768] + xnor_result[0][769] + xnor_result[0][770] + xnor_result[0][771] + xnor_result[0][772] + xnor_result[0][773] + xnor_result[0][774] + xnor_result[0][775] + xnor_result[0][776] + xnor_result[0][777] + xnor_result[0][778] + xnor_result[0][779] + xnor_result[0][780] + xnor_result[0][781] + xnor_result[0][782] + xnor_result[0][783] + xnor_result[0][784] + xnor_result[0][785] + xnor_result[0][786] + xnor_result[0][787] + xnor_result[0][788] + xnor_result[0][789] + xnor_result[0][790] + xnor_result[0][791] + xnor_result[0][792] + xnor_result[0][793] + xnor_result[0][794] + xnor_result[0][795] + xnor_result[0][796] + xnor_result[0][797] + xnor_result[0][798] + xnor_result[0][799] + xnor_result[0][800] + xnor_result[0][801] + xnor_result[0][802] + xnor_result[0][803] + xnor_result[0][804] + xnor_result[0][805] + xnor_result[0][806] + xnor_result[0][807] + xnor_result[0][808] + xnor_result[0][809] + xnor_result[0][810] + xnor_result[0][811] + xnor_result[0][812] + xnor_result[0][813] + xnor_result[0][814] + xnor_result[0][815] + xnor_result[0][816] + xnor_result[0][817] + xnor_result[0][818] + xnor_result[0][819] + xnor_result[0][820] + xnor_result[0][821] + xnor_result[0][822] + xnor_result[0][823] + xnor_result[0][824] + xnor_result[0][825] + xnor_result[0][826] + xnor_result[0][827] + xnor_result[0][828] + xnor_result[0][829] + xnor_result[0][830] + xnor_result[0][831] + xnor_result[0][832] + xnor_result[0][833] + xnor_result[0][834] + xnor_result[0][835] + xnor_result[0][836] + xnor_result[0][837] + xnor_result[0][838] + xnor_result[0][839] + xnor_result[0][840] + xnor_result[0][841] + xnor_result[0][842] + xnor_result[0][843] + xnor_result[0][844] + xnor_result[0][845] + xnor_result[0][846] + xnor_result[0][847] + xnor_result[0][848] + xnor_result[0][849] + xnor_result[0][850] + xnor_result[0][851] + xnor_result[0][852] + xnor_result[0][853] + xnor_result[0][854] + xnor_result[0][855] + xnor_result[0][856] + xnor_result[0][857] + xnor_result[0][858] + xnor_result[0][859] + xnor_result[0][860] + xnor_result[0][861] + xnor_result[0][862] + xnor_result[0][863] + xnor_result[0][864] + xnor_result[0][865] + xnor_result[0][866] + xnor_result[0][867] + xnor_result[0][868] + xnor_result[0][869] + xnor_result[0][870] + xnor_result[0][871] + xnor_result[0][872] + xnor_result[0][873] + xnor_result[0][874] + xnor_result[0][875] + xnor_result[0][876] + xnor_result[0][877] + xnor_result[0][878] + xnor_result[0][879] + xnor_result[0][880] + xnor_result[0][881] + xnor_result[0][882] + xnor_result[0][883] + xnor_result[0][884] + xnor_result[0][885] + xnor_result[0][886] + xnor_result[0][887] + xnor_result[0][888] + xnor_result[0][889] + xnor_result[0][890] + xnor_result[0][891] + xnor_result[0][892] + xnor_result[0][893] + xnor_result[0][894] + xnor_result[0][895] + xnor_result[0][896] + xnor_result[0][897] + xnor_result[0][898] + xnor_result[0][899] + xnor_result[0][900] + xnor_result[0][901] + xnor_result[0][902] + xnor_result[0][903] + xnor_result[0][904] + xnor_result[0][905] + xnor_result[0][906] + xnor_result[0][907] + xnor_result[0][908] + xnor_result[0][909] + xnor_result[0][910] + xnor_result[0][911] + xnor_result[0][912] + xnor_result[0][913] + xnor_result[0][914] + xnor_result[0][915] + xnor_result[0][916] + xnor_result[0][917] + xnor_result[0][918] + xnor_result[0][919] + xnor_result[0][920] + xnor_result[0][921] + xnor_result[0][922] + xnor_result[0][923] + xnor_result[0][924] + xnor_result[0][925] + xnor_result[0][926] + xnor_result[0][927] + xnor_result[0][928] + xnor_result[0][929] + xnor_result[0][930] + xnor_result[0][931] + xnor_result[0][932] + xnor_result[0][933] + xnor_result[0][934] + xnor_result[0][935] + xnor_result[0][936] + xnor_result[0][937] + xnor_result[0][938] + xnor_result[0][939] + xnor_result[0][940] + xnor_result[0][941] + xnor_result[0][942] + xnor_result[0][943] + xnor_result[0][944] + xnor_result[0][945] + xnor_result[0][946] + xnor_result[0][947] + xnor_result[0][948] + xnor_result[0][949] + xnor_result[0][950] + xnor_result[0][951] + xnor_result[0][952] + xnor_result[0][953] + xnor_result[0][954] + xnor_result[0][955] + xnor_result[0][956] + xnor_result[0][957] + xnor_result[0][958] + xnor_result[0][959] ;
assign accumulation_result[1] = xnor_result[1][0] + xnor_result[1][1] + xnor_result[1][2] + xnor_result[1][3] + xnor_result[1][4] + xnor_result[1][5] + xnor_result[1][6] + xnor_result[1][7] + xnor_result[1][8] + xnor_result[1][9] + xnor_result[1][10] + xnor_result[1][11] + xnor_result[1][12] + xnor_result[1][13] + xnor_result[1][14] + xnor_result[1][15] + xnor_result[1][16] + xnor_result[1][17] + xnor_result[1][18] + xnor_result[1][19] + xnor_result[1][20] + xnor_result[1][21] + xnor_result[1][22] + xnor_result[1][23] + xnor_result[1][24] + xnor_result[1][25] + xnor_result[1][26] + xnor_result[1][27] + xnor_result[1][28] + xnor_result[1][29] + xnor_result[1][30] + xnor_result[1][31] + xnor_result[1][32] + xnor_result[1][33] + xnor_result[1][34] + xnor_result[1][35] + xnor_result[1][36] + xnor_result[1][37] + xnor_result[1][38] + xnor_result[1][39] + xnor_result[1][40] + xnor_result[1][41] + xnor_result[1][42] + xnor_result[1][43] + xnor_result[1][44] + xnor_result[1][45] + xnor_result[1][46] + xnor_result[1][47] + xnor_result[1][48] + xnor_result[1][49] + xnor_result[1][50] + xnor_result[1][51] + xnor_result[1][52] + xnor_result[1][53] + xnor_result[1][54] + xnor_result[1][55] + xnor_result[1][56] + xnor_result[1][57] + xnor_result[1][58] + xnor_result[1][59] + xnor_result[1][60] + xnor_result[1][61] + xnor_result[1][62] + xnor_result[1][63] + xnor_result[1][64] + xnor_result[1][65] + xnor_result[1][66] + xnor_result[1][67] + xnor_result[1][68] + xnor_result[1][69] + xnor_result[1][70] + xnor_result[1][71] + xnor_result[1][72] + xnor_result[1][73] + xnor_result[1][74] + xnor_result[1][75] + xnor_result[1][76] + xnor_result[1][77] + xnor_result[1][78] + xnor_result[1][79] + xnor_result[1][80] + xnor_result[1][81] + xnor_result[1][82] + xnor_result[1][83] + xnor_result[1][84] + xnor_result[1][85] + xnor_result[1][86] + xnor_result[1][87] + xnor_result[1][88] + xnor_result[1][89] + xnor_result[1][90] + xnor_result[1][91] + xnor_result[1][92] + xnor_result[1][93] + xnor_result[1][94] + xnor_result[1][95] + xnor_result[1][96] + xnor_result[1][97] + xnor_result[1][98] + xnor_result[1][99] + xnor_result[1][100] + xnor_result[1][101] + xnor_result[1][102] + xnor_result[1][103] + xnor_result[1][104] + xnor_result[1][105] + xnor_result[1][106] + xnor_result[1][107] + xnor_result[1][108] + xnor_result[1][109] + xnor_result[1][110] + xnor_result[1][111] + xnor_result[1][112] + xnor_result[1][113] + xnor_result[1][114] + xnor_result[1][115] + xnor_result[1][116] + xnor_result[1][117] + xnor_result[1][118] + xnor_result[1][119] + xnor_result[1][120] + xnor_result[1][121] + xnor_result[1][122] + xnor_result[1][123] + xnor_result[1][124] + xnor_result[1][125] + xnor_result[1][126] + xnor_result[1][127] + xnor_result[1][128] + xnor_result[1][129] + xnor_result[1][130] + xnor_result[1][131] + xnor_result[1][132] + xnor_result[1][133] + xnor_result[1][134] + xnor_result[1][135] + xnor_result[1][136] + xnor_result[1][137] + xnor_result[1][138] + xnor_result[1][139] + xnor_result[1][140] + xnor_result[1][141] + xnor_result[1][142] + xnor_result[1][143] + xnor_result[1][144] + xnor_result[1][145] + xnor_result[1][146] + xnor_result[1][147] + xnor_result[1][148] + xnor_result[1][149] + xnor_result[1][150] + xnor_result[1][151] + xnor_result[1][152] + xnor_result[1][153] + xnor_result[1][154] + xnor_result[1][155] + xnor_result[1][156] + xnor_result[1][157] + xnor_result[1][158] + xnor_result[1][159] + xnor_result[1][160] + xnor_result[1][161] + xnor_result[1][162] + xnor_result[1][163] + xnor_result[1][164] + xnor_result[1][165] + xnor_result[1][166] + xnor_result[1][167] + xnor_result[1][168] + xnor_result[1][169] + xnor_result[1][170] + xnor_result[1][171] + xnor_result[1][172] + xnor_result[1][173] + xnor_result[1][174] + xnor_result[1][175] + xnor_result[1][176] + xnor_result[1][177] + xnor_result[1][178] + xnor_result[1][179] + xnor_result[1][180] + xnor_result[1][181] + xnor_result[1][182] + xnor_result[1][183] + xnor_result[1][184] + xnor_result[1][185] + xnor_result[1][186] + xnor_result[1][187] + xnor_result[1][188] + xnor_result[1][189] + xnor_result[1][190] + xnor_result[1][191] + xnor_result[1][192] + xnor_result[1][193] + xnor_result[1][194] + xnor_result[1][195] + xnor_result[1][196] + xnor_result[1][197] + xnor_result[1][198] + xnor_result[1][199] + xnor_result[1][200] + xnor_result[1][201] + xnor_result[1][202] + xnor_result[1][203] + xnor_result[1][204] + xnor_result[1][205] + xnor_result[1][206] + xnor_result[1][207] + xnor_result[1][208] + xnor_result[1][209] + xnor_result[1][210] + xnor_result[1][211] + xnor_result[1][212] + xnor_result[1][213] + xnor_result[1][214] + xnor_result[1][215] + xnor_result[1][216] + xnor_result[1][217] + xnor_result[1][218] + xnor_result[1][219] + xnor_result[1][220] + xnor_result[1][221] + xnor_result[1][222] + xnor_result[1][223] + xnor_result[1][224] + xnor_result[1][225] + xnor_result[1][226] + xnor_result[1][227] + xnor_result[1][228] + xnor_result[1][229] + xnor_result[1][230] + xnor_result[1][231] + xnor_result[1][232] + xnor_result[1][233] + xnor_result[1][234] + xnor_result[1][235] + xnor_result[1][236] + xnor_result[1][237] + xnor_result[1][238] + xnor_result[1][239] + xnor_result[1][240] + xnor_result[1][241] + xnor_result[1][242] + xnor_result[1][243] + xnor_result[1][244] + xnor_result[1][245] + xnor_result[1][246] + xnor_result[1][247] + xnor_result[1][248] + xnor_result[1][249] + xnor_result[1][250] + xnor_result[1][251] + xnor_result[1][252] + xnor_result[1][253] + xnor_result[1][254] + xnor_result[1][255] + xnor_result[1][256] + xnor_result[1][257] + xnor_result[1][258] + xnor_result[1][259] + xnor_result[1][260] + xnor_result[1][261] + xnor_result[1][262] + xnor_result[1][263] + xnor_result[1][264] + xnor_result[1][265] + xnor_result[1][266] + xnor_result[1][267] + xnor_result[1][268] + xnor_result[1][269] + xnor_result[1][270] + xnor_result[1][271] + xnor_result[1][272] + xnor_result[1][273] + xnor_result[1][274] + xnor_result[1][275] + xnor_result[1][276] + xnor_result[1][277] + xnor_result[1][278] + xnor_result[1][279] + xnor_result[1][280] + xnor_result[1][281] + xnor_result[1][282] + xnor_result[1][283] + xnor_result[1][284] + xnor_result[1][285] + xnor_result[1][286] + xnor_result[1][287] + xnor_result[1][288] + xnor_result[1][289] + xnor_result[1][290] + xnor_result[1][291] + xnor_result[1][292] + xnor_result[1][293] + xnor_result[1][294] + xnor_result[1][295] + xnor_result[1][296] + xnor_result[1][297] + xnor_result[1][298] + xnor_result[1][299] + xnor_result[1][300] + xnor_result[1][301] + xnor_result[1][302] + xnor_result[1][303] + xnor_result[1][304] + xnor_result[1][305] + xnor_result[1][306] + xnor_result[1][307] + xnor_result[1][308] + xnor_result[1][309] + xnor_result[1][310] + xnor_result[1][311] + xnor_result[1][312] + xnor_result[1][313] + xnor_result[1][314] + xnor_result[1][315] + xnor_result[1][316] + xnor_result[1][317] + xnor_result[1][318] + xnor_result[1][319] + xnor_result[1][320] + xnor_result[1][321] + xnor_result[1][322] + xnor_result[1][323] + xnor_result[1][324] + xnor_result[1][325] + xnor_result[1][326] + xnor_result[1][327] + xnor_result[1][328] + xnor_result[1][329] + xnor_result[1][330] + xnor_result[1][331] + xnor_result[1][332] + xnor_result[1][333] + xnor_result[1][334] + xnor_result[1][335] + xnor_result[1][336] + xnor_result[1][337] + xnor_result[1][338] + xnor_result[1][339] + xnor_result[1][340] + xnor_result[1][341] + xnor_result[1][342] + xnor_result[1][343] + xnor_result[1][344] + xnor_result[1][345] + xnor_result[1][346] + xnor_result[1][347] + xnor_result[1][348] + xnor_result[1][349] + xnor_result[1][350] + xnor_result[1][351] + xnor_result[1][352] + xnor_result[1][353] + xnor_result[1][354] + xnor_result[1][355] + xnor_result[1][356] + xnor_result[1][357] + xnor_result[1][358] + xnor_result[1][359] + xnor_result[1][360] + xnor_result[1][361] + xnor_result[1][362] + xnor_result[1][363] + xnor_result[1][364] + xnor_result[1][365] + xnor_result[1][366] + xnor_result[1][367] + xnor_result[1][368] + xnor_result[1][369] + xnor_result[1][370] + xnor_result[1][371] + xnor_result[1][372] + xnor_result[1][373] + xnor_result[1][374] + xnor_result[1][375] + xnor_result[1][376] + xnor_result[1][377] + xnor_result[1][378] + xnor_result[1][379] + xnor_result[1][380] + xnor_result[1][381] + xnor_result[1][382] + xnor_result[1][383] + xnor_result[1][384] + xnor_result[1][385] + xnor_result[1][386] + xnor_result[1][387] + xnor_result[1][388] + xnor_result[1][389] + xnor_result[1][390] + xnor_result[1][391] + xnor_result[1][392] + xnor_result[1][393] + xnor_result[1][394] + xnor_result[1][395] + xnor_result[1][396] + xnor_result[1][397] + xnor_result[1][398] + xnor_result[1][399] + xnor_result[1][400] + xnor_result[1][401] + xnor_result[1][402] + xnor_result[1][403] + xnor_result[1][404] + xnor_result[1][405] + xnor_result[1][406] + xnor_result[1][407] + xnor_result[1][408] + xnor_result[1][409] + xnor_result[1][410] + xnor_result[1][411] + xnor_result[1][412] + xnor_result[1][413] + xnor_result[1][414] + xnor_result[1][415] + xnor_result[1][416] + xnor_result[1][417] + xnor_result[1][418] + xnor_result[1][419] + xnor_result[1][420] + xnor_result[1][421] + xnor_result[1][422] + xnor_result[1][423] + xnor_result[1][424] + xnor_result[1][425] + xnor_result[1][426] + xnor_result[1][427] + xnor_result[1][428] + xnor_result[1][429] + xnor_result[1][430] + xnor_result[1][431] + xnor_result[1][432] + xnor_result[1][433] + xnor_result[1][434] + xnor_result[1][435] + xnor_result[1][436] + xnor_result[1][437] + xnor_result[1][438] + xnor_result[1][439] + xnor_result[1][440] + xnor_result[1][441] + xnor_result[1][442] + xnor_result[1][443] + xnor_result[1][444] + xnor_result[1][445] + xnor_result[1][446] + xnor_result[1][447] + xnor_result[1][448] + xnor_result[1][449] + xnor_result[1][450] + xnor_result[1][451] + xnor_result[1][452] + xnor_result[1][453] + xnor_result[1][454] + xnor_result[1][455] + xnor_result[1][456] + xnor_result[1][457] + xnor_result[1][458] + xnor_result[1][459] + xnor_result[1][460] + xnor_result[1][461] + xnor_result[1][462] + xnor_result[1][463] + xnor_result[1][464] + xnor_result[1][465] + xnor_result[1][466] + xnor_result[1][467] + xnor_result[1][468] + xnor_result[1][469] + xnor_result[1][470] + xnor_result[1][471] + xnor_result[1][472] + xnor_result[1][473] + xnor_result[1][474] + xnor_result[1][475] + xnor_result[1][476] + xnor_result[1][477] + xnor_result[1][478] + xnor_result[1][479] + xnor_result[1][480] + xnor_result[1][481] + xnor_result[1][482] + xnor_result[1][483] + xnor_result[1][484] + xnor_result[1][485] + xnor_result[1][486] + xnor_result[1][487] + xnor_result[1][488] + xnor_result[1][489] + xnor_result[1][490] + xnor_result[1][491] + xnor_result[1][492] + xnor_result[1][493] + xnor_result[1][494] + xnor_result[1][495] + xnor_result[1][496] + xnor_result[1][497] + xnor_result[1][498] + xnor_result[1][499] + xnor_result[1][500] + xnor_result[1][501] + xnor_result[1][502] + xnor_result[1][503] + xnor_result[1][504] + xnor_result[1][505] + xnor_result[1][506] + xnor_result[1][507] + xnor_result[1][508] + xnor_result[1][509] + xnor_result[1][510] + xnor_result[1][511] + xnor_result[1][512] + xnor_result[1][513] + xnor_result[1][514] + xnor_result[1][515] + xnor_result[1][516] + xnor_result[1][517] + xnor_result[1][518] + xnor_result[1][519] + xnor_result[1][520] + xnor_result[1][521] + xnor_result[1][522] + xnor_result[1][523] + xnor_result[1][524] + xnor_result[1][525] + xnor_result[1][526] + xnor_result[1][527] + xnor_result[1][528] + xnor_result[1][529] + xnor_result[1][530] + xnor_result[1][531] + xnor_result[1][532] + xnor_result[1][533] + xnor_result[1][534] + xnor_result[1][535] + xnor_result[1][536] + xnor_result[1][537] + xnor_result[1][538] + xnor_result[1][539] + xnor_result[1][540] + xnor_result[1][541] + xnor_result[1][542] + xnor_result[1][543] + xnor_result[1][544] + xnor_result[1][545] + xnor_result[1][546] + xnor_result[1][547] + xnor_result[1][548] + xnor_result[1][549] + xnor_result[1][550] + xnor_result[1][551] + xnor_result[1][552] + xnor_result[1][553] + xnor_result[1][554] + xnor_result[1][555] + xnor_result[1][556] + xnor_result[1][557] + xnor_result[1][558] + xnor_result[1][559] + xnor_result[1][560] + xnor_result[1][561] + xnor_result[1][562] + xnor_result[1][563] + xnor_result[1][564] + xnor_result[1][565] + xnor_result[1][566] + xnor_result[1][567] + xnor_result[1][568] + xnor_result[1][569] + xnor_result[1][570] + xnor_result[1][571] + xnor_result[1][572] + xnor_result[1][573] + xnor_result[1][574] + xnor_result[1][575] + xnor_result[1][576] + xnor_result[1][577] + xnor_result[1][578] + xnor_result[1][579] + xnor_result[1][580] + xnor_result[1][581] + xnor_result[1][582] + xnor_result[1][583] + xnor_result[1][584] + xnor_result[1][585] + xnor_result[1][586] + xnor_result[1][587] + xnor_result[1][588] + xnor_result[1][589] + xnor_result[1][590] + xnor_result[1][591] + xnor_result[1][592] + xnor_result[1][593] + xnor_result[1][594] + xnor_result[1][595] + xnor_result[1][596] + xnor_result[1][597] + xnor_result[1][598] + xnor_result[1][599] + xnor_result[1][600] + xnor_result[1][601] + xnor_result[1][602] + xnor_result[1][603] + xnor_result[1][604] + xnor_result[1][605] + xnor_result[1][606] + xnor_result[1][607] + xnor_result[1][608] + xnor_result[1][609] + xnor_result[1][610] + xnor_result[1][611] + xnor_result[1][612] + xnor_result[1][613] + xnor_result[1][614] + xnor_result[1][615] + xnor_result[1][616] + xnor_result[1][617] + xnor_result[1][618] + xnor_result[1][619] + xnor_result[1][620] + xnor_result[1][621] + xnor_result[1][622] + xnor_result[1][623] + xnor_result[1][624] + xnor_result[1][625] + xnor_result[1][626] + xnor_result[1][627] + xnor_result[1][628] + xnor_result[1][629] + xnor_result[1][630] + xnor_result[1][631] + xnor_result[1][632] + xnor_result[1][633] + xnor_result[1][634] + xnor_result[1][635] + xnor_result[1][636] + xnor_result[1][637] + xnor_result[1][638] + xnor_result[1][639] + xnor_result[1][640] + xnor_result[1][641] + xnor_result[1][642] + xnor_result[1][643] + xnor_result[1][644] + xnor_result[1][645] + xnor_result[1][646] + xnor_result[1][647] + xnor_result[1][648] + xnor_result[1][649] + xnor_result[1][650] + xnor_result[1][651] + xnor_result[1][652] + xnor_result[1][653] + xnor_result[1][654] + xnor_result[1][655] + xnor_result[1][656] + xnor_result[1][657] + xnor_result[1][658] + xnor_result[1][659] + xnor_result[1][660] + xnor_result[1][661] + xnor_result[1][662] + xnor_result[1][663] + xnor_result[1][664] + xnor_result[1][665] + xnor_result[1][666] + xnor_result[1][667] + xnor_result[1][668] + xnor_result[1][669] + xnor_result[1][670] + xnor_result[1][671] + xnor_result[1][672] + xnor_result[1][673] + xnor_result[1][674] + xnor_result[1][675] + xnor_result[1][676] + xnor_result[1][677] + xnor_result[1][678] + xnor_result[1][679] + xnor_result[1][680] + xnor_result[1][681] + xnor_result[1][682] + xnor_result[1][683] + xnor_result[1][684] + xnor_result[1][685] + xnor_result[1][686] + xnor_result[1][687] + xnor_result[1][688] + xnor_result[1][689] + xnor_result[1][690] + xnor_result[1][691] + xnor_result[1][692] + xnor_result[1][693] + xnor_result[1][694] + xnor_result[1][695] + xnor_result[1][696] + xnor_result[1][697] + xnor_result[1][698] + xnor_result[1][699] + xnor_result[1][700] + xnor_result[1][701] + xnor_result[1][702] + xnor_result[1][703] + xnor_result[1][704] + xnor_result[1][705] + xnor_result[1][706] + xnor_result[1][707] + xnor_result[1][708] + xnor_result[1][709] + xnor_result[1][710] + xnor_result[1][711] + xnor_result[1][712] + xnor_result[1][713] + xnor_result[1][714] + xnor_result[1][715] + xnor_result[1][716] + xnor_result[1][717] + xnor_result[1][718] + xnor_result[1][719] + xnor_result[1][720] + xnor_result[1][721] + xnor_result[1][722] + xnor_result[1][723] + xnor_result[1][724] + xnor_result[1][725] + xnor_result[1][726] + xnor_result[1][727] + xnor_result[1][728] + xnor_result[1][729] + xnor_result[1][730] + xnor_result[1][731] + xnor_result[1][732] + xnor_result[1][733] + xnor_result[1][734] + xnor_result[1][735] + xnor_result[1][736] + xnor_result[1][737] + xnor_result[1][738] + xnor_result[1][739] + xnor_result[1][740] + xnor_result[1][741] + xnor_result[1][742] + xnor_result[1][743] + xnor_result[1][744] + xnor_result[1][745] + xnor_result[1][746] + xnor_result[1][747] + xnor_result[1][748] + xnor_result[1][749] + xnor_result[1][750] + xnor_result[1][751] + xnor_result[1][752] + xnor_result[1][753] + xnor_result[1][754] + xnor_result[1][755] + xnor_result[1][756] + xnor_result[1][757] + xnor_result[1][758] + xnor_result[1][759] + xnor_result[1][760] + xnor_result[1][761] + xnor_result[1][762] + xnor_result[1][763] + xnor_result[1][764] + xnor_result[1][765] + xnor_result[1][766] + xnor_result[1][767] + xnor_result[1][768] + xnor_result[1][769] + xnor_result[1][770] + xnor_result[1][771] + xnor_result[1][772] + xnor_result[1][773] + xnor_result[1][774] + xnor_result[1][775] + xnor_result[1][776] + xnor_result[1][777] + xnor_result[1][778] + xnor_result[1][779] + xnor_result[1][780] + xnor_result[1][781] + xnor_result[1][782] + xnor_result[1][783] + xnor_result[1][784] + xnor_result[1][785] + xnor_result[1][786] + xnor_result[1][787] + xnor_result[1][788] + xnor_result[1][789] + xnor_result[1][790] + xnor_result[1][791] + xnor_result[1][792] + xnor_result[1][793] + xnor_result[1][794] + xnor_result[1][795] + xnor_result[1][796] + xnor_result[1][797] + xnor_result[1][798] + xnor_result[1][799] + xnor_result[1][800] + xnor_result[1][801] + xnor_result[1][802] + xnor_result[1][803] + xnor_result[1][804] + xnor_result[1][805] + xnor_result[1][806] + xnor_result[1][807] + xnor_result[1][808] + xnor_result[1][809] + xnor_result[1][810] + xnor_result[1][811] + xnor_result[1][812] + xnor_result[1][813] + xnor_result[1][814] + xnor_result[1][815] + xnor_result[1][816] + xnor_result[1][817] + xnor_result[1][818] + xnor_result[1][819] + xnor_result[1][820] + xnor_result[1][821] + xnor_result[1][822] + xnor_result[1][823] + xnor_result[1][824] + xnor_result[1][825] + xnor_result[1][826] + xnor_result[1][827] + xnor_result[1][828] + xnor_result[1][829] + xnor_result[1][830] + xnor_result[1][831] + xnor_result[1][832] + xnor_result[1][833] + xnor_result[1][834] + xnor_result[1][835] + xnor_result[1][836] + xnor_result[1][837] + xnor_result[1][838] + xnor_result[1][839] + xnor_result[1][840] + xnor_result[1][841] + xnor_result[1][842] + xnor_result[1][843] + xnor_result[1][844] + xnor_result[1][845] + xnor_result[1][846] + xnor_result[1][847] + xnor_result[1][848] + xnor_result[1][849] + xnor_result[1][850] + xnor_result[1][851] + xnor_result[1][852] + xnor_result[1][853] + xnor_result[1][854] + xnor_result[1][855] + xnor_result[1][856] + xnor_result[1][857] + xnor_result[1][858] + xnor_result[1][859] + xnor_result[1][860] + xnor_result[1][861] + xnor_result[1][862] + xnor_result[1][863] + xnor_result[1][864] + xnor_result[1][865] + xnor_result[1][866] + xnor_result[1][867] + xnor_result[1][868] + xnor_result[1][869] + xnor_result[1][870] + xnor_result[1][871] + xnor_result[1][872] + xnor_result[1][873] + xnor_result[1][874] + xnor_result[1][875] + xnor_result[1][876] + xnor_result[1][877] + xnor_result[1][878] + xnor_result[1][879] + xnor_result[1][880] + xnor_result[1][881] + xnor_result[1][882] + xnor_result[1][883] + xnor_result[1][884] + xnor_result[1][885] + xnor_result[1][886] + xnor_result[1][887] + xnor_result[1][888] + xnor_result[1][889] + xnor_result[1][890] + xnor_result[1][891] + xnor_result[1][892] + xnor_result[1][893] + xnor_result[1][894] + xnor_result[1][895] + xnor_result[1][896] + xnor_result[1][897] + xnor_result[1][898] + xnor_result[1][899] + xnor_result[1][900] + xnor_result[1][901] + xnor_result[1][902] + xnor_result[1][903] + xnor_result[1][904] + xnor_result[1][905] + xnor_result[1][906] + xnor_result[1][907] + xnor_result[1][908] + xnor_result[1][909] + xnor_result[1][910] + xnor_result[1][911] + xnor_result[1][912] + xnor_result[1][913] + xnor_result[1][914] + xnor_result[1][915] + xnor_result[1][916] + xnor_result[1][917] + xnor_result[1][918] + xnor_result[1][919] + xnor_result[1][920] + xnor_result[1][921] + xnor_result[1][922] + xnor_result[1][923] + xnor_result[1][924] + xnor_result[1][925] + xnor_result[1][926] + xnor_result[1][927] + xnor_result[1][928] + xnor_result[1][929] + xnor_result[1][930] + xnor_result[1][931] + xnor_result[1][932] + xnor_result[1][933] + xnor_result[1][934] + xnor_result[1][935] + xnor_result[1][936] + xnor_result[1][937] + xnor_result[1][938] + xnor_result[1][939] + xnor_result[1][940] + xnor_result[1][941] + xnor_result[1][942] + xnor_result[1][943] + xnor_result[1][944] + xnor_result[1][945] + xnor_result[1][946] + xnor_result[1][947] + xnor_result[1][948] + xnor_result[1][949] + xnor_result[1][950] + xnor_result[1][951] + xnor_result[1][952] + xnor_result[1][953] + xnor_result[1][954] + xnor_result[1][955] + xnor_result[1][956] + xnor_result[1][957] + xnor_result[1][958] + xnor_result[1][959] ;
assign accumulation_result[2] = xnor_result[2][0] + xnor_result[2][1] + xnor_result[2][2] + xnor_result[2][3] + xnor_result[2][4] + xnor_result[2][5] + xnor_result[2][6] + xnor_result[2][7] + xnor_result[2][8] + xnor_result[2][9] + xnor_result[2][10] + xnor_result[2][11] + xnor_result[2][12] + xnor_result[2][13] + xnor_result[2][14] + xnor_result[2][15] + xnor_result[2][16] + xnor_result[2][17] + xnor_result[2][18] + xnor_result[2][19] + xnor_result[2][20] + xnor_result[2][21] + xnor_result[2][22] + xnor_result[2][23] + xnor_result[2][24] + xnor_result[2][25] + xnor_result[2][26] + xnor_result[2][27] + xnor_result[2][28] + xnor_result[2][29] + xnor_result[2][30] + xnor_result[2][31] + xnor_result[2][32] + xnor_result[2][33] + xnor_result[2][34] + xnor_result[2][35] + xnor_result[2][36] + xnor_result[2][37] + xnor_result[2][38] + xnor_result[2][39] + xnor_result[2][40] + xnor_result[2][41] + xnor_result[2][42] + xnor_result[2][43] + xnor_result[2][44] + xnor_result[2][45] + xnor_result[2][46] + xnor_result[2][47] + xnor_result[2][48] + xnor_result[2][49] + xnor_result[2][50] + xnor_result[2][51] + xnor_result[2][52] + xnor_result[2][53] + xnor_result[2][54] + xnor_result[2][55] + xnor_result[2][56] + xnor_result[2][57] + xnor_result[2][58] + xnor_result[2][59] + xnor_result[2][60] + xnor_result[2][61] + xnor_result[2][62] + xnor_result[2][63] + xnor_result[2][64] + xnor_result[2][65] + xnor_result[2][66] + xnor_result[2][67] + xnor_result[2][68] + xnor_result[2][69] + xnor_result[2][70] + xnor_result[2][71] + xnor_result[2][72] + xnor_result[2][73] + xnor_result[2][74] + xnor_result[2][75] + xnor_result[2][76] + xnor_result[2][77] + xnor_result[2][78] + xnor_result[2][79] + xnor_result[2][80] + xnor_result[2][81] + xnor_result[2][82] + xnor_result[2][83] + xnor_result[2][84] + xnor_result[2][85] + xnor_result[2][86] + xnor_result[2][87] + xnor_result[2][88] + xnor_result[2][89] + xnor_result[2][90] + xnor_result[2][91] + xnor_result[2][92] + xnor_result[2][93] + xnor_result[2][94] + xnor_result[2][95] + xnor_result[2][96] + xnor_result[2][97] + xnor_result[2][98] + xnor_result[2][99] + xnor_result[2][100] + xnor_result[2][101] + xnor_result[2][102] + xnor_result[2][103] + xnor_result[2][104] + xnor_result[2][105] + xnor_result[2][106] + xnor_result[2][107] + xnor_result[2][108] + xnor_result[2][109] + xnor_result[2][110] + xnor_result[2][111] + xnor_result[2][112] + xnor_result[2][113] + xnor_result[2][114] + xnor_result[2][115] + xnor_result[2][116] + xnor_result[2][117] + xnor_result[2][118] + xnor_result[2][119] + xnor_result[2][120] + xnor_result[2][121] + xnor_result[2][122] + xnor_result[2][123] + xnor_result[2][124] + xnor_result[2][125] + xnor_result[2][126] + xnor_result[2][127] + xnor_result[2][128] + xnor_result[2][129] + xnor_result[2][130] + xnor_result[2][131] + xnor_result[2][132] + xnor_result[2][133] + xnor_result[2][134] + xnor_result[2][135] + xnor_result[2][136] + xnor_result[2][137] + xnor_result[2][138] + xnor_result[2][139] + xnor_result[2][140] + xnor_result[2][141] + xnor_result[2][142] + xnor_result[2][143] + xnor_result[2][144] + xnor_result[2][145] + xnor_result[2][146] + xnor_result[2][147] + xnor_result[2][148] + xnor_result[2][149] + xnor_result[2][150] + xnor_result[2][151] + xnor_result[2][152] + xnor_result[2][153] + xnor_result[2][154] + xnor_result[2][155] + xnor_result[2][156] + xnor_result[2][157] + xnor_result[2][158] + xnor_result[2][159] + xnor_result[2][160] + xnor_result[2][161] + xnor_result[2][162] + xnor_result[2][163] + xnor_result[2][164] + xnor_result[2][165] + xnor_result[2][166] + xnor_result[2][167] + xnor_result[2][168] + xnor_result[2][169] + xnor_result[2][170] + xnor_result[2][171] + xnor_result[2][172] + xnor_result[2][173] + xnor_result[2][174] + xnor_result[2][175] + xnor_result[2][176] + xnor_result[2][177] + xnor_result[2][178] + xnor_result[2][179] + xnor_result[2][180] + xnor_result[2][181] + xnor_result[2][182] + xnor_result[2][183] + xnor_result[2][184] + xnor_result[2][185] + xnor_result[2][186] + xnor_result[2][187] + xnor_result[2][188] + xnor_result[2][189] + xnor_result[2][190] + xnor_result[2][191] + xnor_result[2][192] + xnor_result[2][193] + xnor_result[2][194] + xnor_result[2][195] + xnor_result[2][196] + xnor_result[2][197] + xnor_result[2][198] + xnor_result[2][199] + xnor_result[2][200] + xnor_result[2][201] + xnor_result[2][202] + xnor_result[2][203] + xnor_result[2][204] + xnor_result[2][205] + xnor_result[2][206] + xnor_result[2][207] + xnor_result[2][208] + xnor_result[2][209] + xnor_result[2][210] + xnor_result[2][211] + xnor_result[2][212] + xnor_result[2][213] + xnor_result[2][214] + xnor_result[2][215] + xnor_result[2][216] + xnor_result[2][217] + xnor_result[2][218] + xnor_result[2][219] + xnor_result[2][220] + xnor_result[2][221] + xnor_result[2][222] + xnor_result[2][223] + xnor_result[2][224] + xnor_result[2][225] + xnor_result[2][226] + xnor_result[2][227] + xnor_result[2][228] + xnor_result[2][229] + xnor_result[2][230] + xnor_result[2][231] + xnor_result[2][232] + xnor_result[2][233] + xnor_result[2][234] + xnor_result[2][235] + xnor_result[2][236] + xnor_result[2][237] + xnor_result[2][238] + xnor_result[2][239] + xnor_result[2][240] + xnor_result[2][241] + xnor_result[2][242] + xnor_result[2][243] + xnor_result[2][244] + xnor_result[2][245] + xnor_result[2][246] + xnor_result[2][247] + xnor_result[2][248] + xnor_result[2][249] + xnor_result[2][250] + xnor_result[2][251] + xnor_result[2][252] + xnor_result[2][253] + xnor_result[2][254] + xnor_result[2][255] + xnor_result[2][256] + xnor_result[2][257] + xnor_result[2][258] + xnor_result[2][259] + xnor_result[2][260] + xnor_result[2][261] + xnor_result[2][262] + xnor_result[2][263] + xnor_result[2][264] + xnor_result[2][265] + xnor_result[2][266] + xnor_result[2][267] + xnor_result[2][268] + xnor_result[2][269] + xnor_result[2][270] + xnor_result[2][271] + xnor_result[2][272] + xnor_result[2][273] + xnor_result[2][274] + xnor_result[2][275] + xnor_result[2][276] + xnor_result[2][277] + xnor_result[2][278] + xnor_result[2][279] + xnor_result[2][280] + xnor_result[2][281] + xnor_result[2][282] + xnor_result[2][283] + xnor_result[2][284] + xnor_result[2][285] + xnor_result[2][286] + xnor_result[2][287] + xnor_result[2][288] + xnor_result[2][289] + xnor_result[2][290] + xnor_result[2][291] + xnor_result[2][292] + xnor_result[2][293] + xnor_result[2][294] + xnor_result[2][295] + xnor_result[2][296] + xnor_result[2][297] + xnor_result[2][298] + xnor_result[2][299] + xnor_result[2][300] + xnor_result[2][301] + xnor_result[2][302] + xnor_result[2][303] + xnor_result[2][304] + xnor_result[2][305] + xnor_result[2][306] + xnor_result[2][307] + xnor_result[2][308] + xnor_result[2][309] + xnor_result[2][310] + xnor_result[2][311] + xnor_result[2][312] + xnor_result[2][313] + xnor_result[2][314] + xnor_result[2][315] + xnor_result[2][316] + xnor_result[2][317] + xnor_result[2][318] + xnor_result[2][319] + xnor_result[2][320] + xnor_result[2][321] + xnor_result[2][322] + xnor_result[2][323] + xnor_result[2][324] + xnor_result[2][325] + xnor_result[2][326] + xnor_result[2][327] + xnor_result[2][328] + xnor_result[2][329] + xnor_result[2][330] + xnor_result[2][331] + xnor_result[2][332] + xnor_result[2][333] + xnor_result[2][334] + xnor_result[2][335] + xnor_result[2][336] + xnor_result[2][337] + xnor_result[2][338] + xnor_result[2][339] + xnor_result[2][340] + xnor_result[2][341] + xnor_result[2][342] + xnor_result[2][343] + xnor_result[2][344] + xnor_result[2][345] + xnor_result[2][346] + xnor_result[2][347] + xnor_result[2][348] + xnor_result[2][349] + xnor_result[2][350] + xnor_result[2][351] + xnor_result[2][352] + xnor_result[2][353] + xnor_result[2][354] + xnor_result[2][355] + xnor_result[2][356] + xnor_result[2][357] + xnor_result[2][358] + xnor_result[2][359] + xnor_result[2][360] + xnor_result[2][361] + xnor_result[2][362] + xnor_result[2][363] + xnor_result[2][364] + xnor_result[2][365] + xnor_result[2][366] + xnor_result[2][367] + xnor_result[2][368] + xnor_result[2][369] + xnor_result[2][370] + xnor_result[2][371] + xnor_result[2][372] + xnor_result[2][373] + xnor_result[2][374] + xnor_result[2][375] + xnor_result[2][376] + xnor_result[2][377] + xnor_result[2][378] + xnor_result[2][379] + xnor_result[2][380] + xnor_result[2][381] + xnor_result[2][382] + xnor_result[2][383] + xnor_result[2][384] + xnor_result[2][385] + xnor_result[2][386] + xnor_result[2][387] + xnor_result[2][388] + xnor_result[2][389] + xnor_result[2][390] + xnor_result[2][391] + xnor_result[2][392] + xnor_result[2][393] + xnor_result[2][394] + xnor_result[2][395] + xnor_result[2][396] + xnor_result[2][397] + xnor_result[2][398] + xnor_result[2][399] + xnor_result[2][400] + xnor_result[2][401] + xnor_result[2][402] + xnor_result[2][403] + xnor_result[2][404] + xnor_result[2][405] + xnor_result[2][406] + xnor_result[2][407] + xnor_result[2][408] + xnor_result[2][409] + xnor_result[2][410] + xnor_result[2][411] + xnor_result[2][412] + xnor_result[2][413] + xnor_result[2][414] + xnor_result[2][415] + xnor_result[2][416] + xnor_result[2][417] + xnor_result[2][418] + xnor_result[2][419] + xnor_result[2][420] + xnor_result[2][421] + xnor_result[2][422] + xnor_result[2][423] + xnor_result[2][424] + xnor_result[2][425] + xnor_result[2][426] + xnor_result[2][427] + xnor_result[2][428] + xnor_result[2][429] + xnor_result[2][430] + xnor_result[2][431] + xnor_result[2][432] + xnor_result[2][433] + xnor_result[2][434] + xnor_result[2][435] + xnor_result[2][436] + xnor_result[2][437] + xnor_result[2][438] + xnor_result[2][439] + xnor_result[2][440] + xnor_result[2][441] + xnor_result[2][442] + xnor_result[2][443] + xnor_result[2][444] + xnor_result[2][445] + xnor_result[2][446] + xnor_result[2][447] + xnor_result[2][448] + xnor_result[2][449] + xnor_result[2][450] + xnor_result[2][451] + xnor_result[2][452] + xnor_result[2][453] + xnor_result[2][454] + xnor_result[2][455] + xnor_result[2][456] + xnor_result[2][457] + xnor_result[2][458] + xnor_result[2][459] + xnor_result[2][460] + xnor_result[2][461] + xnor_result[2][462] + xnor_result[2][463] + xnor_result[2][464] + xnor_result[2][465] + xnor_result[2][466] + xnor_result[2][467] + xnor_result[2][468] + xnor_result[2][469] + xnor_result[2][470] + xnor_result[2][471] + xnor_result[2][472] + xnor_result[2][473] + xnor_result[2][474] + xnor_result[2][475] + xnor_result[2][476] + xnor_result[2][477] + xnor_result[2][478] + xnor_result[2][479] + xnor_result[2][480] + xnor_result[2][481] + xnor_result[2][482] + xnor_result[2][483] + xnor_result[2][484] + xnor_result[2][485] + xnor_result[2][486] + xnor_result[2][487] + xnor_result[2][488] + xnor_result[2][489] + xnor_result[2][490] + xnor_result[2][491] + xnor_result[2][492] + xnor_result[2][493] + xnor_result[2][494] + xnor_result[2][495] + xnor_result[2][496] + xnor_result[2][497] + xnor_result[2][498] + xnor_result[2][499] + xnor_result[2][500] + xnor_result[2][501] + xnor_result[2][502] + xnor_result[2][503] + xnor_result[2][504] + xnor_result[2][505] + xnor_result[2][506] + xnor_result[2][507] + xnor_result[2][508] + xnor_result[2][509] + xnor_result[2][510] + xnor_result[2][511] + xnor_result[2][512] + xnor_result[2][513] + xnor_result[2][514] + xnor_result[2][515] + xnor_result[2][516] + xnor_result[2][517] + xnor_result[2][518] + xnor_result[2][519] + xnor_result[2][520] + xnor_result[2][521] + xnor_result[2][522] + xnor_result[2][523] + xnor_result[2][524] + xnor_result[2][525] + xnor_result[2][526] + xnor_result[2][527] + xnor_result[2][528] + xnor_result[2][529] + xnor_result[2][530] + xnor_result[2][531] + xnor_result[2][532] + xnor_result[2][533] + xnor_result[2][534] + xnor_result[2][535] + xnor_result[2][536] + xnor_result[2][537] + xnor_result[2][538] + xnor_result[2][539] + xnor_result[2][540] + xnor_result[2][541] + xnor_result[2][542] + xnor_result[2][543] + xnor_result[2][544] + xnor_result[2][545] + xnor_result[2][546] + xnor_result[2][547] + xnor_result[2][548] + xnor_result[2][549] + xnor_result[2][550] + xnor_result[2][551] + xnor_result[2][552] + xnor_result[2][553] + xnor_result[2][554] + xnor_result[2][555] + xnor_result[2][556] + xnor_result[2][557] + xnor_result[2][558] + xnor_result[2][559] + xnor_result[2][560] + xnor_result[2][561] + xnor_result[2][562] + xnor_result[2][563] + xnor_result[2][564] + xnor_result[2][565] + xnor_result[2][566] + xnor_result[2][567] + xnor_result[2][568] + xnor_result[2][569] + xnor_result[2][570] + xnor_result[2][571] + xnor_result[2][572] + xnor_result[2][573] + xnor_result[2][574] + xnor_result[2][575] + xnor_result[2][576] + xnor_result[2][577] + xnor_result[2][578] + xnor_result[2][579] + xnor_result[2][580] + xnor_result[2][581] + xnor_result[2][582] + xnor_result[2][583] + xnor_result[2][584] + xnor_result[2][585] + xnor_result[2][586] + xnor_result[2][587] + xnor_result[2][588] + xnor_result[2][589] + xnor_result[2][590] + xnor_result[2][591] + xnor_result[2][592] + xnor_result[2][593] + xnor_result[2][594] + xnor_result[2][595] + xnor_result[2][596] + xnor_result[2][597] + xnor_result[2][598] + xnor_result[2][599] + xnor_result[2][600] + xnor_result[2][601] + xnor_result[2][602] + xnor_result[2][603] + xnor_result[2][604] + xnor_result[2][605] + xnor_result[2][606] + xnor_result[2][607] + xnor_result[2][608] + xnor_result[2][609] + xnor_result[2][610] + xnor_result[2][611] + xnor_result[2][612] + xnor_result[2][613] + xnor_result[2][614] + xnor_result[2][615] + xnor_result[2][616] + xnor_result[2][617] + xnor_result[2][618] + xnor_result[2][619] + xnor_result[2][620] + xnor_result[2][621] + xnor_result[2][622] + xnor_result[2][623] + xnor_result[2][624] + xnor_result[2][625] + xnor_result[2][626] + xnor_result[2][627] + xnor_result[2][628] + xnor_result[2][629] + xnor_result[2][630] + xnor_result[2][631] + xnor_result[2][632] + xnor_result[2][633] + xnor_result[2][634] + xnor_result[2][635] + xnor_result[2][636] + xnor_result[2][637] + xnor_result[2][638] + xnor_result[2][639] + xnor_result[2][640] + xnor_result[2][641] + xnor_result[2][642] + xnor_result[2][643] + xnor_result[2][644] + xnor_result[2][645] + xnor_result[2][646] + xnor_result[2][647] + xnor_result[2][648] + xnor_result[2][649] + xnor_result[2][650] + xnor_result[2][651] + xnor_result[2][652] + xnor_result[2][653] + xnor_result[2][654] + xnor_result[2][655] + xnor_result[2][656] + xnor_result[2][657] + xnor_result[2][658] + xnor_result[2][659] + xnor_result[2][660] + xnor_result[2][661] + xnor_result[2][662] + xnor_result[2][663] + xnor_result[2][664] + xnor_result[2][665] + xnor_result[2][666] + xnor_result[2][667] + xnor_result[2][668] + xnor_result[2][669] + xnor_result[2][670] + xnor_result[2][671] + xnor_result[2][672] + xnor_result[2][673] + xnor_result[2][674] + xnor_result[2][675] + xnor_result[2][676] + xnor_result[2][677] + xnor_result[2][678] + xnor_result[2][679] + xnor_result[2][680] + xnor_result[2][681] + xnor_result[2][682] + xnor_result[2][683] + xnor_result[2][684] + xnor_result[2][685] + xnor_result[2][686] + xnor_result[2][687] + xnor_result[2][688] + xnor_result[2][689] + xnor_result[2][690] + xnor_result[2][691] + xnor_result[2][692] + xnor_result[2][693] + xnor_result[2][694] + xnor_result[2][695] + xnor_result[2][696] + xnor_result[2][697] + xnor_result[2][698] + xnor_result[2][699] + xnor_result[2][700] + xnor_result[2][701] + xnor_result[2][702] + xnor_result[2][703] + xnor_result[2][704] + xnor_result[2][705] + xnor_result[2][706] + xnor_result[2][707] + xnor_result[2][708] + xnor_result[2][709] + xnor_result[2][710] + xnor_result[2][711] + xnor_result[2][712] + xnor_result[2][713] + xnor_result[2][714] + xnor_result[2][715] + xnor_result[2][716] + xnor_result[2][717] + xnor_result[2][718] + xnor_result[2][719] + xnor_result[2][720] + xnor_result[2][721] + xnor_result[2][722] + xnor_result[2][723] + xnor_result[2][724] + xnor_result[2][725] + xnor_result[2][726] + xnor_result[2][727] + xnor_result[2][728] + xnor_result[2][729] + xnor_result[2][730] + xnor_result[2][731] + xnor_result[2][732] + xnor_result[2][733] + xnor_result[2][734] + xnor_result[2][735] + xnor_result[2][736] + xnor_result[2][737] + xnor_result[2][738] + xnor_result[2][739] + xnor_result[2][740] + xnor_result[2][741] + xnor_result[2][742] + xnor_result[2][743] + xnor_result[2][744] + xnor_result[2][745] + xnor_result[2][746] + xnor_result[2][747] + xnor_result[2][748] + xnor_result[2][749] + xnor_result[2][750] + xnor_result[2][751] + xnor_result[2][752] + xnor_result[2][753] + xnor_result[2][754] + xnor_result[2][755] + xnor_result[2][756] + xnor_result[2][757] + xnor_result[2][758] + xnor_result[2][759] + xnor_result[2][760] + xnor_result[2][761] + xnor_result[2][762] + xnor_result[2][763] + xnor_result[2][764] + xnor_result[2][765] + xnor_result[2][766] + xnor_result[2][767] + xnor_result[2][768] + xnor_result[2][769] + xnor_result[2][770] + xnor_result[2][771] + xnor_result[2][772] + xnor_result[2][773] + xnor_result[2][774] + xnor_result[2][775] + xnor_result[2][776] + xnor_result[2][777] + xnor_result[2][778] + xnor_result[2][779] + xnor_result[2][780] + xnor_result[2][781] + xnor_result[2][782] + xnor_result[2][783] + xnor_result[2][784] + xnor_result[2][785] + xnor_result[2][786] + xnor_result[2][787] + xnor_result[2][788] + xnor_result[2][789] + xnor_result[2][790] + xnor_result[2][791] + xnor_result[2][792] + xnor_result[2][793] + xnor_result[2][794] + xnor_result[2][795] + xnor_result[2][796] + xnor_result[2][797] + xnor_result[2][798] + xnor_result[2][799] + xnor_result[2][800] + xnor_result[2][801] + xnor_result[2][802] + xnor_result[2][803] + xnor_result[2][804] + xnor_result[2][805] + xnor_result[2][806] + xnor_result[2][807] + xnor_result[2][808] + xnor_result[2][809] + xnor_result[2][810] + xnor_result[2][811] + xnor_result[2][812] + xnor_result[2][813] + xnor_result[2][814] + xnor_result[2][815] + xnor_result[2][816] + xnor_result[2][817] + xnor_result[2][818] + xnor_result[2][819] + xnor_result[2][820] + xnor_result[2][821] + xnor_result[2][822] + xnor_result[2][823] + xnor_result[2][824] + xnor_result[2][825] + xnor_result[2][826] + xnor_result[2][827] + xnor_result[2][828] + xnor_result[2][829] + xnor_result[2][830] + xnor_result[2][831] + xnor_result[2][832] + xnor_result[2][833] + xnor_result[2][834] + xnor_result[2][835] + xnor_result[2][836] + xnor_result[2][837] + xnor_result[2][838] + xnor_result[2][839] + xnor_result[2][840] + xnor_result[2][841] + xnor_result[2][842] + xnor_result[2][843] + xnor_result[2][844] + xnor_result[2][845] + xnor_result[2][846] + xnor_result[2][847] + xnor_result[2][848] + xnor_result[2][849] + xnor_result[2][850] + xnor_result[2][851] + xnor_result[2][852] + xnor_result[2][853] + xnor_result[2][854] + xnor_result[2][855] + xnor_result[2][856] + xnor_result[2][857] + xnor_result[2][858] + xnor_result[2][859] + xnor_result[2][860] + xnor_result[2][861] + xnor_result[2][862] + xnor_result[2][863] + xnor_result[2][864] + xnor_result[2][865] + xnor_result[2][866] + xnor_result[2][867] + xnor_result[2][868] + xnor_result[2][869] + xnor_result[2][870] + xnor_result[2][871] + xnor_result[2][872] + xnor_result[2][873] + xnor_result[2][874] + xnor_result[2][875] + xnor_result[2][876] + xnor_result[2][877] + xnor_result[2][878] + xnor_result[2][879] + xnor_result[2][880] + xnor_result[2][881] + xnor_result[2][882] + xnor_result[2][883] + xnor_result[2][884] + xnor_result[2][885] + xnor_result[2][886] + xnor_result[2][887] + xnor_result[2][888] + xnor_result[2][889] + xnor_result[2][890] + xnor_result[2][891] + xnor_result[2][892] + xnor_result[2][893] + xnor_result[2][894] + xnor_result[2][895] + xnor_result[2][896] + xnor_result[2][897] + xnor_result[2][898] + xnor_result[2][899] + xnor_result[2][900] + xnor_result[2][901] + xnor_result[2][902] + xnor_result[2][903] + xnor_result[2][904] + xnor_result[2][905] + xnor_result[2][906] + xnor_result[2][907] + xnor_result[2][908] + xnor_result[2][909] + xnor_result[2][910] + xnor_result[2][911] + xnor_result[2][912] + xnor_result[2][913] + xnor_result[2][914] + xnor_result[2][915] + xnor_result[2][916] + xnor_result[2][917] + xnor_result[2][918] + xnor_result[2][919] + xnor_result[2][920] + xnor_result[2][921] + xnor_result[2][922] + xnor_result[2][923] + xnor_result[2][924] + xnor_result[2][925] + xnor_result[2][926] + xnor_result[2][927] + xnor_result[2][928] + xnor_result[2][929] + xnor_result[2][930] + xnor_result[2][931] + xnor_result[2][932] + xnor_result[2][933] + xnor_result[2][934] + xnor_result[2][935] + xnor_result[2][936] + xnor_result[2][937] + xnor_result[2][938] + xnor_result[2][939] + xnor_result[2][940] + xnor_result[2][941] + xnor_result[2][942] + xnor_result[2][943] + xnor_result[2][944] + xnor_result[2][945] + xnor_result[2][946] + xnor_result[2][947] + xnor_result[2][948] + xnor_result[2][949] + xnor_result[2][950] + xnor_result[2][951] + xnor_result[2][952] + xnor_result[2][953] + xnor_result[2][954] + xnor_result[2][955] + xnor_result[2][956] + xnor_result[2][957] + xnor_result[2][958] + xnor_result[2][959] ;
assign accumulation_result[3] = xnor_result[3][0] + xnor_result[3][1] + xnor_result[3][2] + xnor_result[3][3] + xnor_result[3][4] + xnor_result[3][5] + xnor_result[3][6] + xnor_result[3][7] + xnor_result[3][8] + xnor_result[3][9] + xnor_result[3][10] + xnor_result[3][11] + xnor_result[3][12] + xnor_result[3][13] + xnor_result[3][14] + xnor_result[3][15] + xnor_result[3][16] + xnor_result[3][17] + xnor_result[3][18] + xnor_result[3][19] + xnor_result[3][20] + xnor_result[3][21] + xnor_result[3][22] + xnor_result[3][23] + xnor_result[3][24] + xnor_result[3][25] + xnor_result[3][26] + xnor_result[3][27] + xnor_result[3][28] + xnor_result[3][29] + xnor_result[3][30] + xnor_result[3][31] + xnor_result[3][32] + xnor_result[3][33] + xnor_result[3][34] + xnor_result[3][35] + xnor_result[3][36] + xnor_result[3][37] + xnor_result[3][38] + xnor_result[3][39] + xnor_result[3][40] + xnor_result[3][41] + xnor_result[3][42] + xnor_result[3][43] + xnor_result[3][44] + xnor_result[3][45] + xnor_result[3][46] + xnor_result[3][47] + xnor_result[3][48] + xnor_result[3][49] + xnor_result[3][50] + xnor_result[3][51] + xnor_result[3][52] + xnor_result[3][53] + xnor_result[3][54] + xnor_result[3][55] + xnor_result[3][56] + xnor_result[3][57] + xnor_result[3][58] + xnor_result[3][59] + xnor_result[3][60] + xnor_result[3][61] + xnor_result[3][62] + xnor_result[3][63] + xnor_result[3][64] + xnor_result[3][65] + xnor_result[3][66] + xnor_result[3][67] + xnor_result[3][68] + xnor_result[3][69] + xnor_result[3][70] + xnor_result[3][71] + xnor_result[3][72] + xnor_result[3][73] + xnor_result[3][74] + xnor_result[3][75] + xnor_result[3][76] + xnor_result[3][77] + xnor_result[3][78] + xnor_result[3][79] + xnor_result[3][80] + xnor_result[3][81] + xnor_result[3][82] + xnor_result[3][83] + xnor_result[3][84] + xnor_result[3][85] + xnor_result[3][86] + xnor_result[3][87] + xnor_result[3][88] + xnor_result[3][89] + xnor_result[3][90] + xnor_result[3][91] + xnor_result[3][92] + xnor_result[3][93] + xnor_result[3][94] + xnor_result[3][95] + xnor_result[3][96] + xnor_result[3][97] + xnor_result[3][98] + xnor_result[3][99] + xnor_result[3][100] + xnor_result[3][101] + xnor_result[3][102] + xnor_result[3][103] + xnor_result[3][104] + xnor_result[3][105] + xnor_result[3][106] + xnor_result[3][107] + xnor_result[3][108] + xnor_result[3][109] + xnor_result[3][110] + xnor_result[3][111] + xnor_result[3][112] + xnor_result[3][113] + xnor_result[3][114] + xnor_result[3][115] + xnor_result[3][116] + xnor_result[3][117] + xnor_result[3][118] + xnor_result[3][119] + xnor_result[3][120] + xnor_result[3][121] + xnor_result[3][122] + xnor_result[3][123] + xnor_result[3][124] + xnor_result[3][125] + xnor_result[3][126] + xnor_result[3][127] + xnor_result[3][128] + xnor_result[3][129] + xnor_result[3][130] + xnor_result[3][131] + xnor_result[3][132] + xnor_result[3][133] + xnor_result[3][134] + xnor_result[3][135] + xnor_result[3][136] + xnor_result[3][137] + xnor_result[3][138] + xnor_result[3][139] + xnor_result[3][140] + xnor_result[3][141] + xnor_result[3][142] + xnor_result[3][143] + xnor_result[3][144] + xnor_result[3][145] + xnor_result[3][146] + xnor_result[3][147] + xnor_result[3][148] + xnor_result[3][149] + xnor_result[3][150] + xnor_result[3][151] + xnor_result[3][152] + xnor_result[3][153] + xnor_result[3][154] + xnor_result[3][155] + xnor_result[3][156] + xnor_result[3][157] + xnor_result[3][158] + xnor_result[3][159] + xnor_result[3][160] + xnor_result[3][161] + xnor_result[3][162] + xnor_result[3][163] + xnor_result[3][164] + xnor_result[3][165] + xnor_result[3][166] + xnor_result[3][167] + xnor_result[3][168] + xnor_result[3][169] + xnor_result[3][170] + xnor_result[3][171] + xnor_result[3][172] + xnor_result[3][173] + xnor_result[3][174] + xnor_result[3][175] + xnor_result[3][176] + xnor_result[3][177] + xnor_result[3][178] + xnor_result[3][179] + xnor_result[3][180] + xnor_result[3][181] + xnor_result[3][182] + xnor_result[3][183] + xnor_result[3][184] + xnor_result[3][185] + xnor_result[3][186] + xnor_result[3][187] + xnor_result[3][188] + xnor_result[3][189] + xnor_result[3][190] + xnor_result[3][191] + xnor_result[3][192] + xnor_result[3][193] + xnor_result[3][194] + xnor_result[3][195] + xnor_result[3][196] + xnor_result[3][197] + xnor_result[3][198] + xnor_result[3][199] + xnor_result[3][200] + xnor_result[3][201] + xnor_result[3][202] + xnor_result[3][203] + xnor_result[3][204] + xnor_result[3][205] + xnor_result[3][206] + xnor_result[3][207] + xnor_result[3][208] + xnor_result[3][209] + xnor_result[3][210] + xnor_result[3][211] + xnor_result[3][212] + xnor_result[3][213] + xnor_result[3][214] + xnor_result[3][215] + xnor_result[3][216] + xnor_result[3][217] + xnor_result[3][218] + xnor_result[3][219] + xnor_result[3][220] + xnor_result[3][221] + xnor_result[3][222] + xnor_result[3][223] + xnor_result[3][224] + xnor_result[3][225] + xnor_result[3][226] + xnor_result[3][227] + xnor_result[3][228] + xnor_result[3][229] + xnor_result[3][230] + xnor_result[3][231] + xnor_result[3][232] + xnor_result[3][233] + xnor_result[3][234] + xnor_result[3][235] + xnor_result[3][236] + xnor_result[3][237] + xnor_result[3][238] + xnor_result[3][239] + xnor_result[3][240] + xnor_result[3][241] + xnor_result[3][242] + xnor_result[3][243] + xnor_result[3][244] + xnor_result[3][245] + xnor_result[3][246] + xnor_result[3][247] + xnor_result[3][248] + xnor_result[3][249] + xnor_result[3][250] + xnor_result[3][251] + xnor_result[3][252] + xnor_result[3][253] + xnor_result[3][254] + xnor_result[3][255] + xnor_result[3][256] + xnor_result[3][257] + xnor_result[3][258] + xnor_result[3][259] + xnor_result[3][260] + xnor_result[3][261] + xnor_result[3][262] + xnor_result[3][263] + xnor_result[3][264] + xnor_result[3][265] + xnor_result[3][266] + xnor_result[3][267] + xnor_result[3][268] + xnor_result[3][269] + xnor_result[3][270] + xnor_result[3][271] + xnor_result[3][272] + xnor_result[3][273] + xnor_result[3][274] + xnor_result[3][275] + xnor_result[3][276] + xnor_result[3][277] + xnor_result[3][278] + xnor_result[3][279] + xnor_result[3][280] + xnor_result[3][281] + xnor_result[3][282] + xnor_result[3][283] + xnor_result[3][284] + xnor_result[3][285] + xnor_result[3][286] + xnor_result[3][287] + xnor_result[3][288] + xnor_result[3][289] + xnor_result[3][290] + xnor_result[3][291] + xnor_result[3][292] + xnor_result[3][293] + xnor_result[3][294] + xnor_result[3][295] + xnor_result[3][296] + xnor_result[3][297] + xnor_result[3][298] + xnor_result[3][299] + xnor_result[3][300] + xnor_result[3][301] + xnor_result[3][302] + xnor_result[3][303] + xnor_result[3][304] + xnor_result[3][305] + xnor_result[3][306] + xnor_result[3][307] + xnor_result[3][308] + xnor_result[3][309] + xnor_result[3][310] + xnor_result[3][311] + xnor_result[3][312] + xnor_result[3][313] + xnor_result[3][314] + xnor_result[3][315] + xnor_result[3][316] + xnor_result[3][317] + xnor_result[3][318] + xnor_result[3][319] + xnor_result[3][320] + xnor_result[3][321] + xnor_result[3][322] + xnor_result[3][323] + xnor_result[3][324] + xnor_result[3][325] + xnor_result[3][326] + xnor_result[3][327] + xnor_result[3][328] + xnor_result[3][329] + xnor_result[3][330] + xnor_result[3][331] + xnor_result[3][332] + xnor_result[3][333] + xnor_result[3][334] + xnor_result[3][335] + xnor_result[3][336] + xnor_result[3][337] + xnor_result[3][338] + xnor_result[3][339] + xnor_result[3][340] + xnor_result[3][341] + xnor_result[3][342] + xnor_result[3][343] + xnor_result[3][344] + xnor_result[3][345] + xnor_result[3][346] + xnor_result[3][347] + xnor_result[3][348] + xnor_result[3][349] + xnor_result[3][350] + xnor_result[3][351] + xnor_result[3][352] + xnor_result[3][353] + xnor_result[3][354] + xnor_result[3][355] + xnor_result[3][356] + xnor_result[3][357] + xnor_result[3][358] + xnor_result[3][359] + xnor_result[3][360] + xnor_result[3][361] + xnor_result[3][362] + xnor_result[3][363] + xnor_result[3][364] + xnor_result[3][365] + xnor_result[3][366] + xnor_result[3][367] + xnor_result[3][368] + xnor_result[3][369] + xnor_result[3][370] + xnor_result[3][371] + xnor_result[3][372] + xnor_result[3][373] + xnor_result[3][374] + xnor_result[3][375] + xnor_result[3][376] + xnor_result[3][377] + xnor_result[3][378] + xnor_result[3][379] + xnor_result[3][380] + xnor_result[3][381] + xnor_result[3][382] + xnor_result[3][383] + xnor_result[3][384] + xnor_result[3][385] + xnor_result[3][386] + xnor_result[3][387] + xnor_result[3][388] + xnor_result[3][389] + xnor_result[3][390] + xnor_result[3][391] + xnor_result[3][392] + xnor_result[3][393] + xnor_result[3][394] + xnor_result[3][395] + xnor_result[3][396] + xnor_result[3][397] + xnor_result[3][398] + xnor_result[3][399] + xnor_result[3][400] + xnor_result[3][401] + xnor_result[3][402] + xnor_result[3][403] + xnor_result[3][404] + xnor_result[3][405] + xnor_result[3][406] + xnor_result[3][407] + xnor_result[3][408] + xnor_result[3][409] + xnor_result[3][410] + xnor_result[3][411] + xnor_result[3][412] + xnor_result[3][413] + xnor_result[3][414] + xnor_result[3][415] + xnor_result[3][416] + xnor_result[3][417] + xnor_result[3][418] + xnor_result[3][419] + xnor_result[3][420] + xnor_result[3][421] + xnor_result[3][422] + xnor_result[3][423] + xnor_result[3][424] + xnor_result[3][425] + xnor_result[3][426] + xnor_result[3][427] + xnor_result[3][428] + xnor_result[3][429] + xnor_result[3][430] + xnor_result[3][431] + xnor_result[3][432] + xnor_result[3][433] + xnor_result[3][434] + xnor_result[3][435] + xnor_result[3][436] + xnor_result[3][437] + xnor_result[3][438] + xnor_result[3][439] + xnor_result[3][440] + xnor_result[3][441] + xnor_result[3][442] + xnor_result[3][443] + xnor_result[3][444] + xnor_result[3][445] + xnor_result[3][446] + xnor_result[3][447] + xnor_result[3][448] + xnor_result[3][449] + xnor_result[3][450] + xnor_result[3][451] + xnor_result[3][452] + xnor_result[3][453] + xnor_result[3][454] + xnor_result[3][455] + xnor_result[3][456] + xnor_result[3][457] + xnor_result[3][458] + xnor_result[3][459] + xnor_result[3][460] + xnor_result[3][461] + xnor_result[3][462] + xnor_result[3][463] + xnor_result[3][464] + xnor_result[3][465] + xnor_result[3][466] + xnor_result[3][467] + xnor_result[3][468] + xnor_result[3][469] + xnor_result[3][470] + xnor_result[3][471] + xnor_result[3][472] + xnor_result[3][473] + xnor_result[3][474] + xnor_result[3][475] + xnor_result[3][476] + xnor_result[3][477] + xnor_result[3][478] + xnor_result[3][479] + xnor_result[3][480] + xnor_result[3][481] + xnor_result[3][482] + xnor_result[3][483] + xnor_result[3][484] + xnor_result[3][485] + xnor_result[3][486] + xnor_result[3][487] + xnor_result[3][488] + xnor_result[3][489] + xnor_result[3][490] + xnor_result[3][491] + xnor_result[3][492] + xnor_result[3][493] + xnor_result[3][494] + xnor_result[3][495] + xnor_result[3][496] + xnor_result[3][497] + xnor_result[3][498] + xnor_result[3][499] + xnor_result[3][500] + xnor_result[3][501] + xnor_result[3][502] + xnor_result[3][503] + xnor_result[3][504] + xnor_result[3][505] + xnor_result[3][506] + xnor_result[3][507] + xnor_result[3][508] + xnor_result[3][509] + xnor_result[3][510] + xnor_result[3][511] + xnor_result[3][512] + xnor_result[3][513] + xnor_result[3][514] + xnor_result[3][515] + xnor_result[3][516] + xnor_result[3][517] + xnor_result[3][518] + xnor_result[3][519] + xnor_result[3][520] + xnor_result[3][521] + xnor_result[3][522] + xnor_result[3][523] + xnor_result[3][524] + xnor_result[3][525] + xnor_result[3][526] + xnor_result[3][527] + xnor_result[3][528] + xnor_result[3][529] + xnor_result[3][530] + xnor_result[3][531] + xnor_result[3][532] + xnor_result[3][533] + xnor_result[3][534] + xnor_result[3][535] + xnor_result[3][536] + xnor_result[3][537] + xnor_result[3][538] + xnor_result[3][539] + xnor_result[3][540] + xnor_result[3][541] + xnor_result[3][542] + xnor_result[3][543] + xnor_result[3][544] + xnor_result[3][545] + xnor_result[3][546] + xnor_result[3][547] + xnor_result[3][548] + xnor_result[3][549] + xnor_result[3][550] + xnor_result[3][551] + xnor_result[3][552] + xnor_result[3][553] + xnor_result[3][554] + xnor_result[3][555] + xnor_result[3][556] + xnor_result[3][557] + xnor_result[3][558] + xnor_result[3][559] + xnor_result[3][560] + xnor_result[3][561] + xnor_result[3][562] + xnor_result[3][563] + xnor_result[3][564] + xnor_result[3][565] + xnor_result[3][566] + xnor_result[3][567] + xnor_result[3][568] + xnor_result[3][569] + xnor_result[3][570] + xnor_result[3][571] + xnor_result[3][572] + xnor_result[3][573] + xnor_result[3][574] + xnor_result[3][575] + xnor_result[3][576] + xnor_result[3][577] + xnor_result[3][578] + xnor_result[3][579] + xnor_result[3][580] + xnor_result[3][581] + xnor_result[3][582] + xnor_result[3][583] + xnor_result[3][584] + xnor_result[3][585] + xnor_result[3][586] + xnor_result[3][587] + xnor_result[3][588] + xnor_result[3][589] + xnor_result[3][590] + xnor_result[3][591] + xnor_result[3][592] + xnor_result[3][593] + xnor_result[3][594] + xnor_result[3][595] + xnor_result[3][596] + xnor_result[3][597] + xnor_result[3][598] + xnor_result[3][599] + xnor_result[3][600] + xnor_result[3][601] + xnor_result[3][602] + xnor_result[3][603] + xnor_result[3][604] + xnor_result[3][605] + xnor_result[3][606] + xnor_result[3][607] + xnor_result[3][608] + xnor_result[3][609] + xnor_result[3][610] + xnor_result[3][611] + xnor_result[3][612] + xnor_result[3][613] + xnor_result[3][614] + xnor_result[3][615] + xnor_result[3][616] + xnor_result[3][617] + xnor_result[3][618] + xnor_result[3][619] + xnor_result[3][620] + xnor_result[3][621] + xnor_result[3][622] + xnor_result[3][623] + xnor_result[3][624] + xnor_result[3][625] + xnor_result[3][626] + xnor_result[3][627] + xnor_result[3][628] + xnor_result[3][629] + xnor_result[3][630] + xnor_result[3][631] + xnor_result[3][632] + xnor_result[3][633] + xnor_result[3][634] + xnor_result[3][635] + xnor_result[3][636] + xnor_result[3][637] + xnor_result[3][638] + xnor_result[3][639] + xnor_result[3][640] + xnor_result[3][641] + xnor_result[3][642] + xnor_result[3][643] + xnor_result[3][644] + xnor_result[3][645] + xnor_result[3][646] + xnor_result[3][647] + xnor_result[3][648] + xnor_result[3][649] + xnor_result[3][650] + xnor_result[3][651] + xnor_result[3][652] + xnor_result[3][653] + xnor_result[3][654] + xnor_result[3][655] + xnor_result[3][656] + xnor_result[3][657] + xnor_result[3][658] + xnor_result[3][659] + xnor_result[3][660] + xnor_result[3][661] + xnor_result[3][662] + xnor_result[3][663] + xnor_result[3][664] + xnor_result[3][665] + xnor_result[3][666] + xnor_result[3][667] + xnor_result[3][668] + xnor_result[3][669] + xnor_result[3][670] + xnor_result[3][671] + xnor_result[3][672] + xnor_result[3][673] + xnor_result[3][674] + xnor_result[3][675] + xnor_result[3][676] + xnor_result[3][677] + xnor_result[3][678] + xnor_result[3][679] + xnor_result[3][680] + xnor_result[3][681] + xnor_result[3][682] + xnor_result[3][683] + xnor_result[3][684] + xnor_result[3][685] + xnor_result[3][686] + xnor_result[3][687] + xnor_result[3][688] + xnor_result[3][689] + xnor_result[3][690] + xnor_result[3][691] + xnor_result[3][692] + xnor_result[3][693] + xnor_result[3][694] + xnor_result[3][695] + xnor_result[3][696] + xnor_result[3][697] + xnor_result[3][698] + xnor_result[3][699] + xnor_result[3][700] + xnor_result[3][701] + xnor_result[3][702] + xnor_result[3][703] + xnor_result[3][704] + xnor_result[3][705] + xnor_result[3][706] + xnor_result[3][707] + xnor_result[3][708] + xnor_result[3][709] + xnor_result[3][710] + xnor_result[3][711] + xnor_result[3][712] + xnor_result[3][713] + xnor_result[3][714] + xnor_result[3][715] + xnor_result[3][716] + xnor_result[3][717] + xnor_result[3][718] + xnor_result[3][719] + xnor_result[3][720] + xnor_result[3][721] + xnor_result[3][722] + xnor_result[3][723] + xnor_result[3][724] + xnor_result[3][725] + xnor_result[3][726] + xnor_result[3][727] + xnor_result[3][728] + xnor_result[3][729] + xnor_result[3][730] + xnor_result[3][731] + xnor_result[3][732] + xnor_result[3][733] + xnor_result[3][734] + xnor_result[3][735] + xnor_result[3][736] + xnor_result[3][737] + xnor_result[3][738] + xnor_result[3][739] + xnor_result[3][740] + xnor_result[3][741] + xnor_result[3][742] + xnor_result[3][743] + xnor_result[3][744] + xnor_result[3][745] + xnor_result[3][746] + xnor_result[3][747] + xnor_result[3][748] + xnor_result[3][749] + xnor_result[3][750] + xnor_result[3][751] + xnor_result[3][752] + xnor_result[3][753] + xnor_result[3][754] + xnor_result[3][755] + xnor_result[3][756] + xnor_result[3][757] + xnor_result[3][758] + xnor_result[3][759] + xnor_result[3][760] + xnor_result[3][761] + xnor_result[3][762] + xnor_result[3][763] + xnor_result[3][764] + xnor_result[3][765] + xnor_result[3][766] + xnor_result[3][767] + xnor_result[3][768] + xnor_result[3][769] + xnor_result[3][770] + xnor_result[3][771] + xnor_result[3][772] + xnor_result[3][773] + xnor_result[3][774] + xnor_result[3][775] + xnor_result[3][776] + xnor_result[3][777] + xnor_result[3][778] + xnor_result[3][779] + xnor_result[3][780] + xnor_result[3][781] + xnor_result[3][782] + xnor_result[3][783] + xnor_result[3][784] + xnor_result[3][785] + xnor_result[3][786] + xnor_result[3][787] + xnor_result[3][788] + xnor_result[3][789] + xnor_result[3][790] + xnor_result[3][791] + xnor_result[3][792] + xnor_result[3][793] + xnor_result[3][794] + xnor_result[3][795] + xnor_result[3][796] + xnor_result[3][797] + xnor_result[3][798] + xnor_result[3][799] + xnor_result[3][800] + xnor_result[3][801] + xnor_result[3][802] + xnor_result[3][803] + xnor_result[3][804] + xnor_result[3][805] + xnor_result[3][806] + xnor_result[3][807] + xnor_result[3][808] + xnor_result[3][809] + xnor_result[3][810] + xnor_result[3][811] + xnor_result[3][812] + xnor_result[3][813] + xnor_result[3][814] + xnor_result[3][815] + xnor_result[3][816] + xnor_result[3][817] + xnor_result[3][818] + xnor_result[3][819] + xnor_result[3][820] + xnor_result[3][821] + xnor_result[3][822] + xnor_result[3][823] + xnor_result[3][824] + xnor_result[3][825] + xnor_result[3][826] + xnor_result[3][827] + xnor_result[3][828] + xnor_result[3][829] + xnor_result[3][830] + xnor_result[3][831] + xnor_result[3][832] + xnor_result[3][833] + xnor_result[3][834] + xnor_result[3][835] + xnor_result[3][836] + xnor_result[3][837] + xnor_result[3][838] + xnor_result[3][839] + xnor_result[3][840] + xnor_result[3][841] + xnor_result[3][842] + xnor_result[3][843] + xnor_result[3][844] + xnor_result[3][845] + xnor_result[3][846] + xnor_result[3][847] + xnor_result[3][848] + xnor_result[3][849] + xnor_result[3][850] + xnor_result[3][851] + xnor_result[3][852] + xnor_result[3][853] + xnor_result[3][854] + xnor_result[3][855] + xnor_result[3][856] + xnor_result[3][857] + xnor_result[3][858] + xnor_result[3][859] + xnor_result[3][860] + xnor_result[3][861] + xnor_result[3][862] + xnor_result[3][863] + xnor_result[3][864] + xnor_result[3][865] + xnor_result[3][866] + xnor_result[3][867] + xnor_result[3][868] + xnor_result[3][869] + xnor_result[3][870] + xnor_result[3][871] + xnor_result[3][872] + xnor_result[3][873] + xnor_result[3][874] + xnor_result[3][875] + xnor_result[3][876] + xnor_result[3][877] + xnor_result[3][878] + xnor_result[3][879] + xnor_result[3][880] + xnor_result[3][881] + xnor_result[3][882] + xnor_result[3][883] + xnor_result[3][884] + xnor_result[3][885] + xnor_result[3][886] + xnor_result[3][887] + xnor_result[3][888] + xnor_result[3][889] + xnor_result[3][890] + xnor_result[3][891] + xnor_result[3][892] + xnor_result[3][893] + xnor_result[3][894] + xnor_result[3][895] + xnor_result[3][896] + xnor_result[3][897] + xnor_result[3][898] + xnor_result[3][899] + xnor_result[3][900] + xnor_result[3][901] + xnor_result[3][902] + xnor_result[3][903] + xnor_result[3][904] + xnor_result[3][905] + xnor_result[3][906] + xnor_result[3][907] + xnor_result[3][908] + xnor_result[3][909] + xnor_result[3][910] + xnor_result[3][911] + xnor_result[3][912] + xnor_result[3][913] + xnor_result[3][914] + xnor_result[3][915] + xnor_result[3][916] + xnor_result[3][917] + xnor_result[3][918] + xnor_result[3][919] + xnor_result[3][920] + xnor_result[3][921] + xnor_result[3][922] + xnor_result[3][923] + xnor_result[3][924] + xnor_result[3][925] + xnor_result[3][926] + xnor_result[3][927] + xnor_result[3][928] + xnor_result[3][929] + xnor_result[3][930] + xnor_result[3][931] + xnor_result[3][932] + xnor_result[3][933] + xnor_result[3][934] + xnor_result[3][935] + xnor_result[3][936] + xnor_result[3][937] + xnor_result[3][938] + xnor_result[3][939] + xnor_result[3][940] + xnor_result[3][941] + xnor_result[3][942] + xnor_result[3][943] + xnor_result[3][944] + xnor_result[3][945] + xnor_result[3][946] + xnor_result[3][947] + xnor_result[3][948] + xnor_result[3][949] + xnor_result[3][950] + xnor_result[3][951] + xnor_result[3][952] + xnor_result[3][953] + xnor_result[3][954] + xnor_result[3][955] + xnor_result[3][956] + xnor_result[3][957] + xnor_result[3][958] + xnor_result[3][959] ;
assign accumulation_result[4] = xnor_result[4][0] + xnor_result[4][1] + xnor_result[4][2] + xnor_result[4][3] + xnor_result[4][4] + xnor_result[4][5] + xnor_result[4][6] + xnor_result[4][7] + xnor_result[4][8] + xnor_result[4][9] + xnor_result[4][10] + xnor_result[4][11] + xnor_result[4][12] + xnor_result[4][13] + xnor_result[4][14] + xnor_result[4][15] + xnor_result[4][16] + xnor_result[4][17] + xnor_result[4][18] + xnor_result[4][19] + xnor_result[4][20] + xnor_result[4][21] + xnor_result[4][22] + xnor_result[4][23] + xnor_result[4][24] + xnor_result[4][25] + xnor_result[4][26] + xnor_result[4][27] + xnor_result[4][28] + xnor_result[4][29] + xnor_result[4][30] + xnor_result[4][31] + xnor_result[4][32] + xnor_result[4][33] + xnor_result[4][34] + xnor_result[4][35] + xnor_result[4][36] + xnor_result[4][37] + xnor_result[4][38] + xnor_result[4][39] + xnor_result[4][40] + xnor_result[4][41] + xnor_result[4][42] + xnor_result[4][43] + xnor_result[4][44] + xnor_result[4][45] + xnor_result[4][46] + xnor_result[4][47] + xnor_result[4][48] + xnor_result[4][49] + xnor_result[4][50] + xnor_result[4][51] + xnor_result[4][52] + xnor_result[4][53] + xnor_result[4][54] + xnor_result[4][55] + xnor_result[4][56] + xnor_result[4][57] + xnor_result[4][58] + xnor_result[4][59] + xnor_result[4][60] + xnor_result[4][61] + xnor_result[4][62] + xnor_result[4][63] + xnor_result[4][64] + xnor_result[4][65] + xnor_result[4][66] + xnor_result[4][67] + xnor_result[4][68] + xnor_result[4][69] + xnor_result[4][70] + xnor_result[4][71] + xnor_result[4][72] + xnor_result[4][73] + xnor_result[4][74] + xnor_result[4][75] + xnor_result[4][76] + xnor_result[4][77] + xnor_result[4][78] + xnor_result[4][79] + xnor_result[4][80] + xnor_result[4][81] + xnor_result[4][82] + xnor_result[4][83] + xnor_result[4][84] + xnor_result[4][85] + xnor_result[4][86] + xnor_result[4][87] + xnor_result[4][88] + xnor_result[4][89] + xnor_result[4][90] + xnor_result[4][91] + xnor_result[4][92] + xnor_result[4][93] + xnor_result[4][94] + xnor_result[4][95] + xnor_result[4][96] + xnor_result[4][97] + xnor_result[4][98] + xnor_result[4][99] + xnor_result[4][100] + xnor_result[4][101] + xnor_result[4][102] + xnor_result[4][103] + xnor_result[4][104] + xnor_result[4][105] + xnor_result[4][106] + xnor_result[4][107] + xnor_result[4][108] + xnor_result[4][109] + xnor_result[4][110] + xnor_result[4][111] + xnor_result[4][112] + xnor_result[4][113] + xnor_result[4][114] + xnor_result[4][115] + xnor_result[4][116] + xnor_result[4][117] + xnor_result[4][118] + xnor_result[4][119] + xnor_result[4][120] + xnor_result[4][121] + xnor_result[4][122] + xnor_result[4][123] + xnor_result[4][124] + xnor_result[4][125] + xnor_result[4][126] + xnor_result[4][127] + xnor_result[4][128] + xnor_result[4][129] + xnor_result[4][130] + xnor_result[4][131] + xnor_result[4][132] + xnor_result[4][133] + xnor_result[4][134] + xnor_result[4][135] + xnor_result[4][136] + xnor_result[4][137] + xnor_result[4][138] + xnor_result[4][139] + xnor_result[4][140] + xnor_result[4][141] + xnor_result[4][142] + xnor_result[4][143] + xnor_result[4][144] + xnor_result[4][145] + xnor_result[4][146] + xnor_result[4][147] + xnor_result[4][148] + xnor_result[4][149] + xnor_result[4][150] + xnor_result[4][151] + xnor_result[4][152] + xnor_result[4][153] + xnor_result[4][154] + xnor_result[4][155] + xnor_result[4][156] + xnor_result[4][157] + xnor_result[4][158] + xnor_result[4][159] + xnor_result[4][160] + xnor_result[4][161] + xnor_result[4][162] + xnor_result[4][163] + xnor_result[4][164] + xnor_result[4][165] + xnor_result[4][166] + xnor_result[4][167] + xnor_result[4][168] + xnor_result[4][169] + xnor_result[4][170] + xnor_result[4][171] + xnor_result[4][172] + xnor_result[4][173] + xnor_result[4][174] + xnor_result[4][175] + xnor_result[4][176] + xnor_result[4][177] + xnor_result[4][178] + xnor_result[4][179] + xnor_result[4][180] + xnor_result[4][181] + xnor_result[4][182] + xnor_result[4][183] + xnor_result[4][184] + xnor_result[4][185] + xnor_result[4][186] + xnor_result[4][187] + xnor_result[4][188] + xnor_result[4][189] + xnor_result[4][190] + xnor_result[4][191] + xnor_result[4][192] + xnor_result[4][193] + xnor_result[4][194] + xnor_result[4][195] + xnor_result[4][196] + xnor_result[4][197] + xnor_result[4][198] + xnor_result[4][199] + xnor_result[4][200] + xnor_result[4][201] + xnor_result[4][202] + xnor_result[4][203] + xnor_result[4][204] + xnor_result[4][205] + xnor_result[4][206] + xnor_result[4][207] + xnor_result[4][208] + xnor_result[4][209] + xnor_result[4][210] + xnor_result[4][211] + xnor_result[4][212] + xnor_result[4][213] + xnor_result[4][214] + xnor_result[4][215] + xnor_result[4][216] + xnor_result[4][217] + xnor_result[4][218] + xnor_result[4][219] + xnor_result[4][220] + xnor_result[4][221] + xnor_result[4][222] + xnor_result[4][223] + xnor_result[4][224] + xnor_result[4][225] + xnor_result[4][226] + xnor_result[4][227] + xnor_result[4][228] + xnor_result[4][229] + xnor_result[4][230] + xnor_result[4][231] + xnor_result[4][232] + xnor_result[4][233] + xnor_result[4][234] + xnor_result[4][235] + xnor_result[4][236] + xnor_result[4][237] + xnor_result[4][238] + xnor_result[4][239] + xnor_result[4][240] + xnor_result[4][241] + xnor_result[4][242] + xnor_result[4][243] + xnor_result[4][244] + xnor_result[4][245] + xnor_result[4][246] + xnor_result[4][247] + xnor_result[4][248] + xnor_result[4][249] + xnor_result[4][250] + xnor_result[4][251] + xnor_result[4][252] + xnor_result[4][253] + xnor_result[4][254] + xnor_result[4][255] + xnor_result[4][256] + xnor_result[4][257] + xnor_result[4][258] + xnor_result[4][259] + xnor_result[4][260] + xnor_result[4][261] + xnor_result[4][262] + xnor_result[4][263] + xnor_result[4][264] + xnor_result[4][265] + xnor_result[4][266] + xnor_result[4][267] + xnor_result[4][268] + xnor_result[4][269] + xnor_result[4][270] + xnor_result[4][271] + xnor_result[4][272] + xnor_result[4][273] + xnor_result[4][274] + xnor_result[4][275] + xnor_result[4][276] + xnor_result[4][277] + xnor_result[4][278] + xnor_result[4][279] + xnor_result[4][280] + xnor_result[4][281] + xnor_result[4][282] + xnor_result[4][283] + xnor_result[4][284] + xnor_result[4][285] + xnor_result[4][286] + xnor_result[4][287] + xnor_result[4][288] + xnor_result[4][289] + xnor_result[4][290] + xnor_result[4][291] + xnor_result[4][292] + xnor_result[4][293] + xnor_result[4][294] + xnor_result[4][295] + xnor_result[4][296] + xnor_result[4][297] + xnor_result[4][298] + xnor_result[4][299] + xnor_result[4][300] + xnor_result[4][301] + xnor_result[4][302] + xnor_result[4][303] + xnor_result[4][304] + xnor_result[4][305] + xnor_result[4][306] + xnor_result[4][307] + xnor_result[4][308] + xnor_result[4][309] + xnor_result[4][310] + xnor_result[4][311] + xnor_result[4][312] + xnor_result[4][313] + xnor_result[4][314] + xnor_result[4][315] + xnor_result[4][316] + xnor_result[4][317] + xnor_result[4][318] + xnor_result[4][319] + xnor_result[4][320] + xnor_result[4][321] + xnor_result[4][322] + xnor_result[4][323] + xnor_result[4][324] + xnor_result[4][325] + xnor_result[4][326] + xnor_result[4][327] + xnor_result[4][328] + xnor_result[4][329] + xnor_result[4][330] + xnor_result[4][331] + xnor_result[4][332] + xnor_result[4][333] + xnor_result[4][334] + xnor_result[4][335] + xnor_result[4][336] + xnor_result[4][337] + xnor_result[4][338] + xnor_result[4][339] + xnor_result[4][340] + xnor_result[4][341] + xnor_result[4][342] + xnor_result[4][343] + xnor_result[4][344] + xnor_result[4][345] + xnor_result[4][346] + xnor_result[4][347] + xnor_result[4][348] + xnor_result[4][349] + xnor_result[4][350] + xnor_result[4][351] + xnor_result[4][352] + xnor_result[4][353] + xnor_result[4][354] + xnor_result[4][355] + xnor_result[4][356] + xnor_result[4][357] + xnor_result[4][358] + xnor_result[4][359] + xnor_result[4][360] + xnor_result[4][361] + xnor_result[4][362] + xnor_result[4][363] + xnor_result[4][364] + xnor_result[4][365] + xnor_result[4][366] + xnor_result[4][367] + xnor_result[4][368] + xnor_result[4][369] + xnor_result[4][370] + xnor_result[4][371] + xnor_result[4][372] + xnor_result[4][373] + xnor_result[4][374] + xnor_result[4][375] + xnor_result[4][376] + xnor_result[4][377] + xnor_result[4][378] + xnor_result[4][379] + xnor_result[4][380] + xnor_result[4][381] + xnor_result[4][382] + xnor_result[4][383] + xnor_result[4][384] + xnor_result[4][385] + xnor_result[4][386] + xnor_result[4][387] + xnor_result[4][388] + xnor_result[4][389] + xnor_result[4][390] + xnor_result[4][391] + xnor_result[4][392] + xnor_result[4][393] + xnor_result[4][394] + xnor_result[4][395] + xnor_result[4][396] + xnor_result[4][397] + xnor_result[4][398] + xnor_result[4][399] + xnor_result[4][400] + xnor_result[4][401] + xnor_result[4][402] + xnor_result[4][403] + xnor_result[4][404] + xnor_result[4][405] + xnor_result[4][406] + xnor_result[4][407] + xnor_result[4][408] + xnor_result[4][409] + xnor_result[4][410] + xnor_result[4][411] + xnor_result[4][412] + xnor_result[4][413] + xnor_result[4][414] + xnor_result[4][415] + xnor_result[4][416] + xnor_result[4][417] + xnor_result[4][418] + xnor_result[4][419] + xnor_result[4][420] + xnor_result[4][421] + xnor_result[4][422] + xnor_result[4][423] + xnor_result[4][424] + xnor_result[4][425] + xnor_result[4][426] + xnor_result[4][427] + xnor_result[4][428] + xnor_result[4][429] + xnor_result[4][430] + xnor_result[4][431] + xnor_result[4][432] + xnor_result[4][433] + xnor_result[4][434] + xnor_result[4][435] + xnor_result[4][436] + xnor_result[4][437] + xnor_result[4][438] + xnor_result[4][439] + xnor_result[4][440] + xnor_result[4][441] + xnor_result[4][442] + xnor_result[4][443] + xnor_result[4][444] + xnor_result[4][445] + xnor_result[4][446] + xnor_result[4][447] + xnor_result[4][448] + xnor_result[4][449] + xnor_result[4][450] + xnor_result[4][451] + xnor_result[4][452] + xnor_result[4][453] + xnor_result[4][454] + xnor_result[4][455] + xnor_result[4][456] + xnor_result[4][457] + xnor_result[4][458] + xnor_result[4][459] + xnor_result[4][460] + xnor_result[4][461] + xnor_result[4][462] + xnor_result[4][463] + xnor_result[4][464] + xnor_result[4][465] + xnor_result[4][466] + xnor_result[4][467] + xnor_result[4][468] + xnor_result[4][469] + xnor_result[4][470] + xnor_result[4][471] + xnor_result[4][472] + xnor_result[4][473] + xnor_result[4][474] + xnor_result[4][475] + xnor_result[4][476] + xnor_result[4][477] + xnor_result[4][478] + xnor_result[4][479] + xnor_result[4][480] + xnor_result[4][481] + xnor_result[4][482] + xnor_result[4][483] + xnor_result[4][484] + xnor_result[4][485] + xnor_result[4][486] + xnor_result[4][487] + xnor_result[4][488] + xnor_result[4][489] + xnor_result[4][490] + xnor_result[4][491] + xnor_result[4][492] + xnor_result[4][493] + xnor_result[4][494] + xnor_result[4][495] + xnor_result[4][496] + xnor_result[4][497] + xnor_result[4][498] + xnor_result[4][499] + xnor_result[4][500] + xnor_result[4][501] + xnor_result[4][502] + xnor_result[4][503] + xnor_result[4][504] + xnor_result[4][505] + xnor_result[4][506] + xnor_result[4][507] + xnor_result[4][508] + xnor_result[4][509] + xnor_result[4][510] + xnor_result[4][511] + xnor_result[4][512] + xnor_result[4][513] + xnor_result[4][514] + xnor_result[4][515] + xnor_result[4][516] + xnor_result[4][517] + xnor_result[4][518] + xnor_result[4][519] + xnor_result[4][520] + xnor_result[4][521] + xnor_result[4][522] + xnor_result[4][523] + xnor_result[4][524] + xnor_result[4][525] + xnor_result[4][526] + xnor_result[4][527] + xnor_result[4][528] + xnor_result[4][529] + xnor_result[4][530] + xnor_result[4][531] + xnor_result[4][532] + xnor_result[4][533] + xnor_result[4][534] + xnor_result[4][535] + xnor_result[4][536] + xnor_result[4][537] + xnor_result[4][538] + xnor_result[4][539] + xnor_result[4][540] + xnor_result[4][541] + xnor_result[4][542] + xnor_result[4][543] + xnor_result[4][544] + xnor_result[4][545] + xnor_result[4][546] + xnor_result[4][547] + xnor_result[4][548] + xnor_result[4][549] + xnor_result[4][550] + xnor_result[4][551] + xnor_result[4][552] + xnor_result[4][553] + xnor_result[4][554] + xnor_result[4][555] + xnor_result[4][556] + xnor_result[4][557] + xnor_result[4][558] + xnor_result[4][559] + xnor_result[4][560] + xnor_result[4][561] + xnor_result[4][562] + xnor_result[4][563] + xnor_result[4][564] + xnor_result[4][565] + xnor_result[4][566] + xnor_result[4][567] + xnor_result[4][568] + xnor_result[4][569] + xnor_result[4][570] + xnor_result[4][571] + xnor_result[4][572] + xnor_result[4][573] + xnor_result[4][574] + xnor_result[4][575] + xnor_result[4][576] + xnor_result[4][577] + xnor_result[4][578] + xnor_result[4][579] + xnor_result[4][580] + xnor_result[4][581] + xnor_result[4][582] + xnor_result[4][583] + xnor_result[4][584] + xnor_result[4][585] + xnor_result[4][586] + xnor_result[4][587] + xnor_result[4][588] + xnor_result[4][589] + xnor_result[4][590] + xnor_result[4][591] + xnor_result[4][592] + xnor_result[4][593] + xnor_result[4][594] + xnor_result[4][595] + xnor_result[4][596] + xnor_result[4][597] + xnor_result[4][598] + xnor_result[4][599] + xnor_result[4][600] + xnor_result[4][601] + xnor_result[4][602] + xnor_result[4][603] + xnor_result[4][604] + xnor_result[4][605] + xnor_result[4][606] + xnor_result[4][607] + xnor_result[4][608] + xnor_result[4][609] + xnor_result[4][610] + xnor_result[4][611] + xnor_result[4][612] + xnor_result[4][613] + xnor_result[4][614] + xnor_result[4][615] + xnor_result[4][616] + xnor_result[4][617] + xnor_result[4][618] + xnor_result[4][619] + xnor_result[4][620] + xnor_result[4][621] + xnor_result[4][622] + xnor_result[4][623] + xnor_result[4][624] + xnor_result[4][625] + xnor_result[4][626] + xnor_result[4][627] + xnor_result[4][628] + xnor_result[4][629] + xnor_result[4][630] + xnor_result[4][631] + xnor_result[4][632] + xnor_result[4][633] + xnor_result[4][634] + xnor_result[4][635] + xnor_result[4][636] + xnor_result[4][637] + xnor_result[4][638] + xnor_result[4][639] + xnor_result[4][640] + xnor_result[4][641] + xnor_result[4][642] + xnor_result[4][643] + xnor_result[4][644] + xnor_result[4][645] + xnor_result[4][646] + xnor_result[4][647] + xnor_result[4][648] + xnor_result[4][649] + xnor_result[4][650] + xnor_result[4][651] + xnor_result[4][652] + xnor_result[4][653] + xnor_result[4][654] + xnor_result[4][655] + xnor_result[4][656] + xnor_result[4][657] + xnor_result[4][658] + xnor_result[4][659] + xnor_result[4][660] + xnor_result[4][661] + xnor_result[4][662] + xnor_result[4][663] + xnor_result[4][664] + xnor_result[4][665] + xnor_result[4][666] + xnor_result[4][667] + xnor_result[4][668] + xnor_result[4][669] + xnor_result[4][670] + xnor_result[4][671] + xnor_result[4][672] + xnor_result[4][673] + xnor_result[4][674] + xnor_result[4][675] + xnor_result[4][676] + xnor_result[4][677] + xnor_result[4][678] + xnor_result[4][679] + xnor_result[4][680] + xnor_result[4][681] + xnor_result[4][682] + xnor_result[4][683] + xnor_result[4][684] + xnor_result[4][685] + xnor_result[4][686] + xnor_result[4][687] + xnor_result[4][688] + xnor_result[4][689] + xnor_result[4][690] + xnor_result[4][691] + xnor_result[4][692] + xnor_result[4][693] + xnor_result[4][694] + xnor_result[4][695] + xnor_result[4][696] + xnor_result[4][697] + xnor_result[4][698] + xnor_result[4][699] + xnor_result[4][700] + xnor_result[4][701] + xnor_result[4][702] + xnor_result[4][703] + xnor_result[4][704] + xnor_result[4][705] + xnor_result[4][706] + xnor_result[4][707] + xnor_result[4][708] + xnor_result[4][709] + xnor_result[4][710] + xnor_result[4][711] + xnor_result[4][712] + xnor_result[4][713] + xnor_result[4][714] + xnor_result[4][715] + xnor_result[4][716] + xnor_result[4][717] + xnor_result[4][718] + xnor_result[4][719] + xnor_result[4][720] + xnor_result[4][721] + xnor_result[4][722] + xnor_result[4][723] + xnor_result[4][724] + xnor_result[4][725] + xnor_result[4][726] + xnor_result[4][727] + xnor_result[4][728] + xnor_result[4][729] + xnor_result[4][730] + xnor_result[4][731] + xnor_result[4][732] + xnor_result[4][733] + xnor_result[4][734] + xnor_result[4][735] + xnor_result[4][736] + xnor_result[4][737] + xnor_result[4][738] + xnor_result[4][739] + xnor_result[4][740] + xnor_result[4][741] + xnor_result[4][742] + xnor_result[4][743] + xnor_result[4][744] + xnor_result[4][745] + xnor_result[4][746] + xnor_result[4][747] + xnor_result[4][748] + xnor_result[4][749] + xnor_result[4][750] + xnor_result[4][751] + xnor_result[4][752] + xnor_result[4][753] + xnor_result[4][754] + xnor_result[4][755] + xnor_result[4][756] + xnor_result[4][757] + xnor_result[4][758] + xnor_result[4][759] + xnor_result[4][760] + xnor_result[4][761] + xnor_result[4][762] + xnor_result[4][763] + xnor_result[4][764] + xnor_result[4][765] + xnor_result[4][766] + xnor_result[4][767] + xnor_result[4][768] + xnor_result[4][769] + xnor_result[4][770] + xnor_result[4][771] + xnor_result[4][772] + xnor_result[4][773] + xnor_result[4][774] + xnor_result[4][775] + xnor_result[4][776] + xnor_result[4][777] + xnor_result[4][778] + xnor_result[4][779] + xnor_result[4][780] + xnor_result[4][781] + xnor_result[4][782] + xnor_result[4][783] + xnor_result[4][784] + xnor_result[4][785] + xnor_result[4][786] + xnor_result[4][787] + xnor_result[4][788] + xnor_result[4][789] + xnor_result[4][790] + xnor_result[4][791] + xnor_result[4][792] + xnor_result[4][793] + xnor_result[4][794] + xnor_result[4][795] + xnor_result[4][796] + xnor_result[4][797] + xnor_result[4][798] + xnor_result[4][799] + xnor_result[4][800] + xnor_result[4][801] + xnor_result[4][802] + xnor_result[4][803] + xnor_result[4][804] + xnor_result[4][805] + xnor_result[4][806] + xnor_result[4][807] + xnor_result[4][808] + xnor_result[4][809] + xnor_result[4][810] + xnor_result[4][811] + xnor_result[4][812] + xnor_result[4][813] + xnor_result[4][814] + xnor_result[4][815] + xnor_result[4][816] + xnor_result[4][817] + xnor_result[4][818] + xnor_result[4][819] + xnor_result[4][820] + xnor_result[4][821] + xnor_result[4][822] + xnor_result[4][823] + xnor_result[4][824] + xnor_result[4][825] + xnor_result[4][826] + xnor_result[4][827] + xnor_result[4][828] + xnor_result[4][829] + xnor_result[4][830] + xnor_result[4][831] + xnor_result[4][832] + xnor_result[4][833] + xnor_result[4][834] + xnor_result[4][835] + xnor_result[4][836] + xnor_result[4][837] + xnor_result[4][838] + xnor_result[4][839] + xnor_result[4][840] + xnor_result[4][841] + xnor_result[4][842] + xnor_result[4][843] + xnor_result[4][844] + xnor_result[4][845] + xnor_result[4][846] + xnor_result[4][847] + xnor_result[4][848] + xnor_result[4][849] + xnor_result[4][850] + xnor_result[4][851] + xnor_result[4][852] + xnor_result[4][853] + xnor_result[4][854] + xnor_result[4][855] + xnor_result[4][856] + xnor_result[4][857] + xnor_result[4][858] + xnor_result[4][859] + xnor_result[4][860] + xnor_result[4][861] + xnor_result[4][862] + xnor_result[4][863] + xnor_result[4][864] + xnor_result[4][865] + xnor_result[4][866] + xnor_result[4][867] + xnor_result[4][868] + xnor_result[4][869] + xnor_result[4][870] + xnor_result[4][871] + xnor_result[4][872] + xnor_result[4][873] + xnor_result[4][874] + xnor_result[4][875] + xnor_result[4][876] + xnor_result[4][877] + xnor_result[4][878] + xnor_result[4][879] + xnor_result[4][880] + xnor_result[4][881] + xnor_result[4][882] + xnor_result[4][883] + xnor_result[4][884] + xnor_result[4][885] + xnor_result[4][886] + xnor_result[4][887] + xnor_result[4][888] + xnor_result[4][889] + xnor_result[4][890] + xnor_result[4][891] + xnor_result[4][892] + xnor_result[4][893] + xnor_result[4][894] + xnor_result[4][895] + xnor_result[4][896] + xnor_result[4][897] + xnor_result[4][898] + xnor_result[4][899] + xnor_result[4][900] + xnor_result[4][901] + xnor_result[4][902] + xnor_result[4][903] + xnor_result[4][904] + xnor_result[4][905] + xnor_result[4][906] + xnor_result[4][907] + xnor_result[4][908] + xnor_result[4][909] + xnor_result[4][910] + xnor_result[4][911] + xnor_result[4][912] + xnor_result[4][913] + xnor_result[4][914] + xnor_result[4][915] + xnor_result[4][916] + xnor_result[4][917] + xnor_result[4][918] + xnor_result[4][919] + xnor_result[4][920] + xnor_result[4][921] + xnor_result[4][922] + xnor_result[4][923] + xnor_result[4][924] + xnor_result[4][925] + xnor_result[4][926] + xnor_result[4][927] + xnor_result[4][928] + xnor_result[4][929] + xnor_result[4][930] + xnor_result[4][931] + xnor_result[4][932] + xnor_result[4][933] + xnor_result[4][934] + xnor_result[4][935] + xnor_result[4][936] + xnor_result[4][937] + xnor_result[4][938] + xnor_result[4][939] + xnor_result[4][940] + xnor_result[4][941] + xnor_result[4][942] + xnor_result[4][943] + xnor_result[4][944] + xnor_result[4][945] + xnor_result[4][946] + xnor_result[4][947] + xnor_result[4][948] + xnor_result[4][949] + xnor_result[4][950] + xnor_result[4][951] + xnor_result[4][952] + xnor_result[4][953] + xnor_result[4][954] + xnor_result[4][955] + xnor_result[4][956] + xnor_result[4][957] + xnor_result[4][958] + xnor_result[4][959] ;
assign accumulation_result[5] = xnor_result[5][0] + xnor_result[5][1] + xnor_result[5][2] + xnor_result[5][3] + xnor_result[5][4] + xnor_result[5][5] + xnor_result[5][6] + xnor_result[5][7] + xnor_result[5][8] + xnor_result[5][9] + xnor_result[5][10] + xnor_result[5][11] + xnor_result[5][12] + xnor_result[5][13] + xnor_result[5][14] + xnor_result[5][15] + xnor_result[5][16] + xnor_result[5][17] + xnor_result[5][18] + xnor_result[5][19] + xnor_result[5][20] + xnor_result[5][21] + xnor_result[5][22] + xnor_result[5][23] + xnor_result[5][24] + xnor_result[5][25] + xnor_result[5][26] + xnor_result[5][27] + xnor_result[5][28] + xnor_result[5][29] + xnor_result[5][30] + xnor_result[5][31] + xnor_result[5][32] + xnor_result[5][33] + xnor_result[5][34] + xnor_result[5][35] + xnor_result[5][36] + xnor_result[5][37] + xnor_result[5][38] + xnor_result[5][39] + xnor_result[5][40] + xnor_result[5][41] + xnor_result[5][42] + xnor_result[5][43] + xnor_result[5][44] + xnor_result[5][45] + xnor_result[5][46] + xnor_result[5][47] + xnor_result[5][48] + xnor_result[5][49] + xnor_result[5][50] + xnor_result[5][51] + xnor_result[5][52] + xnor_result[5][53] + xnor_result[5][54] + xnor_result[5][55] + xnor_result[5][56] + xnor_result[5][57] + xnor_result[5][58] + xnor_result[5][59] + xnor_result[5][60] + xnor_result[5][61] + xnor_result[5][62] + xnor_result[5][63] + xnor_result[5][64] + xnor_result[5][65] + xnor_result[5][66] + xnor_result[5][67] + xnor_result[5][68] + xnor_result[5][69] + xnor_result[5][70] + xnor_result[5][71] + xnor_result[5][72] + xnor_result[5][73] + xnor_result[5][74] + xnor_result[5][75] + xnor_result[5][76] + xnor_result[5][77] + xnor_result[5][78] + xnor_result[5][79] + xnor_result[5][80] + xnor_result[5][81] + xnor_result[5][82] + xnor_result[5][83] + xnor_result[5][84] + xnor_result[5][85] + xnor_result[5][86] + xnor_result[5][87] + xnor_result[5][88] + xnor_result[5][89] + xnor_result[5][90] + xnor_result[5][91] + xnor_result[5][92] + xnor_result[5][93] + xnor_result[5][94] + xnor_result[5][95] + xnor_result[5][96] + xnor_result[5][97] + xnor_result[5][98] + xnor_result[5][99] + xnor_result[5][100] + xnor_result[5][101] + xnor_result[5][102] + xnor_result[5][103] + xnor_result[5][104] + xnor_result[5][105] + xnor_result[5][106] + xnor_result[5][107] + xnor_result[5][108] + xnor_result[5][109] + xnor_result[5][110] + xnor_result[5][111] + xnor_result[5][112] + xnor_result[5][113] + xnor_result[5][114] + xnor_result[5][115] + xnor_result[5][116] + xnor_result[5][117] + xnor_result[5][118] + xnor_result[5][119] + xnor_result[5][120] + xnor_result[5][121] + xnor_result[5][122] + xnor_result[5][123] + xnor_result[5][124] + xnor_result[5][125] + xnor_result[5][126] + xnor_result[5][127] + xnor_result[5][128] + xnor_result[5][129] + xnor_result[5][130] + xnor_result[5][131] + xnor_result[5][132] + xnor_result[5][133] + xnor_result[5][134] + xnor_result[5][135] + xnor_result[5][136] + xnor_result[5][137] + xnor_result[5][138] + xnor_result[5][139] + xnor_result[5][140] + xnor_result[5][141] + xnor_result[5][142] + xnor_result[5][143] + xnor_result[5][144] + xnor_result[5][145] + xnor_result[5][146] + xnor_result[5][147] + xnor_result[5][148] + xnor_result[5][149] + xnor_result[5][150] + xnor_result[5][151] + xnor_result[5][152] + xnor_result[5][153] + xnor_result[5][154] + xnor_result[5][155] + xnor_result[5][156] + xnor_result[5][157] + xnor_result[5][158] + xnor_result[5][159] + xnor_result[5][160] + xnor_result[5][161] + xnor_result[5][162] + xnor_result[5][163] + xnor_result[5][164] + xnor_result[5][165] + xnor_result[5][166] + xnor_result[5][167] + xnor_result[5][168] + xnor_result[5][169] + xnor_result[5][170] + xnor_result[5][171] + xnor_result[5][172] + xnor_result[5][173] + xnor_result[5][174] + xnor_result[5][175] + xnor_result[5][176] + xnor_result[5][177] + xnor_result[5][178] + xnor_result[5][179] + xnor_result[5][180] + xnor_result[5][181] + xnor_result[5][182] + xnor_result[5][183] + xnor_result[5][184] + xnor_result[5][185] + xnor_result[5][186] + xnor_result[5][187] + xnor_result[5][188] + xnor_result[5][189] + xnor_result[5][190] + xnor_result[5][191] + xnor_result[5][192] + xnor_result[5][193] + xnor_result[5][194] + xnor_result[5][195] + xnor_result[5][196] + xnor_result[5][197] + xnor_result[5][198] + xnor_result[5][199] + xnor_result[5][200] + xnor_result[5][201] + xnor_result[5][202] + xnor_result[5][203] + xnor_result[5][204] + xnor_result[5][205] + xnor_result[5][206] + xnor_result[5][207] + xnor_result[5][208] + xnor_result[5][209] + xnor_result[5][210] + xnor_result[5][211] + xnor_result[5][212] + xnor_result[5][213] + xnor_result[5][214] + xnor_result[5][215] + xnor_result[5][216] + xnor_result[5][217] + xnor_result[5][218] + xnor_result[5][219] + xnor_result[5][220] + xnor_result[5][221] + xnor_result[5][222] + xnor_result[5][223] + xnor_result[5][224] + xnor_result[5][225] + xnor_result[5][226] + xnor_result[5][227] + xnor_result[5][228] + xnor_result[5][229] + xnor_result[5][230] + xnor_result[5][231] + xnor_result[5][232] + xnor_result[5][233] + xnor_result[5][234] + xnor_result[5][235] + xnor_result[5][236] + xnor_result[5][237] + xnor_result[5][238] + xnor_result[5][239] + xnor_result[5][240] + xnor_result[5][241] + xnor_result[5][242] + xnor_result[5][243] + xnor_result[5][244] + xnor_result[5][245] + xnor_result[5][246] + xnor_result[5][247] + xnor_result[5][248] + xnor_result[5][249] + xnor_result[5][250] + xnor_result[5][251] + xnor_result[5][252] + xnor_result[5][253] + xnor_result[5][254] + xnor_result[5][255] + xnor_result[5][256] + xnor_result[5][257] + xnor_result[5][258] + xnor_result[5][259] + xnor_result[5][260] + xnor_result[5][261] + xnor_result[5][262] + xnor_result[5][263] + xnor_result[5][264] + xnor_result[5][265] + xnor_result[5][266] + xnor_result[5][267] + xnor_result[5][268] + xnor_result[5][269] + xnor_result[5][270] + xnor_result[5][271] + xnor_result[5][272] + xnor_result[5][273] + xnor_result[5][274] + xnor_result[5][275] + xnor_result[5][276] + xnor_result[5][277] + xnor_result[5][278] + xnor_result[5][279] + xnor_result[5][280] + xnor_result[5][281] + xnor_result[5][282] + xnor_result[5][283] + xnor_result[5][284] + xnor_result[5][285] + xnor_result[5][286] + xnor_result[5][287] + xnor_result[5][288] + xnor_result[5][289] + xnor_result[5][290] + xnor_result[5][291] + xnor_result[5][292] + xnor_result[5][293] + xnor_result[5][294] + xnor_result[5][295] + xnor_result[5][296] + xnor_result[5][297] + xnor_result[5][298] + xnor_result[5][299] + xnor_result[5][300] + xnor_result[5][301] + xnor_result[5][302] + xnor_result[5][303] + xnor_result[5][304] + xnor_result[5][305] + xnor_result[5][306] + xnor_result[5][307] + xnor_result[5][308] + xnor_result[5][309] + xnor_result[5][310] + xnor_result[5][311] + xnor_result[5][312] + xnor_result[5][313] + xnor_result[5][314] + xnor_result[5][315] + xnor_result[5][316] + xnor_result[5][317] + xnor_result[5][318] + xnor_result[5][319] + xnor_result[5][320] + xnor_result[5][321] + xnor_result[5][322] + xnor_result[5][323] + xnor_result[5][324] + xnor_result[5][325] + xnor_result[5][326] + xnor_result[5][327] + xnor_result[5][328] + xnor_result[5][329] + xnor_result[5][330] + xnor_result[5][331] + xnor_result[5][332] + xnor_result[5][333] + xnor_result[5][334] + xnor_result[5][335] + xnor_result[5][336] + xnor_result[5][337] + xnor_result[5][338] + xnor_result[5][339] + xnor_result[5][340] + xnor_result[5][341] + xnor_result[5][342] + xnor_result[5][343] + xnor_result[5][344] + xnor_result[5][345] + xnor_result[5][346] + xnor_result[5][347] + xnor_result[5][348] + xnor_result[5][349] + xnor_result[5][350] + xnor_result[5][351] + xnor_result[5][352] + xnor_result[5][353] + xnor_result[5][354] + xnor_result[5][355] + xnor_result[5][356] + xnor_result[5][357] + xnor_result[5][358] + xnor_result[5][359] + xnor_result[5][360] + xnor_result[5][361] + xnor_result[5][362] + xnor_result[5][363] + xnor_result[5][364] + xnor_result[5][365] + xnor_result[5][366] + xnor_result[5][367] + xnor_result[5][368] + xnor_result[5][369] + xnor_result[5][370] + xnor_result[5][371] + xnor_result[5][372] + xnor_result[5][373] + xnor_result[5][374] + xnor_result[5][375] + xnor_result[5][376] + xnor_result[5][377] + xnor_result[5][378] + xnor_result[5][379] + xnor_result[5][380] + xnor_result[5][381] + xnor_result[5][382] + xnor_result[5][383] + xnor_result[5][384] + xnor_result[5][385] + xnor_result[5][386] + xnor_result[5][387] + xnor_result[5][388] + xnor_result[5][389] + xnor_result[5][390] + xnor_result[5][391] + xnor_result[5][392] + xnor_result[5][393] + xnor_result[5][394] + xnor_result[5][395] + xnor_result[5][396] + xnor_result[5][397] + xnor_result[5][398] + xnor_result[5][399] + xnor_result[5][400] + xnor_result[5][401] + xnor_result[5][402] + xnor_result[5][403] + xnor_result[5][404] + xnor_result[5][405] + xnor_result[5][406] + xnor_result[5][407] + xnor_result[5][408] + xnor_result[5][409] + xnor_result[5][410] + xnor_result[5][411] + xnor_result[5][412] + xnor_result[5][413] + xnor_result[5][414] + xnor_result[5][415] + xnor_result[5][416] + xnor_result[5][417] + xnor_result[5][418] + xnor_result[5][419] + xnor_result[5][420] + xnor_result[5][421] + xnor_result[5][422] + xnor_result[5][423] + xnor_result[5][424] + xnor_result[5][425] + xnor_result[5][426] + xnor_result[5][427] + xnor_result[5][428] + xnor_result[5][429] + xnor_result[5][430] + xnor_result[5][431] + xnor_result[5][432] + xnor_result[5][433] + xnor_result[5][434] + xnor_result[5][435] + xnor_result[5][436] + xnor_result[5][437] + xnor_result[5][438] + xnor_result[5][439] + xnor_result[5][440] + xnor_result[5][441] + xnor_result[5][442] + xnor_result[5][443] + xnor_result[5][444] + xnor_result[5][445] + xnor_result[5][446] + xnor_result[5][447] + xnor_result[5][448] + xnor_result[5][449] + xnor_result[5][450] + xnor_result[5][451] + xnor_result[5][452] + xnor_result[5][453] + xnor_result[5][454] + xnor_result[5][455] + xnor_result[5][456] + xnor_result[5][457] + xnor_result[5][458] + xnor_result[5][459] + xnor_result[5][460] + xnor_result[5][461] + xnor_result[5][462] + xnor_result[5][463] + xnor_result[5][464] + xnor_result[5][465] + xnor_result[5][466] + xnor_result[5][467] + xnor_result[5][468] + xnor_result[5][469] + xnor_result[5][470] + xnor_result[5][471] + xnor_result[5][472] + xnor_result[5][473] + xnor_result[5][474] + xnor_result[5][475] + xnor_result[5][476] + xnor_result[5][477] + xnor_result[5][478] + xnor_result[5][479] + xnor_result[5][480] + xnor_result[5][481] + xnor_result[5][482] + xnor_result[5][483] + xnor_result[5][484] + xnor_result[5][485] + xnor_result[5][486] + xnor_result[5][487] + xnor_result[5][488] + xnor_result[5][489] + xnor_result[5][490] + xnor_result[5][491] + xnor_result[5][492] + xnor_result[5][493] + xnor_result[5][494] + xnor_result[5][495] + xnor_result[5][496] + xnor_result[5][497] + xnor_result[5][498] + xnor_result[5][499] + xnor_result[5][500] + xnor_result[5][501] + xnor_result[5][502] + xnor_result[5][503] + xnor_result[5][504] + xnor_result[5][505] + xnor_result[5][506] + xnor_result[5][507] + xnor_result[5][508] + xnor_result[5][509] + xnor_result[5][510] + xnor_result[5][511] + xnor_result[5][512] + xnor_result[5][513] + xnor_result[5][514] + xnor_result[5][515] + xnor_result[5][516] + xnor_result[5][517] + xnor_result[5][518] + xnor_result[5][519] + xnor_result[5][520] + xnor_result[5][521] + xnor_result[5][522] + xnor_result[5][523] + xnor_result[5][524] + xnor_result[5][525] + xnor_result[5][526] + xnor_result[5][527] + xnor_result[5][528] + xnor_result[5][529] + xnor_result[5][530] + xnor_result[5][531] + xnor_result[5][532] + xnor_result[5][533] + xnor_result[5][534] + xnor_result[5][535] + xnor_result[5][536] + xnor_result[5][537] + xnor_result[5][538] + xnor_result[5][539] + xnor_result[5][540] + xnor_result[5][541] + xnor_result[5][542] + xnor_result[5][543] + xnor_result[5][544] + xnor_result[5][545] + xnor_result[5][546] + xnor_result[5][547] + xnor_result[5][548] + xnor_result[5][549] + xnor_result[5][550] + xnor_result[5][551] + xnor_result[5][552] + xnor_result[5][553] + xnor_result[5][554] + xnor_result[5][555] + xnor_result[5][556] + xnor_result[5][557] + xnor_result[5][558] + xnor_result[5][559] + xnor_result[5][560] + xnor_result[5][561] + xnor_result[5][562] + xnor_result[5][563] + xnor_result[5][564] + xnor_result[5][565] + xnor_result[5][566] + xnor_result[5][567] + xnor_result[5][568] + xnor_result[5][569] + xnor_result[5][570] + xnor_result[5][571] + xnor_result[5][572] + xnor_result[5][573] + xnor_result[5][574] + xnor_result[5][575] + xnor_result[5][576] + xnor_result[5][577] + xnor_result[5][578] + xnor_result[5][579] + xnor_result[5][580] + xnor_result[5][581] + xnor_result[5][582] + xnor_result[5][583] + xnor_result[5][584] + xnor_result[5][585] + xnor_result[5][586] + xnor_result[5][587] + xnor_result[5][588] + xnor_result[5][589] + xnor_result[5][590] + xnor_result[5][591] + xnor_result[5][592] + xnor_result[5][593] + xnor_result[5][594] + xnor_result[5][595] + xnor_result[5][596] + xnor_result[5][597] + xnor_result[5][598] + xnor_result[5][599] + xnor_result[5][600] + xnor_result[5][601] + xnor_result[5][602] + xnor_result[5][603] + xnor_result[5][604] + xnor_result[5][605] + xnor_result[5][606] + xnor_result[5][607] + xnor_result[5][608] + xnor_result[5][609] + xnor_result[5][610] + xnor_result[5][611] + xnor_result[5][612] + xnor_result[5][613] + xnor_result[5][614] + xnor_result[5][615] + xnor_result[5][616] + xnor_result[5][617] + xnor_result[5][618] + xnor_result[5][619] + xnor_result[5][620] + xnor_result[5][621] + xnor_result[5][622] + xnor_result[5][623] + xnor_result[5][624] + xnor_result[5][625] + xnor_result[5][626] + xnor_result[5][627] + xnor_result[5][628] + xnor_result[5][629] + xnor_result[5][630] + xnor_result[5][631] + xnor_result[5][632] + xnor_result[5][633] + xnor_result[5][634] + xnor_result[5][635] + xnor_result[5][636] + xnor_result[5][637] + xnor_result[5][638] + xnor_result[5][639] + xnor_result[5][640] + xnor_result[5][641] + xnor_result[5][642] + xnor_result[5][643] + xnor_result[5][644] + xnor_result[5][645] + xnor_result[5][646] + xnor_result[5][647] + xnor_result[5][648] + xnor_result[5][649] + xnor_result[5][650] + xnor_result[5][651] + xnor_result[5][652] + xnor_result[5][653] + xnor_result[5][654] + xnor_result[5][655] + xnor_result[5][656] + xnor_result[5][657] + xnor_result[5][658] + xnor_result[5][659] + xnor_result[5][660] + xnor_result[5][661] + xnor_result[5][662] + xnor_result[5][663] + xnor_result[5][664] + xnor_result[5][665] + xnor_result[5][666] + xnor_result[5][667] + xnor_result[5][668] + xnor_result[5][669] + xnor_result[5][670] + xnor_result[5][671] + xnor_result[5][672] + xnor_result[5][673] + xnor_result[5][674] + xnor_result[5][675] + xnor_result[5][676] + xnor_result[5][677] + xnor_result[5][678] + xnor_result[5][679] + xnor_result[5][680] + xnor_result[5][681] + xnor_result[5][682] + xnor_result[5][683] + xnor_result[5][684] + xnor_result[5][685] + xnor_result[5][686] + xnor_result[5][687] + xnor_result[5][688] + xnor_result[5][689] + xnor_result[5][690] + xnor_result[5][691] + xnor_result[5][692] + xnor_result[5][693] + xnor_result[5][694] + xnor_result[5][695] + xnor_result[5][696] + xnor_result[5][697] + xnor_result[5][698] + xnor_result[5][699] + xnor_result[5][700] + xnor_result[5][701] + xnor_result[5][702] + xnor_result[5][703] + xnor_result[5][704] + xnor_result[5][705] + xnor_result[5][706] + xnor_result[5][707] + xnor_result[5][708] + xnor_result[5][709] + xnor_result[5][710] + xnor_result[5][711] + xnor_result[5][712] + xnor_result[5][713] + xnor_result[5][714] + xnor_result[5][715] + xnor_result[5][716] + xnor_result[5][717] + xnor_result[5][718] + xnor_result[5][719] + xnor_result[5][720] + xnor_result[5][721] + xnor_result[5][722] + xnor_result[5][723] + xnor_result[5][724] + xnor_result[5][725] + xnor_result[5][726] + xnor_result[5][727] + xnor_result[5][728] + xnor_result[5][729] + xnor_result[5][730] + xnor_result[5][731] + xnor_result[5][732] + xnor_result[5][733] + xnor_result[5][734] + xnor_result[5][735] + xnor_result[5][736] + xnor_result[5][737] + xnor_result[5][738] + xnor_result[5][739] + xnor_result[5][740] + xnor_result[5][741] + xnor_result[5][742] + xnor_result[5][743] + xnor_result[5][744] + xnor_result[5][745] + xnor_result[5][746] + xnor_result[5][747] + xnor_result[5][748] + xnor_result[5][749] + xnor_result[5][750] + xnor_result[5][751] + xnor_result[5][752] + xnor_result[5][753] + xnor_result[5][754] + xnor_result[5][755] + xnor_result[5][756] + xnor_result[5][757] + xnor_result[5][758] + xnor_result[5][759] + xnor_result[5][760] + xnor_result[5][761] + xnor_result[5][762] + xnor_result[5][763] + xnor_result[5][764] + xnor_result[5][765] + xnor_result[5][766] + xnor_result[5][767] + xnor_result[5][768] + xnor_result[5][769] + xnor_result[5][770] + xnor_result[5][771] + xnor_result[5][772] + xnor_result[5][773] + xnor_result[5][774] + xnor_result[5][775] + xnor_result[5][776] + xnor_result[5][777] + xnor_result[5][778] + xnor_result[5][779] + xnor_result[5][780] + xnor_result[5][781] + xnor_result[5][782] + xnor_result[5][783] + xnor_result[5][784] + xnor_result[5][785] + xnor_result[5][786] + xnor_result[5][787] + xnor_result[5][788] + xnor_result[5][789] + xnor_result[5][790] + xnor_result[5][791] + xnor_result[5][792] + xnor_result[5][793] + xnor_result[5][794] + xnor_result[5][795] + xnor_result[5][796] + xnor_result[5][797] + xnor_result[5][798] + xnor_result[5][799] + xnor_result[5][800] + xnor_result[5][801] + xnor_result[5][802] + xnor_result[5][803] + xnor_result[5][804] + xnor_result[5][805] + xnor_result[5][806] + xnor_result[5][807] + xnor_result[5][808] + xnor_result[5][809] + xnor_result[5][810] + xnor_result[5][811] + xnor_result[5][812] + xnor_result[5][813] + xnor_result[5][814] + xnor_result[5][815] + xnor_result[5][816] + xnor_result[5][817] + xnor_result[5][818] + xnor_result[5][819] + xnor_result[5][820] + xnor_result[5][821] + xnor_result[5][822] + xnor_result[5][823] + xnor_result[5][824] + xnor_result[5][825] + xnor_result[5][826] + xnor_result[5][827] + xnor_result[5][828] + xnor_result[5][829] + xnor_result[5][830] + xnor_result[5][831] + xnor_result[5][832] + xnor_result[5][833] + xnor_result[5][834] + xnor_result[5][835] + xnor_result[5][836] + xnor_result[5][837] + xnor_result[5][838] + xnor_result[5][839] + xnor_result[5][840] + xnor_result[5][841] + xnor_result[5][842] + xnor_result[5][843] + xnor_result[5][844] + xnor_result[5][845] + xnor_result[5][846] + xnor_result[5][847] + xnor_result[5][848] + xnor_result[5][849] + xnor_result[5][850] + xnor_result[5][851] + xnor_result[5][852] + xnor_result[5][853] + xnor_result[5][854] + xnor_result[5][855] + xnor_result[5][856] + xnor_result[5][857] + xnor_result[5][858] + xnor_result[5][859] + xnor_result[5][860] + xnor_result[5][861] + xnor_result[5][862] + xnor_result[5][863] + xnor_result[5][864] + xnor_result[5][865] + xnor_result[5][866] + xnor_result[5][867] + xnor_result[5][868] + xnor_result[5][869] + xnor_result[5][870] + xnor_result[5][871] + xnor_result[5][872] + xnor_result[5][873] + xnor_result[5][874] + xnor_result[5][875] + xnor_result[5][876] + xnor_result[5][877] + xnor_result[5][878] + xnor_result[5][879] + xnor_result[5][880] + xnor_result[5][881] + xnor_result[5][882] + xnor_result[5][883] + xnor_result[5][884] + xnor_result[5][885] + xnor_result[5][886] + xnor_result[5][887] + xnor_result[5][888] + xnor_result[5][889] + xnor_result[5][890] + xnor_result[5][891] + xnor_result[5][892] + xnor_result[5][893] + xnor_result[5][894] + xnor_result[5][895] + xnor_result[5][896] + xnor_result[5][897] + xnor_result[5][898] + xnor_result[5][899] + xnor_result[5][900] + xnor_result[5][901] + xnor_result[5][902] + xnor_result[5][903] + xnor_result[5][904] + xnor_result[5][905] + xnor_result[5][906] + xnor_result[5][907] + xnor_result[5][908] + xnor_result[5][909] + xnor_result[5][910] + xnor_result[5][911] + xnor_result[5][912] + xnor_result[5][913] + xnor_result[5][914] + xnor_result[5][915] + xnor_result[5][916] + xnor_result[5][917] + xnor_result[5][918] + xnor_result[5][919] + xnor_result[5][920] + xnor_result[5][921] + xnor_result[5][922] + xnor_result[5][923] + xnor_result[5][924] + xnor_result[5][925] + xnor_result[5][926] + xnor_result[5][927] + xnor_result[5][928] + xnor_result[5][929] + xnor_result[5][930] + xnor_result[5][931] + xnor_result[5][932] + xnor_result[5][933] + xnor_result[5][934] + xnor_result[5][935] + xnor_result[5][936] + xnor_result[5][937] + xnor_result[5][938] + xnor_result[5][939] + xnor_result[5][940] + xnor_result[5][941] + xnor_result[5][942] + xnor_result[5][943] + xnor_result[5][944] + xnor_result[5][945] + xnor_result[5][946] + xnor_result[5][947] + xnor_result[5][948] + xnor_result[5][949] + xnor_result[5][950] + xnor_result[5][951] + xnor_result[5][952] + xnor_result[5][953] + xnor_result[5][954] + xnor_result[5][955] + xnor_result[5][956] + xnor_result[5][957] + xnor_result[5][958] + xnor_result[5][959] ;
assign accumulation_result[6] = xnor_result[6][0] + xnor_result[6][1] + xnor_result[6][2] + xnor_result[6][3] + xnor_result[6][4] + xnor_result[6][5] + xnor_result[6][6] + xnor_result[6][7] + xnor_result[6][8] + xnor_result[6][9] + xnor_result[6][10] + xnor_result[6][11] + xnor_result[6][12] + xnor_result[6][13] + xnor_result[6][14] + xnor_result[6][15] + xnor_result[6][16] + xnor_result[6][17] + xnor_result[6][18] + xnor_result[6][19] + xnor_result[6][20] + xnor_result[6][21] + xnor_result[6][22] + xnor_result[6][23] + xnor_result[6][24] + xnor_result[6][25] + xnor_result[6][26] + xnor_result[6][27] + xnor_result[6][28] + xnor_result[6][29] + xnor_result[6][30] + xnor_result[6][31] + xnor_result[6][32] + xnor_result[6][33] + xnor_result[6][34] + xnor_result[6][35] + xnor_result[6][36] + xnor_result[6][37] + xnor_result[6][38] + xnor_result[6][39] + xnor_result[6][40] + xnor_result[6][41] + xnor_result[6][42] + xnor_result[6][43] + xnor_result[6][44] + xnor_result[6][45] + xnor_result[6][46] + xnor_result[6][47] + xnor_result[6][48] + xnor_result[6][49] + xnor_result[6][50] + xnor_result[6][51] + xnor_result[6][52] + xnor_result[6][53] + xnor_result[6][54] + xnor_result[6][55] + xnor_result[6][56] + xnor_result[6][57] + xnor_result[6][58] + xnor_result[6][59] + xnor_result[6][60] + xnor_result[6][61] + xnor_result[6][62] + xnor_result[6][63] + xnor_result[6][64] + xnor_result[6][65] + xnor_result[6][66] + xnor_result[6][67] + xnor_result[6][68] + xnor_result[6][69] + xnor_result[6][70] + xnor_result[6][71] + xnor_result[6][72] + xnor_result[6][73] + xnor_result[6][74] + xnor_result[6][75] + xnor_result[6][76] + xnor_result[6][77] + xnor_result[6][78] + xnor_result[6][79] + xnor_result[6][80] + xnor_result[6][81] + xnor_result[6][82] + xnor_result[6][83] + xnor_result[6][84] + xnor_result[6][85] + xnor_result[6][86] + xnor_result[6][87] + xnor_result[6][88] + xnor_result[6][89] + xnor_result[6][90] + xnor_result[6][91] + xnor_result[6][92] + xnor_result[6][93] + xnor_result[6][94] + xnor_result[6][95] + xnor_result[6][96] + xnor_result[6][97] + xnor_result[6][98] + xnor_result[6][99] + xnor_result[6][100] + xnor_result[6][101] + xnor_result[6][102] + xnor_result[6][103] + xnor_result[6][104] + xnor_result[6][105] + xnor_result[6][106] + xnor_result[6][107] + xnor_result[6][108] + xnor_result[6][109] + xnor_result[6][110] + xnor_result[6][111] + xnor_result[6][112] + xnor_result[6][113] + xnor_result[6][114] + xnor_result[6][115] + xnor_result[6][116] + xnor_result[6][117] + xnor_result[6][118] + xnor_result[6][119] + xnor_result[6][120] + xnor_result[6][121] + xnor_result[6][122] + xnor_result[6][123] + xnor_result[6][124] + xnor_result[6][125] + xnor_result[6][126] + xnor_result[6][127] + xnor_result[6][128] + xnor_result[6][129] + xnor_result[6][130] + xnor_result[6][131] + xnor_result[6][132] + xnor_result[6][133] + xnor_result[6][134] + xnor_result[6][135] + xnor_result[6][136] + xnor_result[6][137] + xnor_result[6][138] + xnor_result[6][139] + xnor_result[6][140] + xnor_result[6][141] + xnor_result[6][142] + xnor_result[6][143] + xnor_result[6][144] + xnor_result[6][145] + xnor_result[6][146] + xnor_result[6][147] + xnor_result[6][148] + xnor_result[6][149] + xnor_result[6][150] + xnor_result[6][151] + xnor_result[6][152] + xnor_result[6][153] + xnor_result[6][154] + xnor_result[6][155] + xnor_result[6][156] + xnor_result[6][157] + xnor_result[6][158] + xnor_result[6][159] + xnor_result[6][160] + xnor_result[6][161] + xnor_result[6][162] + xnor_result[6][163] + xnor_result[6][164] + xnor_result[6][165] + xnor_result[6][166] + xnor_result[6][167] + xnor_result[6][168] + xnor_result[6][169] + xnor_result[6][170] + xnor_result[6][171] + xnor_result[6][172] + xnor_result[6][173] + xnor_result[6][174] + xnor_result[6][175] + xnor_result[6][176] + xnor_result[6][177] + xnor_result[6][178] + xnor_result[6][179] + xnor_result[6][180] + xnor_result[6][181] + xnor_result[6][182] + xnor_result[6][183] + xnor_result[6][184] + xnor_result[6][185] + xnor_result[6][186] + xnor_result[6][187] + xnor_result[6][188] + xnor_result[6][189] + xnor_result[6][190] + xnor_result[6][191] + xnor_result[6][192] + xnor_result[6][193] + xnor_result[6][194] + xnor_result[6][195] + xnor_result[6][196] + xnor_result[6][197] + xnor_result[6][198] + xnor_result[6][199] + xnor_result[6][200] + xnor_result[6][201] + xnor_result[6][202] + xnor_result[6][203] + xnor_result[6][204] + xnor_result[6][205] + xnor_result[6][206] + xnor_result[6][207] + xnor_result[6][208] + xnor_result[6][209] + xnor_result[6][210] + xnor_result[6][211] + xnor_result[6][212] + xnor_result[6][213] + xnor_result[6][214] + xnor_result[6][215] + xnor_result[6][216] + xnor_result[6][217] + xnor_result[6][218] + xnor_result[6][219] + xnor_result[6][220] + xnor_result[6][221] + xnor_result[6][222] + xnor_result[6][223] + xnor_result[6][224] + xnor_result[6][225] + xnor_result[6][226] + xnor_result[6][227] + xnor_result[6][228] + xnor_result[6][229] + xnor_result[6][230] + xnor_result[6][231] + xnor_result[6][232] + xnor_result[6][233] + xnor_result[6][234] + xnor_result[6][235] + xnor_result[6][236] + xnor_result[6][237] + xnor_result[6][238] + xnor_result[6][239] + xnor_result[6][240] + xnor_result[6][241] + xnor_result[6][242] + xnor_result[6][243] + xnor_result[6][244] + xnor_result[6][245] + xnor_result[6][246] + xnor_result[6][247] + xnor_result[6][248] + xnor_result[6][249] + xnor_result[6][250] + xnor_result[6][251] + xnor_result[6][252] + xnor_result[6][253] + xnor_result[6][254] + xnor_result[6][255] + xnor_result[6][256] + xnor_result[6][257] + xnor_result[6][258] + xnor_result[6][259] + xnor_result[6][260] + xnor_result[6][261] + xnor_result[6][262] + xnor_result[6][263] + xnor_result[6][264] + xnor_result[6][265] + xnor_result[6][266] + xnor_result[6][267] + xnor_result[6][268] + xnor_result[6][269] + xnor_result[6][270] + xnor_result[6][271] + xnor_result[6][272] + xnor_result[6][273] + xnor_result[6][274] + xnor_result[6][275] + xnor_result[6][276] + xnor_result[6][277] + xnor_result[6][278] + xnor_result[6][279] + xnor_result[6][280] + xnor_result[6][281] + xnor_result[6][282] + xnor_result[6][283] + xnor_result[6][284] + xnor_result[6][285] + xnor_result[6][286] + xnor_result[6][287] + xnor_result[6][288] + xnor_result[6][289] + xnor_result[6][290] + xnor_result[6][291] + xnor_result[6][292] + xnor_result[6][293] + xnor_result[6][294] + xnor_result[6][295] + xnor_result[6][296] + xnor_result[6][297] + xnor_result[6][298] + xnor_result[6][299] + xnor_result[6][300] + xnor_result[6][301] + xnor_result[6][302] + xnor_result[6][303] + xnor_result[6][304] + xnor_result[6][305] + xnor_result[6][306] + xnor_result[6][307] + xnor_result[6][308] + xnor_result[6][309] + xnor_result[6][310] + xnor_result[6][311] + xnor_result[6][312] + xnor_result[6][313] + xnor_result[6][314] + xnor_result[6][315] + xnor_result[6][316] + xnor_result[6][317] + xnor_result[6][318] + xnor_result[6][319] + xnor_result[6][320] + xnor_result[6][321] + xnor_result[6][322] + xnor_result[6][323] + xnor_result[6][324] + xnor_result[6][325] + xnor_result[6][326] + xnor_result[6][327] + xnor_result[6][328] + xnor_result[6][329] + xnor_result[6][330] + xnor_result[6][331] + xnor_result[6][332] + xnor_result[6][333] + xnor_result[6][334] + xnor_result[6][335] + xnor_result[6][336] + xnor_result[6][337] + xnor_result[6][338] + xnor_result[6][339] + xnor_result[6][340] + xnor_result[6][341] + xnor_result[6][342] + xnor_result[6][343] + xnor_result[6][344] + xnor_result[6][345] + xnor_result[6][346] + xnor_result[6][347] + xnor_result[6][348] + xnor_result[6][349] + xnor_result[6][350] + xnor_result[6][351] + xnor_result[6][352] + xnor_result[6][353] + xnor_result[6][354] + xnor_result[6][355] + xnor_result[6][356] + xnor_result[6][357] + xnor_result[6][358] + xnor_result[6][359] + xnor_result[6][360] + xnor_result[6][361] + xnor_result[6][362] + xnor_result[6][363] + xnor_result[6][364] + xnor_result[6][365] + xnor_result[6][366] + xnor_result[6][367] + xnor_result[6][368] + xnor_result[6][369] + xnor_result[6][370] + xnor_result[6][371] + xnor_result[6][372] + xnor_result[6][373] + xnor_result[6][374] + xnor_result[6][375] + xnor_result[6][376] + xnor_result[6][377] + xnor_result[6][378] + xnor_result[6][379] + xnor_result[6][380] + xnor_result[6][381] + xnor_result[6][382] + xnor_result[6][383] + xnor_result[6][384] + xnor_result[6][385] + xnor_result[6][386] + xnor_result[6][387] + xnor_result[6][388] + xnor_result[6][389] + xnor_result[6][390] + xnor_result[6][391] + xnor_result[6][392] + xnor_result[6][393] + xnor_result[6][394] + xnor_result[6][395] + xnor_result[6][396] + xnor_result[6][397] + xnor_result[6][398] + xnor_result[6][399] + xnor_result[6][400] + xnor_result[6][401] + xnor_result[6][402] + xnor_result[6][403] + xnor_result[6][404] + xnor_result[6][405] + xnor_result[6][406] + xnor_result[6][407] + xnor_result[6][408] + xnor_result[6][409] + xnor_result[6][410] + xnor_result[6][411] + xnor_result[6][412] + xnor_result[6][413] + xnor_result[6][414] + xnor_result[6][415] + xnor_result[6][416] + xnor_result[6][417] + xnor_result[6][418] + xnor_result[6][419] + xnor_result[6][420] + xnor_result[6][421] + xnor_result[6][422] + xnor_result[6][423] + xnor_result[6][424] + xnor_result[6][425] + xnor_result[6][426] + xnor_result[6][427] + xnor_result[6][428] + xnor_result[6][429] + xnor_result[6][430] + xnor_result[6][431] + xnor_result[6][432] + xnor_result[6][433] + xnor_result[6][434] + xnor_result[6][435] + xnor_result[6][436] + xnor_result[6][437] + xnor_result[6][438] + xnor_result[6][439] + xnor_result[6][440] + xnor_result[6][441] + xnor_result[6][442] + xnor_result[6][443] + xnor_result[6][444] + xnor_result[6][445] + xnor_result[6][446] + xnor_result[6][447] + xnor_result[6][448] + xnor_result[6][449] + xnor_result[6][450] + xnor_result[6][451] + xnor_result[6][452] + xnor_result[6][453] + xnor_result[6][454] + xnor_result[6][455] + xnor_result[6][456] + xnor_result[6][457] + xnor_result[6][458] + xnor_result[6][459] + xnor_result[6][460] + xnor_result[6][461] + xnor_result[6][462] + xnor_result[6][463] + xnor_result[6][464] + xnor_result[6][465] + xnor_result[6][466] + xnor_result[6][467] + xnor_result[6][468] + xnor_result[6][469] + xnor_result[6][470] + xnor_result[6][471] + xnor_result[6][472] + xnor_result[6][473] + xnor_result[6][474] + xnor_result[6][475] + xnor_result[6][476] + xnor_result[6][477] + xnor_result[6][478] + xnor_result[6][479] + xnor_result[6][480] + xnor_result[6][481] + xnor_result[6][482] + xnor_result[6][483] + xnor_result[6][484] + xnor_result[6][485] + xnor_result[6][486] + xnor_result[6][487] + xnor_result[6][488] + xnor_result[6][489] + xnor_result[6][490] + xnor_result[6][491] + xnor_result[6][492] + xnor_result[6][493] + xnor_result[6][494] + xnor_result[6][495] + xnor_result[6][496] + xnor_result[6][497] + xnor_result[6][498] + xnor_result[6][499] + xnor_result[6][500] + xnor_result[6][501] + xnor_result[6][502] + xnor_result[6][503] + xnor_result[6][504] + xnor_result[6][505] + xnor_result[6][506] + xnor_result[6][507] + xnor_result[6][508] + xnor_result[6][509] + xnor_result[6][510] + xnor_result[6][511] + xnor_result[6][512] + xnor_result[6][513] + xnor_result[6][514] + xnor_result[6][515] + xnor_result[6][516] + xnor_result[6][517] + xnor_result[6][518] + xnor_result[6][519] + xnor_result[6][520] + xnor_result[6][521] + xnor_result[6][522] + xnor_result[6][523] + xnor_result[6][524] + xnor_result[6][525] + xnor_result[6][526] + xnor_result[6][527] + xnor_result[6][528] + xnor_result[6][529] + xnor_result[6][530] + xnor_result[6][531] + xnor_result[6][532] + xnor_result[6][533] + xnor_result[6][534] + xnor_result[6][535] + xnor_result[6][536] + xnor_result[6][537] + xnor_result[6][538] + xnor_result[6][539] + xnor_result[6][540] + xnor_result[6][541] + xnor_result[6][542] + xnor_result[6][543] + xnor_result[6][544] + xnor_result[6][545] + xnor_result[6][546] + xnor_result[6][547] + xnor_result[6][548] + xnor_result[6][549] + xnor_result[6][550] + xnor_result[6][551] + xnor_result[6][552] + xnor_result[6][553] + xnor_result[6][554] + xnor_result[6][555] + xnor_result[6][556] + xnor_result[6][557] + xnor_result[6][558] + xnor_result[6][559] + xnor_result[6][560] + xnor_result[6][561] + xnor_result[6][562] + xnor_result[6][563] + xnor_result[6][564] + xnor_result[6][565] + xnor_result[6][566] + xnor_result[6][567] + xnor_result[6][568] + xnor_result[6][569] + xnor_result[6][570] + xnor_result[6][571] + xnor_result[6][572] + xnor_result[6][573] + xnor_result[6][574] + xnor_result[6][575] + xnor_result[6][576] + xnor_result[6][577] + xnor_result[6][578] + xnor_result[6][579] + xnor_result[6][580] + xnor_result[6][581] + xnor_result[6][582] + xnor_result[6][583] + xnor_result[6][584] + xnor_result[6][585] + xnor_result[6][586] + xnor_result[6][587] + xnor_result[6][588] + xnor_result[6][589] + xnor_result[6][590] + xnor_result[6][591] + xnor_result[6][592] + xnor_result[6][593] + xnor_result[6][594] + xnor_result[6][595] + xnor_result[6][596] + xnor_result[6][597] + xnor_result[6][598] + xnor_result[6][599] + xnor_result[6][600] + xnor_result[6][601] + xnor_result[6][602] + xnor_result[6][603] + xnor_result[6][604] + xnor_result[6][605] + xnor_result[6][606] + xnor_result[6][607] + xnor_result[6][608] + xnor_result[6][609] + xnor_result[6][610] + xnor_result[6][611] + xnor_result[6][612] + xnor_result[6][613] + xnor_result[6][614] + xnor_result[6][615] + xnor_result[6][616] + xnor_result[6][617] + xnor_result[6][618] + xnor_result[6][619] + xnor_result[6][620] + xnor_result[6][621] + xnor_result[6][622] + xnor_result[6][623] + xnor_result[6][624] + xnor_result[6][625] + xnor_result[6][626] + xnor_result[6][627] + xnor_result[6][628] + xnor_result[6][629] + xnor_result[6][630] + xnor_result[6][631] + xnor_result[6][632] + xnor_result[6][633] + xnor_result[6][634] + xnor_result[6][635] + xnor_result[6][636] + xnor_result[6][637] + xnor_result[6][638] + xnor_result[6][639] + xnor_result[6][640] + xnor_result[6][641] + xnor_result[6][642] + xnor_result[6][643] + xnor_result[6][644] + xnor_result[6][645] + xnor_result[6][646] + xnor_result[6][647] + xnor_result[6][648] + xnor_result[6][649] + xnor_result[6][650] + xnor_result[6][651] + xnor_result[6][652] + xnor_result[6][653] + xnor_result[6][654] + xnor_result[6][655] + xnor_result[6][656] + xnor_result[6][657] + xnor_result[6][658] + xnor_result[6][659] + xnor_result[6][660] + xnor_result[6][661] + xnor_result[6][662] + xnor_result[6][663] + xnor_result[6][664] + xnor_result[6][665] + xnor_result[6][666] + xnor_result[6][667] + xnor_result[6][668] + xnor_result[6][669] + xnor_result[6][670] + xnor_result[6][671] + xnor_result[6][672] + xnor_result[6][673] + xnor_result[6][674] + xnor_result[6][675] + xnor_result[6][676] + xnor_result[6][677] + xnor_result[6][678] + xnor_result[6][679] + xnor_result[6][680] + xnor_result[6][681] + xnor_result[6][682] + xnor_result[6][683] + xnor_result[6][684] + xnor_result[6][685] + xnor_result[6][686] + xnor_result[6][687] + xnor_result[6][688] + xnor_result[6][689] + xnor_result[6][690] + xnor_result[6][691] + xnor_result[6][692] + xnor_result[6][693] + xnor_result[6][694] + xnor_result[6][695] + xnor_result[6][696] + xnor_result[6][697] + xnor_result[6][698] + xnor_result[6][699] + xnor_result[6][700] + xnor_result[6][701] + xnor_result[6][702] + xnor_result[6][703] + xnor_result[6][704] + xnor_result[6][705] + xnor_result[6][706] + xnor_result[6][707] + xnor_result[6][708] + xnor_result[6][709] + xnor_result[6][710] + xnor_result[6][711] + xnor_result[6][712] + xnor_result[6][713] + xnor_result[6][714] + xnor_result[6][715] + xnor_result[6][716] + xnor_result[6][717] + xnor_result[6][718] + xnor_result[6][719] + xnor_result[6][720] + xnor_result[6][721] + xnor_result[6][722] + xnor_result[6][723] + xnor_result[6][724] + xnor_result[6][725] + xnor_result[6][726] + xnor_result[6][727] + xnor_result[6][728] + xnor_result[6][729] + xnor_result[6][730] + xnor_result[6][731] + xnor_result[6][732] + xnor_result[6][733] + xnor_result[6][734] + xnor_result[6][735] + xnor_result[6][736] + xnor_result[6][737] + xnor_result[6][738] + xnor_result[6][739] + xnor_result[6][740] + xnor_result[6][741] + xnor_result[6][742] + xnor_result[6][743] + xnor_result[6][744] + xnor_result[6][745] + xnor_result[6][746] + xnor_result[6][747] + xnor_result[6][748] + xnor_result[6][749] + xnor_result[6][750] + xnor_result[6][751] + xnor_result[6][752] + xnor_result[6][753] + xnor_result[6][754] + xnor_result[6][755] + xnor_result[6][756] + xnor_result[6][757] + xnor_result[6][758] + xnor_result[6][759] + xnor_result[6][760] + xnor_result[6][761] + xnor_result[6][762] + xnor_result[6][763] + xnor_result[6][764] + xnor_result[6][765] + xnor_result[6][766] + xnor_result[6][767] + xnor_result[6][768] + xnor_result[6][769] + xnor_result[6][770] + xnor_result[6][771] + xnor_result[6][772] + xnor_result[6][773] + xnor_result[6][774] + xnor_result[6][775] + xnor_result[6][776] + xnor_result[6][777] + xnor_result[6][778] + xnor_result[6][779] + xnor_result[6][780] + xnor_result[6][781] + xnor_result[6][782] + xnor_result[6][783] + xnor_result[6][784] + xnor_result[6][785] + xnor_result[6][786] + xnor_result[6][787] + xnor_result[6][788] + xnor_result[6][789] + xnor_result[6][790] + xnor_result[6][791] + xnor_result[6][792] + xnor_result[6][793] + xnor_result[6][794] + xnor_result[6][795] + xnor_result[6][796] + xnor_result[6][797] + xnor_result[6][798] + xnor_result[6][799] + xnor_result[6][800] + xnor_result[6][801] + xnor_result[6][802] + xnor_result[6][803] + xnor_result[6][804] + xnor_result[6][805] + xnor_result[6][806] + xnor_result[6][807] + xnor_result[6][808] + xnor_result[6][809] + xnor_result[6][810] + xnor_result[6][811] + xnor_result[6][812] + xnor_result[6][813] + xnor_result[6][814] + xnor_result[6][815] + xnor_result[6][816] + xnor_result[6][817] + xnor_result[6][818] + xnor_result[6][819] + xnor_result[6][820] + xnor_result[6][821] + xnor_result[6][822] + xnor_result[6][823] + xnor_result[6][824] + xnor_result[6][825] + xnor_result[6][826] + xnor_result[6][827] + xnor_result[6][828] + xnor_result[6][829] + xnor_result[6][830] + xnor_result[6][831] + xnor_result[6][832] + xnor_result[6][833] + xnor_result[6][834] + xnor_result[6][835] + xnor_result[6][836] + xnor_result[6][837] + xnor_result[6][838] + xnor_result[6][839] + xnor_result[6][840] + xnor_result[6][841] + xnor_result[6][842] + xnor_result[6][843] + xnor_result[6][844] + xnor_result[6][845] + xnor_result[6][846] + xnor_result[6][847] + xnor_result[6][848] + xnor_result[6][849] + xnor_result[6][850] + xnor_result[6][851] + xnor_result[6][852] + xnor_result[6][853] + xnor_result[6][854] + xnor_result[6][855] + xnor_result[6][856] + xnor_result[6][857] + xnor_result[6][858] + xnor_result[6][859] + xnor_result[6][860] + xnor_result[6][861] + xnor_result[6][862] + xnor_result[6][863] + xnor_result[6][864] + xnor_result[6][865] + xnor_result[6][866] + xnor_result[6][867] + xnor_result[6][868] + xnor_result[6][869] + xnor_result[6][870] + xnor_result[6][871] + xnor_result[6][872] + xnor_result[6][873] + xnor_result[6][874] + xnor_result[6][875] + xnor_result[6][876] + xnor_result[6][877] + xnor_result[6][878] + xnor_result[6][879] + xnor_result[6][880] + xnor_result[6][881] + xnor_result[6][882] + xnor_result[6][883] + xnor_result[6][884] + xnor_result[6][885] + xnor_result[6][886] + xnor_result[6][887] + xnor_result[6][888] + xnor_result[6][889] + xnor_result[6][890] + xnor_result[6][891] + xnor_result[6][892] + xnor_result[6][893] + xnor_result[6][894] + xnor_result[6][895] + xnor_result[6][896] + xnor_result[6][897] + xnor_result[6][898] + xnor_result[6][899] + xnor_result[6][900] + xnor_result[6][901] + xnor_result[6][902] + xnor_result[6][903] + xnor_result[6][904] + xnor_result[6][905] + xnor_result[6][906] + xnor_result[6][907] + xnor_result[6][908] + xnor_result[6][909] + xnor_result[6][910] + xnor_result[6][911] + xnor_result[6][912] + xnor_result[6][913] + xnor_result[6][914] + xnor_result[6][915] + xnor_result[6][916] + xnor_result[6][917] + xnor_result[6][918] + xnor_result[6][919] + xnor_result[6][920] + xnor_result[6][921] + xnor_result[6][922] + xnor_result[6][923] + xnor_result[6][924] + xnor_result[6][925] + xnor_result[6][926] + xnor_result[6][927] + xnor_result[6][928] + xnor_result[6][929] + xnor_result[6][930] + xnor_result[6][931] + xnor_result[6][932] + xnor_result[6][933] + xnor_result[6][934] + xnor_result[6][935] + xnor_result[6][936] + xnor_result[6][937] + xnor_result[6][938] + xnor_result[6][939] + xnor_result[6][940] + xnor_result[6][941] + xnor_result[6][942] + xnor_result[6][943] + xnor_result[6][944] + xnor_result[6][945] + xnor_result[6][946] + xnor_result[6][947] + xnor_result[6][948] + xnor_result[6][949] + xnor_result[6][950] + xnor_result[6][951] + xnor_result[6][952] + xnor_result[6][953] + xnor_result[6][954] + xnor_result[6][955] + xnor_result[6][956] + xnor_result[6][957] + xnor_result[6][958] + xnor_result[6][959] ;
assign accumulation_result[7] = xnor_result[7][0] + xnor_result[7][1] + xnor_result[7][2] + xnor_result[7][3] + xnor_result[7][4] + xnor_result[7][5] + xnor_result[7][6] + xnor_result[7][7] + xnor_result[7][8] + xnor_result[7][9] + xnor_result[7][10] + xnor_result[7][11] + xnor_result[7][12] + xnor_result[7][13] + xnor_result[7][14] + xnor_result[7][15] + xnor_result[7][16] + xnor_result[7][17] + xnor_result[7][18] + xnor_result[7][19] + xnor_result[7][20] + xnor_result[7][21] + xnor_result[7][22] + xnor_result[7][23] + xnor_result[7][24] + xnor_result[7][25] + xnor_result[7][26] + xnor_result[7][27] + xnor_result[7][28] + xnor_result[7][29] + xnor_result[7][30] + xnor_result[7][31] + xnor_result[7][32] + xnor_result[7][33] + xnor_result[7][34] + xnor_result[7][35] + xnor_result[7][36] + xnor_result[7][37] + xnor_result[7][38] + xnor_result[7][39] + xnor_result[7][40] + xnor_result[7][41] + xnor_result[7][42] + xnor_result[7][43] + xnor_result[7][44] + xnor_result[7][45] + xnor_result[7][46] + xnor_result[7][47] + xnor_result[7][48] + xnor_result[7][49] + xnor_result[7][50] + xnor_result[7][51] + xnor_result[7][52] + xnor_result[7][53] + xnor_result[7][54] + xnor_result[7][55] + xnor_result[7][56] + xnor_result[7][57] + xnor_result[7][58] + xnor_result[7][59] + xnor_result[7][60] + xnor_result[7][61] + xnor_result[7][62] + xnor_result[7][63] + xnor_result[7][64] + xnor_result[7][65] + xnor_result[7][66] + xnor_result[7][67] + xnor_result[7][68] + xnor_result[7][69] + xnor_result[7][70] + xnor_result[7][71] + xnor_result[7][72] + xnor_result[7][73] + xnor_result[7][74] + xnor_result[7][75] + xnor_result[7][76] + xnor_result[7][77] + xnor_result[7][78] + xnor_result[7][79] + xnor_result[7][80] + xnor_result[7][81] + xnor_result[7][82] + xnor_result[7][83] + xnor_result[7][84] + xnor_result[7][85] + xnor_result[7][86] + xnor_result[7][87] + xnor_result[7][88] + xnor_result[7][89] + xnor_result[7][90] + xnor_result[7][91] + xnor_result[7][92] + xnor_result[7][93] + xnor_result[7][94] + xnor_result[7][95] + xnor_result[7][96] + xnor_result[7][97] + xnor_result[7][98] + xnor_result[7][99] + xnor_result[7][100] + xnor_result[7][101] + xnor_result[7][102] + xnor_result[7][103] + xnor_result[7][104] + xnor_result[7][105] + xnor_result[7][106] + xnor_result[7][107] + xnor_result[7][108] + xnor_result[7][109] + xnor_result[7][110] + xnor_result[7][111] + xnor_result[7][112] + xnor_result[7][113] + xnor_result[7][114] + xnor_result[7][115] + xnor_result[7][116] + xnor_result[7][117] + xnor_result[7][118] + xnor_result[7][119] + xnor_result[7][120] + xnor_result[7][121] + xnor_result[7][122] + xnor_result[7][123] + xnor_result[7][124] + xnor_result[7][125] + xnor_result[7][126] + xnor_result[7][127] + xnor_result[7][128] + xnor_result[7][129] + xnor_result[7][130] + xnor_result[7][131] + xnor_result[7][132] + xnor_result[7][133] + xnor_result[7][134] + xnor_result[7][135] + xnor_result[7][136] + xnor_result[7][137] + xnor_result[7][138] + xnor_result[7][139] + xnor_result[7][140] + xnor_result[7][141] + xnor_result[7][142] + xnor_result[7][143] + xnor_result[7][144] + xnor_result[7][145] + xnor_result[7][146] + xnor_result[7][147] + xnor_result[7][148] + xnor_result[7][149] + xnor_result[7][150] + xnor_result[7][151] + xnor_result[7][152] + xnor_result[7][153] + xnor_result[7][154] + xnor_result[7][155] + xnor_result[7][156] + xnor_result[7][157] + xnor_result[7][158] + xnor_result[7][159] + xnor_result[7][160] + xnor_result[7][161] + xnor_result[7][162] + xnor_result[7][163] + xnor_result[7][164] + xnor_result[7][165] + xnor_result[7][166] + xnor_result[7][167] + xnor_result[7][168] + xnor_result[7][169] + xnor_result[7][170] + xnor_result[7][171] + xnor_result[7][172] + xnor_result[7][173] + xnor_result[7][174] + xnor_result[7][175] + xnor_result[7][176] + xnor_result[7][177] + xnor_result[7][178] + xnor_result[7][179] + xnor_result[7][180] + xnor_result[7][181] + xnor_result[7][182] + xnor_result[7][183] + xnor_result[7][184] + xnor_result[7][185] + xnor_result[7][186] + xnor_result[7][187] + xnor_result[7][188] + xnor_result[7][189] + xnor_result[7][190] + xnor_result[7][191] + xnor_result[7][192] + xnor_result[7][193] + xnor_result[7][194] + xnor_result[7][195] + xnor_result[7][196] + xnor_result[7][197] + xnor_result[7][198] + xnor_result[7][199] + xnor_result[7][200] + xnor_result[7][201] + xnor_result[7][202] + xnor_result[7][203] + xnor_result[7][204] + xnor_result[7][205] + xnor_result[7][206] + xnor_result[7][207] + xnor_result[7][208] + xnor_result[7][209] + xnor_result[7][210] + xnor_result[7][211] + xnor_result[7][212] + xnor_result[7][213] + xnor_result[7][214] + xnor_result[7][215] + xnor_result[7][216] + xnor_result[7][217] + xnor_result[7][218] + xnor_result[7][219] + xnor_result[7][220] + xnor_result[7][221] + xnor_result[7][222] + xnor_result[7][223] + xnor_result[7][224] + xnor_result[7][225] + xnor_result[7][226] + xnor_result[7][227] + xnor_result[7][228] + xnor_result[7][229] + xnor_result[7][230] + xnor_result[7][231] + xnor_result[7][232] + xnor_result[7][233] + xnor_result[7][234] + xnor_result[7][235] + xnor_result[7][236] + xnor_result[7][237] + xnor_result[7][238] + xnor_result[7][239] + xnor_result[7][240] + xnor_result[7][241] + xnor_result[7][242] + xnor_result[7][243] + xnor_result[7][244] + xnor_result[7][245] + xnor_result[7][246] + xnor_result[7][247] + xnor_result[7][248] + xnor_result[7][249] + xnor_result[7][250] + xnor_result[7][251] + xnor_result[7][252] + xnor_result[7][253] + xnor_result[7][254] + xnor_result[7][255] + xnor_result[7][256] + xnor_result[7][257] + xnor_result[7][258] + xnor_result[7][259] + xnor_result[7][260] + xnor_result[7][261] + xnor_result[7][262] + xnor_result[7][263] + xnor_result[7][264] + xnor_result[7][265] + xnor_result[7][266] + xnor_result[7][267] + xnor_result[7][268] + xnor_result[7][269] + xnor_result[7][270] + xnor_result[7][271] + xnor_result[7][272] + xnor_result[7][273] + xnor_result[7][274] + xnor_result[7][275] + xnor_result[7][276] + xnor_result[7][277] + xnor_result[7][278] + xnor_result[7][279] + xnor_result[7][280] + xnor_result[7][281] + xnor_result[7][282] + xnor_result[7][283] + xnor_result[7][284] + xnor_result[7][285] + xnor_result[7][286] + xnor_result[7][287] + xnor_result[7][288] + xnor_result[7][289] + xnor_result[7][290] + xnor_result[7][291] + xnor_result[7][292] + xnor_result[7][293] + xnor_result[7][294] + xnor_result[7][295] + xnor_result[7][296] + xnor_result[7][297] + xnor_result[7][298] + xnor_result[7][299] + xnor_result[7][300] + xnor_result[7][301] + xnor_result[7][302] + xnor_result[7][303] + xnor_result[7][304] + xnor_result[7][305] + xnor_result[7][306] + xnor_result[7][307] + xnor_result[7][308] + xnor_result[7][309] + xnor_result[7][310] + xnor_result[7][311] + xnor_result[7][312] + xnor_result[7][313] + xnor_result[7][314] + xnor_result[7][315] + xnor_result[7][316] + xnor_result[7][317] + xnor_result[7][318] + xnor_result[7][319] + xnor_result[7][320] + xnor_result[7][321] + xnor_result[7][322] + xnor_result[7][323] + xnor_result[7][324] + xnor_result[7][325] + xnor_result[7][326] + xnor_result[7][327] + xnor_result[7][328] + xnor_result[7][329] + xnor_result[7][330] + xnor_result[7][331] + xnor_result[7][332] + xnor_result[7][333] + xnor_result[7][334] + xnor_result[7][335] + xnor_result[7][336] + xnor_result[7][337] + xnor_result[7][338] + xnor_result[7][339] + xnor_result[7][340] + xnor_result[7][341] + xnor_result[7][342] + xnor_result[7][343] + xnor_result[7][344] + xnor_result[7][345] + xnor_result[7][346] + xnor_result[7][347] + xnor_result[7][348] + xnor_result[7][349] + xnor_result[7][350] + xnor_result[7][351] + xnor_result[7][352] + xnor_result[7][353] + xnor_result[7][354] + xnor_result[7][355] + xnor_result[7][356] + xnor_result[7][357] + xnor_result[7][358] + xnor_result[7][359] + xnor_result[7][360] + xnor_result[7][361] + xnor_result[7][362] + xnor_result[7][363] + xnor_result[7][364] + xnor_result[7][365] + xnor_result[7][366] + xnor_result[7][367] + xnor_result[7][368] + xnor_result[7][369] + xnor_result[7][370] + xnor_result[7][371] + xnor_result[7][372] + xnor_result[7][373] + xnor_result[7][374] + xnor_result[7][375] + xnor_result[7][376] + xnor_result[7][377] + xnor_result[7][378] + xnor_result[7][379] + xnor_result[7][380] + xnor_result[7][381] + xnor_result[7][382] + xnor_result[7][383] + xnor_result[7][384] + xnor_result[7][385] + xnor_result[7][386] + xnor_result[7][387] + xnor_result[7][388] + xnor_result[7][389] + xnor_result[7][390] + xnor_result[7][391] + xnor_result[7][392] + xnor_result[7][393] + xnor_result[7][394] + xnor_result[7][395] + xnor_result[7][396] + xnor_result[7][397] + xnor_result[7][398] + xnor_result[7][399] + xnor_result[7][400] + xnor_result[7][401] + xnor_result[7][402] + xnor_result[7][403] + xnor_result[7][404] + xnor_result[7][405] + xnor_result[7][406] + xnor_result[7][407] + xnor_result[7][408] + xnor_result[7][409] + xnor_result[7][410] + xnor_result[7][411] + xnor_result[7][412] + xnor_result[7][413] + xnor_result[7][414] + xnor_result[7][415] + xnor_result[7][416] + xnor_result[7][417] + xnor_result[7][418] + xnor_result[7][419] + xnor_result[7][420] + xnor_result[7][421] + xnor_result[7][422] + xnor_result[7][423] + xnor_result[7][424] + xnor_result[7][425] + xnor_result[7][426] + xnor_result[7][427] + xnor_result[7][428] + xnor_result[7][429] + xnor_result[7][430] + xnor_result[7][431] + xnor_result[7][432] + xnor_result[7][433] + xnor_result[7][434] + xnor_result[7][435] + xnor_result[7][436] + xnor_result[7][437] + xnor_result[7][438] + xnor_result[7][439] + xnor_result[7][440] + xnor_result[7][441] + xnor_result[7][442] + xnor_result[7][443] + xnor_result[7][444] + xnor_result[7][445] + xnor_result[7][446] + xnor_result[7][447] + xnor_result[7][448] + xnor_result[7][449] + xnor_result[7][450] + xnor_result[7][451] + xnor_result[7][452] + xnor_result[7][453] + xnor_result[7][454] + xnor_result[7][455] + xnor_result[7][456] + xnor_result[7][457] + xnor_result[7][458] + xnor_result[7][459] + xnor_result[7][460] + xnor_result[7][461] + xnor_result[7][462] + xnor_result[7][463] + xnor_result[7][464] + xnor_result[7][465] + xnor_result[7][466] + xnor_result[7][467] + xnor_result[7][468] + xnor_result[7][469] + xnor_result[7][470] + xnor_result[7][471] + xnor_result[7][472] + xnor_result[7][473] + xnor_result[7][474] + xnor_result[7][475] + xnor_result[7][476] + xnor_result[7][477] + xnor_result[7][478] + xnor_result[7][479] + xnor_result[7][480] + xnor_result[7][481] + xnor_result[7][482] + xnor_result[7][483] + xnor_result[7][484] + xnor_result[7][485] + xnor_result[7][486] + xnor_result[7][487] + xnor_result[7][488] + xnor_result[7][489] + xnor_result[7][490] + xnor_result[7][491] + xnor_result[7][492] + xnor_result[7][493] + xnor_result[7][494] + xnor_result[7][495] + xnor_result[7][496] + xnor_result[7][497] + xnor_result[7][498] + xnor_result[7][499] + xnor_result[7][500] + xnor_result[7][501] + xnor_result[7][502] + xnor_result[7][503] + xnor_result[7][504] + xnor_result[7][505] + xnor_result[7][506] + xnor_result[7][507] + xnor_result[7][508] + xnor_result[7][509] + xnor_result[7][510] + xnor_result[7][511] + xnor_result[7][512] + xnor_result[7][513] + xnor_result[7][514] + xnor_result[7][515] + xnor_result[7][516] + xnor_result[7][517] + xnor_result[7][518] + xnor_result[7][519] + xnor_result[7][520] + xnor_result[7][521] + xnor_result[7][522] + xnor_result[7][523] + xnor_result[7][524] + xnor_result[7][525] + xnor_result[7][526] + xnor_result[7][527] + xnor_result[7][528] + xnor_result[7][529] + xnor_result[7][530] + xnor_result[7][531] + xnor_result[7][532] + xnor_result[7][533] + xnor_result[7][534] + xnor_result[7][535] + xnor_result[7][536] + xnor_result[7][537] + xnor_result[7][538] + xnor_result[7][539] + xnor_result[7][540] + xnor_result[7][541] + xnor_result[7][542] + xnor_result[7][543] + xnor_result[7][544] + xnor_result[7][545] + xnor_result[7][546] + xnor_result[7][547] + xnor_result[7][548] + xnor_result[7][549] + xnor_result[7][550] + xnor_result[7][551] + xnor_result[7][552] + xnor_result[7][553] + xnor_result[7][554] + xnor_result[7][555] + xnor_result[7][556] + xnor_result[7][557] + xnor_result[7][558] + xnor_result[7][559] + xnor_result[7][560] + xnor_result[7][561] + xnor_result[7][562] + xnor_result[7][563] + xnor_result[7][564] + xnor_result[7][565] + xnor_result[7][566] + xnor_result[7][567] + xnor_result[7][568] + xnor_result[7][569] + xnor_result[7][570] + xnor_result[7][571] + xnor_result[7][572] + xnor_result[7][573] + xnor_result[7][574] + xnor_result[7][575] + xnor_result[7][576] + xnor_result[7][577] + xnor_result[7][578] + xnor_result[7][579] + xnor_result[7][580] + xnor_result[7][581] + xnor_result[7][582] + xnor_result[7][583] + xnor_result[7][584] + xnor_result[7][585] + xnor_result[7][586] + xnor_result[7][587] + xnor_result[7][588] + xnor_result[7][589] + xnor_result[7][590] + xnor_result[7][591] + xnor_result[7][592] + xnor_result[7][593] + xnor_result[7][594] + xnor_result[7][595] + xnor_result[7][596] + xnor_result[7][597] + xnor_result[7][598] + xnor_result[7][599] + xnor_result[7][600] + xnor_result[7][601] + xnor_result[7][602] + xnor_result[7][603] + xnor_result[7][604] + xnor_result[7][605] + xnor_result[7][606] + xnor_result[7][607] + xnor_result[7][608] + xnor_result[7][609] + xnor_result[7][610] + xnor_result[7][611] + xnor_result[7][612] + xnor_result[7][613] + xnor_result[7][614] + xnor_result[7][615] + xnor_result[7][616] + xnor_result[7][617] + xnor_result[7][618] + xnor_result[7][619] + xnor_result[7][620] + xnor_result[7][621] + xnor_result[7][622] + xnor_result[7][623] + xnor_result[7][624] + xnor_result[7][625] + xnor_result[7][626] + xnor_result[7][627] + xnor_result[7][628] + xnor_result[7][629] + xnor_result[7][630] + xnor_result[7][631] + xnor_result[7][632] + xnor_result[7][633] + xnor_result[7][634] + xnor_result[7][635] + xnor_result[7][636] + xnor_result[7][637] + xnor_result[7][638] + xnor_result[7][639] + xnor_result[7][640] + xnor_result[7][641] + xnor_result[7][642] + xnor_result[7][643] + xnor_result[7][644] + xnor_result[7][645] + xnor_result[7][646] + xnor_result[7][647] + xnor_result[7][648] + xnor_result[7][649] + xnor_result[7][650] + xnor_result[7][651] + xnor_result[7][652] + xnor_result[7][653] + xnor_result[7][654] + xnor_result[7][655] + xnor_result[7][656] + xnor_result[7][657] + xnor_result[7][658] + xnor_result[7][659] + xnor_result[7][660] + xnor_result[7][661] + xnor_result[7][662] + xnor_result[7][663] + xnor_result[7][664] + xnor_result[7][665] + xnor_result[7][666] + xnor_result[7][667] + xnor_result[7][668] + xnor_result[7][669] + xnor_result[7][670] + xnor_result[7][671] + xnor_result[7][672] + xnor_result[7][673] + xnor_result[7][674] + xnor_result[7][675] + xnor_result[7][676] + xnor_result[7][677] + xnor_result[7][678] + xnor_result[7][679] + xnor_result[7][680] + xnor_result[7][681] + xnor_result[7][682] + xnor_result[7][683] + xnor_result[7][684] + xnor_result[7][685] + xnor_result[7][686] + xnor_result[7][687] + xnor_result[7][688] + xnor_result[7][689] + xnor_result[7][690] + xnor_result[7][691] + xnor_result[7][692] + xnor_result[7][693] + xnor_result[7][694] + xnor_result[7][695] + xnor_result[7][696] + xnor_result[7][697] + xnor_result[7][698] + xnor_result[7][699] + xnor_result[7][700] + xnor_result[7][701] + xnor_result[7][702] + xnor_result[7][703] + xnor_result[7][704] + xnor_result[7][705] + xnor_result[7][706] + xnor_result[7][707] + xnor_result[7][708] + xnor_result[7][709] + xnor_result[7][710] + xnor_result[7][711] + xnor_result[7][712] + xnor_result[7][713] + xnor_result[7][714] + xnor_result[7][715] + xnor_result[7][716] + xnor_result[7][717] + xnor_result[7][718] + xnor_result[7][719] + xnor_result[7][720] + xnor_result[7][721] + xnor_result[7][722] + xnor_result[7][723] + xnor_result[7][724] + xnor_result[7][725] + xnor_result[7][726] + xnor_result[7][727] + xnor_result[7][728] + xnor_result[7][729] + xnor_result[7][730] + xnor_result[7][731] + xnor_result[7][732] + xnor_result[7][733] + xnor_result[7][734] + xnor_result[7][735] + xnor_result[7][736] + xnor_result[7][737] + xnor_result[7][738] + xnor_result[7][739] + xnor_result[7][740] + xnor_result[7][741] + xnor_result[7][742] + xnor_result[7][743] + xnor_result[7][744] + xnor_result[7][745] + xnor_result[7][746] + xnor_result[7][747] + xnor_result[7][748] + xnor_result[7][749] + xnor_result[7][750] + xnor_result[7][751] + xnor_result[7][752] + xnor_result[7][753] + xnor_result[7][754] + xnor_result[7][755] + xnor_result[7][756] + xnor_result[7][757] + xnor_result[7][758] + xnor_result[7][759] + xnor_result[7][760] + xnor_result[7][761] + xnor_result[7][762] + xnor_result[7][763] + xnor_result[7][764] + xnor_result[7][765] + xnor_result[7][766] + xnor_result[7][767] + xnor_result[7][768] + xnor_result[7][769] + xnor_result[7][770] + xnor_result[7][771] + xnor_result[7][772] + xnor_result[7][773] + xnor_result[7][774] + xnor_result[7][775] + xnor_result[7][776] + xnor_result[7][777] + xnor_result[7][778] + xnor_result[7][779] + xnor_result[7][780] + xnor_result[7][781] + xnor_result[7][782] + xnor_result[7][783] + xnor_result[7][784] + xnor_result[7][785] + xnor_result[7][786] + xnor_result[7][787] + xnor_result[7][788] + xnor_result[7][789] + xnor_result[7][790] + xnor_result[7][791] + xnor_result[7][792] + xnor_result[7][793] + xnor_result[7][794] + xnor_result[7][795] + xnor_result[7][796] + xnor_result[7][797] + xnor_result[7][798] + xnor_result[7][799] + xnor_result[7][800] + xnor_result[7][801] + xnor_result[7][802] + xnor_result[7][803] + xnor_result[7][804] + xnor_result[7][805] + xnor_result[7][806] + xnor_result[7][807] + xnor_result[7][808] + xnor_result[7][809] + xnor_result[7][810] + xnor_result[7][811] + xnor_result[7][812] + xnor_result[7][813] + xnor_result[7][814] + xnor_result[7][815] + xnor_result[7][816] + xnor_result[7][817] + xnor_result[7][818] + xnor_result[7][819] + xnor_result[7][820] + xnor_result[7][821] + xnor_result[7][822] + xnor_result[7][823] + xnor_result[7][824] + xnor_result[7][825] + xnor_result[7][826] + xnor_result[7][827] + xnor_result[7][828] + xnor_result[7][829] + xnor_result[7][830] + xnor_result[7][831] + xnor_result[7][832] + xnor_result[7][833] + xnor_result[7][834] + xnor_result[7][835] + xnor_result[7][836] + xnor_result[7][837] + xnor_result[7][838] + xnor_result[7][839] + xnor_result[7][840] + xnor_result[7][841] + xnor_result[7][842] + xnor_result[7][843] + xnor_result[7][844] + xnor_result[7][845] + xnor_result[7][846] + xnor_result[7][847] + xnor_result[7][848] + xnor_result[7][849] + xnor_result[7][850] + xnor_result[7][851] + xnor_result[7][852] + xnor_result[7][853] + xnor_result[7][854] + xnor_result[7][855] + xnor_result[7][856] + xnor_result[7][857] + xnor_result[7][858] + xnor_result[7][859] + xnor_result[7][860] + xnor_result[7][861] + xnor_result[7][862] + xnor_result[7][863] + xnor_result[7][864] + xnor_result[7][865] + xnor_result[7][866] + xnor_result[7][867] + xnor_result[7][868] + xnor_result[7][869] + xnor_result[7][870] + xnor_result[7][871] + xnor_result[7][872] + xnor_result[7][873] + xnor_result[7][874] + xnor_result[7][875] + xnor_result[7][876] + xnor_result[7][877] + xnor_result[7][878] + xnor_result[7][879] + xnor_result[7][880] + xnor_result[7][881] + xnor_result[7][882] + xnor_result[7][883] + xnor_result[7][884] + xnor_result[7][885] + xnor_result[7][886] + xnor_result[7][887] + xnor_result[7][888] + xnor_result[7][889] + xnor_result[7][890] + xnor_result[7][891] + xnor_result[7][892] + xnor_result[7][893] + xnor_result[7][894] + xnor_result[7][895] + xnor_result[7][896] + xnor_result[7][897] + xnor_result[7][898] + xnor_result[7][899] + xnor_result[7][900] + xnor_result[7][901] + xnor_result[7][902] + xnor_result[7][903] + xnor_result[7][904] + xnor_result[7][905] + xnor_result[7][906] + xnor_result[7][907] + xnor_result[7][908] + xnor_result[7][909] + xnor_result[7][910] + xnor_result[7][911] + xnor_result[7][912] + xnor_result[7][913] + xnor_result[7][914] + xnor_result[7][915] + xnor_result[7][916] + xnor_result[7][917] + xnor_result[7][918] + xnor_result[7][919] + xnor_result[7][920] + xnor_result[7][921] + xnor_result[7][922] + xnor_result[7][923] + xnor_result[7][924] + xnor_result[7][925] + xnor_result[7][926] + xnor_result[7][927] + xnor_result[7][928] + xnor_result[7][929] + xnor_result[7][930] + xnor_result[7][931] + xnor_result[7][932] + xnor_result[7][933] + xnor_result[7][934] + xnor_result[7][935] + xnor_result[7][936] + xnor_result[7][937] + xnor_result[7][938] + xnor_result[7][939] + xnor_result[7][940] + xnor_result[7][941] + xnor_result[7][942] + xnor_result[7][943] + xnor_result[7][944] + xnor_result[7][945] + xnor_result[7][946] + xnor_result[7][947] + xnor_result[7][948] + xnor_result[7][949] + xnor_result[7][950] + xnor_result[7][951] + xnor_result[7][952] + xnor_result[7][953] + xnor_result[7][954] + xnor_result[7][955] + xnor_result[7][956] + xnor_result[7][957] + xnor_result[7][958] + xnor_result[7][959] ;
assign accumulation_result[8] = xnor_result[8][0] + xnor_result[8][1] + xnor_result[8][2] + xnor_result[8][3] + xnor_result[8][4] + xnor_result[8][5] + xnor_result[8][6] + xnor_result[8][7] + xnor_result[8][8] + xnor_result[8][9] + xnor_result[8][10] + xnor_result[8][11] + xnor_result[8][12] + xnor_result[8][13] + xnor_result[8][14] + xnor_result[8][15] + xnor_result[8][16] + xnor_result[8][17] + xnor_result[8][18] + xnor_result[8][19] + xnor_result[8][20] + xnor_result[8][21] + xnor_result[8][22] + xnor_result[8][23] + xnor_result[8][24] + xnor_result[8][25] + xnor_result[8][26] + xnor_result[8][27] + xnor_result[8][28] + xnor_result[8][29] + xnor_result[8][30] + xnor_result[8][31] + xnor_result[8][32] + xnor_result[8][33] + xnor_result[8][34] + xnor_result[8][35] + xnor_result[8][36] + xnor_result[8][37] + xnor_result[8][38] + xnor_result[8][39] + xnor_result[8][40] + xnor_result[8][41] + xnor_result[8][42] + xnor_result[8][43] + xnor_result[8][44] + xnor_result[8][45] + xnor_result[8][46] + xnor_result[8][47] + xnor_result[8][48] + xnor_result[8][49] + xnor_result[8][50] + xnor_result[8][51] + xnor_result[8][52] + xnor_result[8][53] + xnor_result[8][54] + xnor_result[8][55] + xnor_result[8][56] + xnor_result[8][57] + xnor_result[8][58] + xnor_result[8][59] + xnor_result[8][60] + xnor_result[8][61] + xnor_result[8][62] + xnor_result[8][63] + xnor_result[8][64] + xnor_result[8][65] + xnor_result[8][66] + xnor_result[8][67] + xnor_result[8][68] + xnor_result[8][69] + xnor_result[8][70] + xnor_result[8][71] + xnor_result[8][72] + xnor_result[8][73] + xnor_result[8][74] + xnor_result[8][75] + xnor_result[8][76] + xnor_result[8][77] + xnor_result[8][78] + xnor_result[8][79] + xnor_result[8][80] + xnor_result[8][81] + xnor_result[8][82] + xnor_result[8][83] + xnor_result[8][84] + xnor_result[8][85] + xnor_result[8][86] + xnor_result[8][87] + xnor_result[8][88] + xnor_result[8][89] + xnor_result[8][90] + xnor_result[8][91] + xnor_result[8][92] + xnor_result[8][93] + xnor_result[8][94] + xnor_result[8][95] + xnor_result[8][96] + xnor_result[8][97] + xnor_result[8][98] + xnor_result[8][99] + xnor_result[8][100] + xnor_result[8][101] + xnor_result[8][102] + xnor_result[8][103] + xnor_result[8][104] + xnor_result[8][105] + xnor_result[8][106] + xnor_result[8][107] + xnor_result[8][108] + xnor_result[8][109] + xnor_result[8][110] + xnor_result[8][111] + xnor_result[8][112] + xnor_result[8][113] + xnor_result[8][114] + xnor_result[8][115] + xnor_result[8][116] + xnor_result[8][117] + xnor_result[8][118] + xnor_result[8][119] + xnor_result[8][120] + xnor_result[8][121] + xnor_result[8][122] + xnor_result[8][123] + xnor_result[8][124] + xnor_result[8][125] + xnor_result[8][126] + xnor_result[8][127] + xnor_result[8][128] + xnor_result[8][129] + xnor_result[8][130] + xnor_result[8][131] + xnor_result[8][132] + xnor_result[8][133] + xnor_result[8][134] + xnor_result[8][135] + xnor_result[8][136] + xnor_result[8][137] + xnor_result[8][138] + xnor_result[8][139] + xnor_result[8][140] + xnor_result[8][141] + xnor_result[8][142] + xnor_result[8][143] + xnor_result[8][144] + xnor_result[8][145] + xnor_result[8][146] + xnor_result[8][147] + xnor_result[8][148] + xnor_result[8][149] + xnor_result[8][150] + xnor_result[8][151] + xnor_result[8][152] + xnor_result[8][153] + xnor_result[8][154] + xnor_result[8][155] + xnor_result[8][156] + xnor_result[8][157] + xnor_result[8][158] + xnor_result[8][159] + xnor_result[8][160] + xnor_result[8][161] + xnor_result[8][162] + xnor_result[8][163] + xnor_result[8][164] + xnor_result[8][165] + xnor_result[8][166] + xnor_result[8][167] + xnor_result[8][168] + xnor_result[8][169] + xnor_result[8][170] + xnor_result[8][171] + xnor_result[8][172] + xnor_result[8][173] + xnor_result[8][174] + xnor_result[8][175] + xnor_result[8][176] + xnor_result[8][177] + xnor_result[8][178] + xnor_result[8][179] + xnor_result[8][180] + xnor_result[8][181] + xnor_result[8][182] + xnor_result[8][183] + xnor_result[8][184] + xnor_result[8][185] + xnor_result[8][186] + xnor_result[8][187] + xnor_result[8][188] + xnor_result[8][189] + xnor_result[8][190] + xnor_result[8][191] + xnor_result[8][192] + xnor_result[8][193] + xnor_result[8][194] + xnor_result[8][195] + xnor_result[8][196] + xnor_result[8][197] + xnor_result[8][198] + xnor_result[8][199] + xnor_result[8][200] + xnor_result[8][201] + xnor_result[8][202] + xnor_result[8][203] + xnor_result[8][204] + xnor_result[8][205] + xnor_result[8][206] + xnor_result[8][207] + xnor_result[8][208] + xnor_result[8][209] + xnor_result[8][210] + xnor_result[8][211] + xnor_result[8][212] + xnor_result[8][213] + xnor_result[8][214] + xnor_result[8][215] + xnor_result[8][216] + xnor_result[8][217] + xnor_result[8][218] + xnor_result[8][219] + xnor_result[8][220] + xnor_result[8][221] + xnor_result[8][222] + xnor_result[8][223] + xnor_result[8][224] + xnor_result[8][225] + xnor_result[8][226] + xnor_result[8][227] + xnor_result[8][228] + xnor_result[8][229] + xnor_result[8][230] + xnor_result[8][231] + xnor_result[8][232] + xnor_result[8][233] + xnor_result[8][234] + xnor_result[8][235] + xnor_result[8][236] + xnor_result[8][237] + xnor_result[8][238] + xnor_result[8][239] + xnor_result[8][240] + xnor_result[8][241] + xnor_result[8][242] + xnor_result[8][243] + xnor_result[8][244] + xnor_result[8][245] + xnor_result[8][246] + xnor_result[8][247] + xnor_result[8][248] + xnor_result[8][249] + xnor_result[8][250] + xnor_result[8][251] + xnor_result[8][252] + xnor_result[8][253] + xnor_result[8][254] + xnor_result[8][255] + xnor_result[8][256] + xnor_result[8][257] + xnor_result[8][258] + xnor_result[8][259] + xnor_result[8][260] + xnor_result[8][261] + xnor_result[8][262] + xnor_result[8][263] + xnor_result[8][264] + xnor_result[8][265] + xnor_result[8][266] + xnor_result[8][267] + xnor_result[8][268] + xnor_result[8][269] + xnor_result[8][270] + xnor_result[8][271] + xnor_result[8][272] + xnor_result[8][273] + xnor_result[8][274] + xnor_result[8][275] + xnor_result[8][276] + xnor_result[8][277] + xnor_result[8][278] + xnor_result[8][279] + xnor_result[8][280] + xnor_result[8][281] + xnor_result[8][282] + xnor_result[8][283] + xnor_result[8][284] + xnor_result[8][285] + xnor_result[8][286] + xnor_result[8][287] + xnor_result[8][288] + xnor_result[8][289] + xnor_result[8][290] + xnor_result[8][291] + xnor_result[8][292] + xnor_result[8][293] + xnor_result[8][294] + xnor_result[8][295] + xnor_result[8][296] + xnor_result[8][297] + xnor_result[8][298] + xnor_result[8][299] + xnor_result[8][300] + xnor_result[8][301] + xnor_result[8][302] + xnor_result[8][303] + xnor_result[8][304] + xnor_result[8][305] + xnor_result[8][306] + xnor_result[8][307] + xnor_result[8][308] + xnor_result[8][309] + xnor_result[8][310] + xnor_result[8][311] + xnor_result[8][312] + xnor_result[8][313] + xnor_result[8][314] + xnor_result[8][315] + xnor_result[8][316] + xnor_result[8][317] + xnor_result[8][318] + xnor_result[8][319] + xnor_result[8][320] + xnor_result[8][321] + xnor_result[8][322] + xnor_result[8][323] + xnor_result[8][324] + xnor_result[8][325] + xnor_result[8][326] + xnor_result[8][327] + xnor_result[8][328] + xnor_result[8][329] + xnor_result[8][330] + xnor_result[8][331] + xnor_result[8][332] + xnor_result[8][333] + xnor_result[8][334] + xnor_result[8][335] + xnor_result[8][336] + xnor_result[8][337] + xnor_result[8][338] + xnor_result[8][339] + xnor_result[8][340] + xnor_result[8][341] + xnor_result[8][342] + xnor_result[8][343] + xnor_result[8][344] + xnor_result[8][345] + xnor_result[8][346] + xnor_result[8][347] + xnor_result[8][348] + xnor_result[8][349] + xnor_result[8][350] + xnor_result[8][351] + xnor_result[8][352] + xnor_result[8][353] + xnor_result[8][354] + xnor_result[8][355] + xnor_result[8][356] + xnor_result[8][357] + xnor_result[8][358] + xnor_result[8][359] + xnor_result[8][360] + xnor_result[8][361] + xnor_result[8][362] + xnor_result[8][363] + xnor_result[8][364] + xnor_result[8][365] + xnor_result[8][366] + xnor_result[8][367] + xnor_result[8][368] + xnor_result[8][369] + xnor_result[8][370] + xnor_result[8][371] + xnor_result[8][372] + xnor_result[8][373] + xnor_result[8][374] + xnor_result[8][375] + xnor_result[8][376] + xnor_result[8][377] + xnor_result[8][378] + xnor_result[8][379] + xnor_result[8][380] + xnor_result[8][381] + xnor_result[8][382] + xnor_result[8][383] + xnor_result[8][384] + xnor_result[8][385] + xnor_result[8][386] + xnor_result[8][387] + xnor_result[8][388] + xnor_result[8][389] + xnor_result[8][390] + xnor_result[8][391] + xnor_result[8][392] + xnor_result[8][393] + xnor_result[8][394] + xnor_result[8][395] + xnor_result[8][396] + xnor_result[8][397] + xnor_result[8][398] + xnor_result[8][399] + xnor_result[8][400] + xnor_result[8][401] + xnor_result[8][402] + xnor_result[8][403] + xnor_result[8][404] + xnor_result[8][405] + xnor_result[8][406] + xnor_result[8][407] + xnor_result[8][408] + xnor_result[8][409] + xnor_result[8][410] + xnor_result[8][411] + xnor_result[8][412] + xnor_result[8][413] + xnor_result[8][414] + xnor_result[8][415] + xnor_result[8][416] + xnor_result[8][417] + xnor_result[8][418] + xnor_result[8][419] + xnor_result[8][420] + xnor_result[8][421] + xnor_result[8][422] + xnor_result[8][423] + xnor_result[8][424] + xnor_result[8][425] + xnor_result[8][426] + xnor_result[8][427] + xnor_result[8][428] + xnor_result[8][429] + xnor_result[8][430] + xnor_result[8][431] + xnor_result[8][432] + xnor_result[8][433] + xnor_result[8][434] + xnor_result[8][435] + xnor_result[8][436] + xnor_result[8][437] + xnor_result[8][438] + xnor_result[8][439] + xnor_result[8][440] + xnor_result[8][441] + xnor_result[8][442] + xnor_result[8][443] + xnor_result[8][444] + xnor_result[8][445] + xnor_result[8][446] + xnor_result[8][447] + xnor_result[8][448] + xnor_result[8][449] + xnor_result[8][450] + xnor_result[8][451] + xnor_result[8][452] + xnor_result[8][453] + xnor_result[8][454] + xnor_result[8][455] + xnor_result[8][456] + xnor_result[8][457] + xnor_result[8][458] + xnor_result[8][459] + xnor_result[8][460] + xnor_result[8][461] + xnor_result[8][462] + xnor_result[8][463] + xnor_result[8][464] + xnor_result[8][465] + xnor_result[8][466] + xnor_result[8][467] + xnor_result[8][468] + xnor_result[8][469] + xnor_result[8][470] + xnor_result[8][471] + xnor_result[8][472] + xnor_result[8][473] + xnor_result[8][474] + xnor_result[8][475] + xnor_result[8][476] + xnor_result[8][477] + xnor_result[8][478] + xnor_result[8][479] + xnor_result[8][480] + xnor_result[8][481] + xnor_result[8][482] + xnor_result[8][483] + xnor_result[8][484] + xnor_result[8][485] + xnor_result[8][486] + xnor_result[8][487] + xnor_result[8][488] + xnor_result[8][489] + xnor_result[8][490] + xnor_result[8][491] + xnor_result[8][492] + xnor_result[8][493] + xnor_result[8][494] + xnor_result[8][495] + xnor_result[8][496] + xnor_result[8][497] + xnor_result[8][498] + xnor_result[8][499] + xnor_result[8][500] + xnor_result[8][501] + xnor_result[8][502] + xnor_result[8][503] + xnor_result[8][504] + xnor_result[8][505] + xnor_result[8][506] + xnor_result[8][507] + xnor_result[8][508] + xnor_result[8][509] + xnor_result[8][510] + xnor_result[8][511] + xnor_result[8][512] + xnor_result[8][513] + xnor_result[8][514] + xnor_result[8][515] + xnor_result[8][516] + xnor_result[8][517] + xnor_result[8][518] + xnor_result[8][519] + xnor_result[8][520] + xnor_result[8][521] + xnor_result[8][522] + xnor_result[8][523] + xnor_result[8][524] + xnor_result[8][525] + xnor_result[8][526] + xnor_result[8][527] + xnor_result[8][528] + xnor_result[8][529] + xnor_result[8][530] + xnor_result[8][531] + xnor_result[8][532] + xnor_result[8][533] + xnor_result[8][534] + xnor_result[8][535] + xnor_result[8][536] + xnor_result[8][537] + xnor_result[8][538] + xnor_result[8][539] + xnor_result[8][540] + xnor_result[8][541] + xnor_result[8][542] + xnor_result[8][543] + xnor_result[8][544] + xnor_result[8][545] + xnor_result[8][546] + xnor_result[8][547] + xnor_result[8][548] + xnor_result[8][549] + xnor_result[8][550] + xnor_result[8][551] + xnor_result[8][552] + xnor_result[8][553] + xnor_result[8][554] + xnor_result[8][555] + xnor_result[8][556] + xnor_result[8][557] + xnor_result[8][558] + xnor_result[8][559] + xnor_result[8][560] + xnor_result[8][561] + xnor_result[8][562] + xnor_result[8][563] + xnor_result[8][564] + xnor_result[8][565] + xnor_result[8][566] + xnor_result[8][567] + xnor_result[8][568] + xnor_result[8][569] + xnor_result[8][570] + xnor_result[8][571] + xnor_result[8][572] + xnor_result[8][573] + xnor_result[8][574] + xnor_result[8][575] + xnor_result[8][576] + xnor_result[8][577] + xnor_result[8][578] + xnor_result[8][579] + xnor_result[8][580] + xnor_result[8][581] + xnor_result[8][582] + xnor_result[8][583] + xnor_result[8][584] + xnor_result[8][585] + xnor_result[8][586] + xnor_result[8][587] + xnor_result[8][588] + xnor_result[8][589] + xnor_result[8][590] + xnor_result[8][591] + xnor_result[8][592] + xnor_result[8][593] + xnor_result[8][594] + xnor_result[8][595] + xnor_result[8][596] + xnor_result[8][597] + xnor_result[8][598] + xnor_result[8][599] + xnor_result[8][600] + xnor_result[8][601] + xnor_result[8][602] + xnor_result[8][603] + xnor_result[8][604] + xnor_result[8][605] + xnor_result[8][606] + xnor_result[8][607] + xnor_result[8][608] + xnor_result[8][609] + xnor_result[8][610] + xnor_result[8][611] + xnor_result[8][612] + xnor_result[8][613] + xnor_result[8][614] + xnor_result[8][615] + xnor_result[8][616] + xnor_result[8][617] + xnor_result[8][618] + xnor_result[8][619] + xnor_result[8][620] + xnor_result[8][621] + xnor_result[8][622] + xnor_result[8][623] + xnor_result[8][624] + xnor_result[8][625] + xnor_result[8][626] + xnor_result[8][627] + xnor_result[8][628] + xnor_result[8][629] + xnor_result[8][630] + xnor_result[8][631] + xnor_result[8][632] + xnor_result[8][633] + xnor_result[8][634] + xnor_result[8][635] + xnor_result[8][636] + xnor_result[8][637] + xnor_result[8][638] + xnor_result[8][639] + xnor_result[8][640] + xnor_result[8][641] + xnor_result[8][642] + xnor_result[8][643] + xnor_result[8][644] + xnor_result[8][645] + xnor_result[8][646] + xnor_result[8][647] + xnor_result[8][648] + xnor_result[8][649] + xnor_result[8][650] + xnor_result[8][651] + xnor_result[8][652] + xnor_result[8][653] + xnor_result[8][654] + xnor_result[8][655] + xnor_result[8][656] + xnor_result[8][657] + xnor_result[8][658] + xnor_result[8][659] + xnor_result[8][660] + xnor_result[8][661] + xnor_result[8][662] + xnor_result[8][663] + xnor_result[8][664] + xnor_result[8][665] + xnor_result[8][666] + xnor_result[8][667] + xnor_result[8][668] + xnor_result[8][669] + xnor_result[8][670] + xnor_result[8][671] + xnor_result[8][672] + xnor_result[8][673] + xnor_result[8][674] + xnor_result[8][675] + xnor_result[8][676] + xnor_result[8][677] + xnor_result[8][678] + xnor_result[8][679] + xnor_result[8][680] + xnor_result[8][681] + xnor_result[8][682] + xnor_result[8][683] + xnor_result[8][684] + xnor_result[8][685] + xnor_result[8][686] + xnor_result[8][687] + xnor_result[8][688] + xnor_result[8][689] + xnor_result[8][690] + xnor_result[8][691] + xnor_result[8][692] + xnor_result[8][693] + xnor_result[8][694] + xnor_result[8][695] + xnor_result[8][696] + xnor_result[8][697] + xnor_result[8][698] + xnor_result[8][699] + xnor_result[8][700] + xnor_result[8][701] + xnor_result[8][702] + xnor_result[8][703] + xnor_result[8][704] + xnor_result[8][705] + xnor_result[8][706] + xnor_result[8][707] + xnor_result[8][708] + xnor_result[8][709] + xnor_result[8][710] + xnor_result[8][711] + xnor_result[8][712] + xnor_result[8][713] + xnor_result[8][714] + xnor_result[8][715] + xnor_result[8][716] + xnor_result[8][717] + xnor_result[8][718] + xnor_result[8][719] + xnor_result[8][720] + xnor_result[8][721] + xnor_result[8][722] + xnor_result[8][723] + xnor_result[8][724] + xnor_result[8][725] + xnor_result[8][726] + xnor_result[8][727] + xnor_result[8][728] + xnor_result[8][729] + xnor_result[8][730] + xnor_result[8][731] + xnor_result[8][732] + xnor_result[8][733] + xnor_result[8][734] + xnor_result[8][735] + xnor_result[8][736] + xnor_result[8][737] + xnor_result[8][738] + xnor_result[8][739] + xnor_result[8][740] + xnor_result[8][741] + xnor_result[8][742] + xnor_result[8][743] + xnor_result[8][744] + xnor_result[8][745] + xnor_result[8][746] + xnor_result[8][747] + xnor_result[8][748] + xnor_result[8][749] + xnor_result[8][750] + xnor_result[8][751] + xnor_result[8][752] + xnor_result[8][753] + xnor_result[8][754] + xnor_result[8][755] + xnor_result[8][756] + xnor_result[8][757] + xnor_result[8][758] + xnor_result[8][759] + xnor_result[8][760] + xnor_result[8][761] + xnor_result[8][762] + xnor_result[8][763] + xnor_result[8][764] + xnor_result[8][765] + xnor_result[8][766] + xnor_result[8][767] + xnor_result[8][768] + xnor_result[8][769] + xnor_result[8][770] + xnor_result[8][771] + xnor_result[8][772] + xnor_result[8][773] + xnor_result[8][774] + xnor_result[8][775] + xnor_result[8][776] + xnor_result[8][777] + xnor_result[8][778] + xnor_result[8][779] + xnor_result[8][780] + xnor_result[8][781] + xnor_result[8][782] + xnor_result[8][783] + xnor_result[8][784] + xnor_result[8][785] + xnor_result[8][786] + xnor_result[8][787] + xnor_result[8][788] + xnor_result[8][789] + xnor_result[8][790] + xnor_result[8][791] + xnor_result[8][792] + xnor_result[8][793] + xnor_result[8][794] + xnor_result[8][795] + xnor_result[8][796] + xnor_result[8][797] + xnor_result[8][798] + xnor_result[8][799] + xnor_result[8][800] + xnor_result[8][801] + xnor_result[8][802] + xnor_result[8][803] + xnor_result[8][804] + xnor_result[8][805] + xnor_result[8][806] + xnor_result[8][807] + xnor_result[8][808] + xnor_result[8][809] + xnor_result[8][810] + xnor_result[8][811] + xnor_result[8][812] + xnor_result[8][813] + xnor_result[8][814] + xnor_result[8][815] + xnor_result[8][816] + xnor_result[8][817] + xnor_result[8][818] + xnor_result[8][819] + xnor_result[8][820] + xnor_result[8][821] + xnor_result[8][822] + xnor_result[8][823] + xnor_result[8][824] + xnor_result[8][825] + xnor_result[8][826] + xnor_result[8][827] + xnor_result[8][828] + xnor_result[8][829] + xnor_result[8][830] + xnor_result[8][831] + xnor_result[8][832] + xnor_result[8][833] + xnor_result[8][834] + xnor_result[8][835] + xnor_result[8][836] + xnor_result[8][837] + xnor_result[8][838] + xnor_result[8][839] + xnor_result[8][840] + xnor_result[8][841] + xnor_result[8][842] + xnor_result[8][843] + xnor_result[8][844] + xnor_result[8][845] + xnor_result[8][846] + xnor_result[8][847] + xnor_result[8][848] + xnor_result[8][849] + xnor_result[8][850] + xnor_result[8][851] + xnor_result[8][852] + xnor_result[8][853] + xnor_result[8][854] + xnor_result[8][855] + xnor_result[8][856] + xnor_result[8][857] + xnor_result[8][858] + xnor_result[8][859] + xnor_result[8][860] + xnor_result[8][861] + xnor_result[8][862] + xnor_result[8][863] + xnor_result[8][864] + xnor_result[8][865] + xnor_result[8][866] + xnor_result[8][867] + xnor_result[8][868] + xnor_result[8][869] + xnor_result[8][870] + xnor_result[8][871] + xnor_result[8][872] + xnor_result[8][873] + xnor_result[8][874] + xnor_result[8][875] + xnor_result[8][876] + xnor_result[8][877] + xnor_result[8][878] + xnor_result[8][879] + xnor_result[8][880] + xnor_result[8][881] + xnor_result[8][882] + xnor_result[8][883] + xnor_result[8][884] + xnor_result[8][885] + xnor_result[8][886] + xnor_result[8][887] + xnor_result[8][888] + xnor_result[8][889] + xnor_result[8][890] + xnor_result[8][891] + xnor_result[8][892] + xnor_result[8][893] + xnor_result[8][894] + xnor_result[8][895] + xnor_result[8][896] + xnor_result[8][897] + xnor_result[8][898] + xnor_result[8][899] + xnor_result[8][900] + xnor_result[8][901] + xnor_result[8][902] + xnor_result[8][903] + xnor_result[8][904] + xnor_result[8][905] + xnor_result[8][906] + xnor_result[8][907] + xnor_result[8][908] + xnor_result[8][909] + xnor_result[8][910] + xnor_result[8][911] + xnor_result[8][912] + xnor_result[8][913] + xnor_result[8][914] + xnor_result[8][915] + xnor_result[8][916] + xnor_result[8][917] + xnor_result[8][918] + xnor_result[8][919] + xnor_result[8][920] + xnor_result[8][921] + xnor_result[8][922] + xnor_result[8][923] + xnor_result[8][924] + xnor_result[8][925] + xnor_result[8][926] + xnor_result[8][927] + xnor_result[8][928] + xnor_result[8][929] + xnor_result[8][930] + xnor_result[8][931] + xnor_result[8][932] + xnor_result[8][933] + xnor_result[8][934] + xnor_result[8][935] + xnor_result[8][936] + xnor_result[8][937] + xnor_result[8][938] + xnor_result[8][939] + xnor_result[8][940] + xnor_result[8][941] + xnor_result[8][942] + xnor_result[8][943] + xnor_result[8][944] + xnor_result[8][945] + xnor_result[8][946] + xnor_result[8][947] + xnor_result[8][948] + xnor_result[8][949] + xnor_result[8][950] + xnor_result[8][951] + xnor_result[8][952] + xnor_result[8][953] + xnor_result[8][954] + xnor_result[8][955] + xnor_result[8][956] + xnor_result[8][957] + xnor_result[8][958] + xnor_result[8][959] ;
assign accumulation_result[9] = xnor_result[9][0] + xnor_result[9][1] + xnor_result[9][2] + xnor_result[9][3] + xnor_result[9][4] + xnor_result[9][5] + xnor_result[9][6] + xnor_result[9][7] + xnor_result[9][8] + xnor_result[9][9] + xnor_result[9][10] + xnor_result[9][11] + xnor_result[9][12] + xnor_result[9][13] + xnor_result[9][14] + xnor_result[9][15] + xnor_result[9][16] + xnor_result[9][17] + xnor_result[9][18] + xnor_result[9][19] + xnor_result[9][20] + xnor_result[9][21] + xnor_result[9][22] + xnor_result[9][23] + xnor_result[9][24] + xnor_result[9][25] + xnor_result[9][26] + xnor_result[9][27] + xnor_result[9][28] + xnor_result[9][29] + xnor_result[9][30] + xnor_result[9][31] + xnor_result[9][32] + xnor_result[9][33] + xnor_result[9][34] + xnor_result[9][35] + xnor_result[9][36] + xnor_result[9][37] + xnor_result[9][38] + xnor_result[9][39] + xnor_result[9][40] + xnor_result[9][41] + xnor_result[9][42] + xnor_result[9][43] + xnor_result[9][44] + xnor_result[9][45] + xnor_result[9][46] + xnor_result[9][47] + xnor_result[9][48] + xnor_result[9][49] + xnor_result[9][50] + xnor_result[9][51] + xnor_result[9][52] + xnor_result[9][53] + xnor_result[9][54] + xnor_result[9][55] + xnor_result[9][56] + xnor_result[9][57] + xnor_result[9][58] + xnor_result[9][59] + xnor_result[9][60] + xnor_result[9][61] + xnor_result[9][62] + xnor_result[9][63] + xnor_result[9][64] + xnor_result[9][65] + xnor_result[9][66] + xnor_result[9][67] + xnor_result[9][68] + xnor_result[9][69] + xnor_result[9][70] + xnor_result[9][71] + xnor_result[9][72] + xnor_result[9][73] + xnor_result[9][74] + xnor_result[9][75] + xnor_result[9][76] + xnor_result[9][77] + xnor_result[9][78] + xnor_result[9][79] + xnor_result[9][80] + xnor_result[9][81] + xnor_result[9][82] + xnor_result[9][83] + xnor_result[9][84] + xnor_result[9][85] + xnor_result[9][86] + xnor_result[9][87] + xnor_result[9][88] + xnor_result[9][89] + xnor_result[9][90] + xnor_result[9][91] + xnor_result[9][92] + xnor_result[9][93] + xnor_result[9][94] + xnor_result[9][95] + xnor_result[9][96] + xnor_result[9][97] + xnor_result[9][98] + xnor_result[9][99] + xnor_result[9][100] + xnor_result[9][101] + xnor_result[9][102] + xnor_result[9][103] + xnor_result[9][104] + xnor_result[9][105] + xnor_result[9][106] + xnor_result[9][107] + xnor_result[9][108] + xnor_result[9][109] + xnor_result[9][110] + xnor_result[9][111] + xnor_result[9][112] + xnor_result[9][113] + xnor_result[9][114] + xnor_result[9][115] + xnor_result[9][116] + xnor_result[9][117] + xnor_result[9][118] + xnor_result[9][119] + xnor_result[9][120] + xnor_result[9][121] + xnor_result[9][122] + xnor_result[9][123] + xnor_result[9][124] + xnor_result[9][125] + xnor_result[9][126] + xnor_result[9][127] + xnor_result[9][128] + xnor_result[9][129] + xnor_result[9][130] + xnor_result[9][131] + xnor_result[9][132] + xnor_result[9][133] + xnor_result[9][134] + xnor_result[9][135] + xnor_result[9][136] + xnor_result[9][137] + xnor_result[9][138] + xnor_result[9][139] + xnor_result[9][140] + xnor_result[9][141] + xnor_result[9][142] + xnor_result[9][143] + xnor_result[9][144] + xnor_result[9][145] + xnor_result[9][146] + xnor_result[9][147] + xnor_result[9][148] + xnor_result[9][149] + xnor_result[9][150] + xnor_result[9][151] + xnor_result[9][152] + xnor_result[9][153] + xnor_result[9][154] + xnor_result[9][155] + xnor_result[9][156] + xnor_result[9][157] + xnor_result[9][158] + xnor_result[9][159] + xnor_result[9][160] + xnor_result[9][161] + xnor_result[9][162] + xnor_result[9][163] + xnor_result[9][164] + xnor_result[9][165] + xnor_result[9][166] + xnor_result[9][167] + xnor_result[9][168] + xnor_result[9][169] + xnor_result[9][170] + xnor_result[9][171] + xnor_result[9][172] + xnor_result[9][173] + xnor_result[9][174] + xnor_result[9][175] + xnor_result[9][176] + xnor_result[9][177] + xnor_result[9][178] + xnor_result[9][179] + xnor_result[9][180] + xnor_result[9][181] + xnor_result[9][182] + xnor_result[9][183] + xnor_result[9][184] + xnor_result[9][185] + xnor_result[9][186] + xnor_result[9][187] + xnor_result[9][188] + xnor_result[9][189] + xnor_result[9][190] + xnor_result[9][191] + xnor_result[9][192] + xnor_result[9][193] + xnor_result[9][194] + xnor_result[9][195] + xnor_result[9][196] + xnor_result[9][197] + xnor_result[9][198] + xnor_result[9][199] + xnor_result[9][200] + xnor_result[9][201] + xnor_result[9][202] + xnor_result[9][203] + xnor_result[9][204] + xnor_result[9][205] + xnor_result[9][206] + xnor_result[9][207] + xnor_result[9][208] + xnor_result[9][209] + xnor_result[9][210] + xnor_result[9][211] + xnor_result[9][212] + xnor_result[9][213] + xnor_result[9][214] + xnor_result[9][215] + xnor_result[9][216] + xnor_result[9][217] + xnor_result[9][218] + xnor_result[9][219] + xnor_result[9][220] + xnor_result[9][221] + xnor_result[9][222] + xnor_result[9][223] + xnor_result[9][224] + xnor_result[9][225] + xnor_result[9][226] + xnor_result[9][227] + xnor_result[9][228] + xnor_result[9][229] + xnor_result[9][230] + xnor_result[9][231] + xnor_result[9][232] + xnor_result[9][233] + xnor_result[9][234] + xnor_result[9][235] + xnor_result[9][236] + xnor_result[9][237] + xnor_result[9][238] + xnor_result[9][239] + xnor_result[9][240] + xnor_result[9][241] + xnor_result[9][242] + xnor_result[9][243] + xnor_result[9][244] + xnor_result[9][245] + xnor_result[9][246] + xnor_result[9][247] + xnor_result[9][248] + xnor_result[9][249] + xnor_result[9][250] + xnor_result[9][251] + xnor_result[9][252] + xnor_result[9][253] + xnor_result[9][254] + xnor_result[9][255] + xnor_result[9][256] + xnor_result[9][257] + xnor_result[9][258] + xnor_result[9][259] + xnor_result[9][260] + xnor_result[9][261] + xnor_result[9][262] + xnor_result[9][263] + xnor_result[9][264] + xnor_result[9][265] + xnor_result[9][266] + xnor_result[9][267] + xnor_result[9][268] + xnor_result[9][269] + xnor_result[9][270] + xnor_result[9][271] + xnor_result[9][272] + xnor_result[9][273] + xnor_result[9][274] + xnor_result[9][275] + xnor_result[9][276] + xnor_result[9][277] + xnor_result[9][278] + xnor_result[9][279] + xnor_result[9][280] + xnor_result[9][281] + xnor_result[9][282] + xnor_result[9][283] + xnor_result[9][284] + xnor_result[9][285] + xnor_result[9][286] + xnor_result[9][287] + xnor_result[9][288] + xnor_result[9][289] + xnor_result[9][290] + xnor_result[9][291] + xnor_result[9][292] + xnor_result[9][293] + xnor_result[9][294] + xnor_result[9][295] + xnor_result[9][296] + xnor_result[9][297] + xnor_result[9][298] + xnor_result[9][299] + xnor_result[9][300] + xnor_result[9][301] + xnor_result[9][302] + xnor_result[9][303] + xnor_result[9][304] + xnor_result[9][305] + xnor_result[9][306] + xnor_result[9][307] + xnor_result[9][308] + xnor_result[9][309] + xnor_result[9][310] + xnor_result[9][311] + xnor_result[9][312] + xnor_result[9][313] + xnor_result[9][314] + xnor_result[9][315] + xnor_result[9][316] + xnor_result[9][317] + xnor_result[9][318] + xnor_result[9][319] + xnor_result[9][320] + xnor_result[9][321] + xnor_result[9][322] + xnor_result[9][323] + xnor_result[9][324] + xnor_result[9][325] + xnor_result[9][326] + xnor_result[9][327] + xnor_result[9][328] + xnor_result[9][329] + xnor_result[9][330] + xnor_result[9][331] + xnor_result[9][332] + xnor_result[9][333] + xnor_result[9][334] + xnor_result[9][335] + xnor_result[9][336] + xnor_result[9][337] + xnor_result[9][338] + xnor_result[9][339] + xnor_result[9][340] + xnor_result[9][341] + xnor_result[9][342] + xnor_result[9][343] + xnor_result[9][344] + xnor_result[9][345] + xnor_result[9][346] + xnor_result[9][347] + xnor_result[9][348] + xnor_result[9][349] + xnor_result[9][350] + xnor_result[9][351] + xnor_result[9][352] + xnor_result[9][353] + xnor_result[9][354] + xnor_result[9][355] + xnor_result[9][356] + xnor_result[9][357] + xnor_result[9][358] + xnor_result[9][359] + xnor_result[9][360] + xnor_result[9][361] + xnor_result[9][362] + xnor_result[9][363] + xnor_result[9][364] + xnor_result[9][365] + xnor_result[9][366] + xnor_result[9][367] + xnor_result[9][368] + xnor_result[9][369] + xnor_result[9][370] + xnor_result[9][371] + xnor_result[9][372] + xnor_result[9][373] + xnor_result[9][374] + xnor_result[9][375] + xnor_result[9][376] + xnor_result[9][377] + xnor_result[9][378] + xnor_result[9][379] + xnor_result[9][380] + xnor_result[9][381] + xnor_result[9][382] + xnor_result[9][383] + xnor_result[9][384] + xnor_result[9][385] + xnor_result[9][386] + xnor_result[9][387] + xnor_result[9][388] + xnor_result[9][389] + xnor_result[9][390] + xnor_result[9][391] + xnor_result[9][392] + xnor_result[9][393] + xnor_result[9][394] + xnor_result[9][395] + xnor_result[9][396] + xnor_result[9][397] + xnor_result[9][398] + xnor_result[9][399] + xnor_result[9][400] + xnor_result[9][401] + xnor_result[9][402] + xnor_result[9][403] + xnor_result[9][404] + xnor_result[9][405] + xnor_result[9][406] + xnor_result[9][407] + xnor_result[9][408] + xnor_result[9][409] + xnor_result[9][410] + xnor_result[9][411] + xnor_result[9][412] + xnor_result[9][413] + xnor_result[9][414] + xnor_result[9][415] + xnor_result[9][416] + xnor_result[9][417] + xnor_result[9][418] + xnor_result[9][419] + xnor_result[9][420] + xnor_result[9][421] + xnor_result[9][422] + xnor_result[9][423] + xnor_result[9][424] + xnor_result[9][425] + xnor_result[9][426] + xnor_result[9][427] + xnor_result[9][428] + xnor_result[9][429] + xnor_result[9][430] + xnor_result[9][431] + xnor_result[9][432] + xnor_result[9][433] + xnor_result[9][434] + xnor_result[9][435] + xnor_result[9][436] + xnor_result[9][437] + xnor_result[9][438] + xnor_result[9][439] + xnor_result[9][440] + xnor_result[9][441] + xnor_result[9][442] + xnor_result[9][443] + xnor_result[9][444] + xnor_result[9][445] + xnor_result[9][446] + xnor_result[9][447] + xnor_result[9][448] + xnor_result[9][449] + xnor_result[9][450] + xnor_result[9][451] + xnor_result[9][452] + xnor_result[9][453] + xnor_result[9][454] + xnor_result[9][455] + xnor_result[9][456] + xnor_result[9][457] + xnor_result[9][458] + xnor_result[9][459] + xnor_result[9][460] + xnor_result[9][461] + xnor_result[9][462] + xnor_result[9][463] + xnor_result[9][464] + xnor_result[9][465] + xnor_result[9][466] + xnor_result[9][467] + xnor_result[9][468] + xnor_result[9][469] + xnor_result[9][470] + xnor_result[9][471] + xnor_result[9][472] + xnor_result[9][473] + xnor_result[9][474] + xnor_result[9][475] + xnor_result[9][476] + xnor_result[9][477] + xnor_result[9][478] + xnor_result[9][479] + xnor_result[9][480] + xnor_result[9][481] + xnor_result[9][482] + xnor_result[9][483] + xnor_result[9][484] + xnor_result[9][485] + xnor_result[9][486] + xnor_result[9][487] + xnor_result[9][488] + xnor_result[9][489] + xnor_result[9][490] + xnor_result[9][491] + xnor_result[9][492] + xnor_result[9][493] + xnor_result[9][494] + xnor_result[9][495] + xnor_result[9][496] + xnor_result[9][497] + xnor_result[9][498] + xnor_result[9][499] + xnor_result[9][500] + xnor_result[9][501] + xnor_result[9][502] + xnor_result[9][503] + xnor_result[9][504] + xnor_result[9][505] + xnor_result[9][506] + xnor_result[9][507] + xnor_result[9][508] + xnor_result[9][509] + xnor_result[9][510] + xnor_result[9][511] + xnor_result[9][512] + xnor_result[9][513] + xnor_result[9][514] + xnor_result[9][515] + xnor_result[9][516] + xnor_result[9][517] + xnor_result[9][518] + xnor_result[9][519] + xnor_result[9][520] + xnor_result[9][521] + xnor_result[9][522] + xnor_result[9][523] + xnor_result[9][524] + xnor_result[9][525] + xnor_result[9][526] + xnor_result[9][527] + xnor_result[9][528] + xnor_result[9][529] + xnor_result[9][530] + xnor_result[9][531] + xnor_result[9][532] + xnor_result[9][533] + xnor_result[9][534] + xnor_result[9][535] + xnor_result[9][536] + xnor_result[9][537] + xnor_result[9][538] + xnor_result[9][539] + xnor_result[9][540] + xnor_result[9][541] + xnor_result[9][542] + xnor_result[9][543] + xnor_result[9][544] + xnor_result[9][545] + xnor_result[9][546] + xnor_result[9][547] + xnor_result[9][548] + xnor_result[9][549] + xnor_result[9][550] + xnor_result[9][551] + xnor_result[9][552] + xnor_result[9][553] + xnor_result[9][554] + xnor_result[9][555] + xnor_result[9][556] + xnor_result[9][557] + xnor_result[9][558] + xnor_result[9][559] + xnor_result[9][560] + xnor_result[9][561] + xnor_result[9][562] + xnor_result[9][563] + xnor_result[9][564] + xnor_result[9][565] + xnor_result[9][566] + xnor_result[9][567] + xnor_result[9][568] + xnor_result[9][569] + xnor_result[9][570] + xnor_result[9][571] + xnor_result[9][572] + xnor_result[9][573] + xnor_result[9][574] + xnor_result[9][575] + xnor_result[9][576] + xnor_result[9][577] + xnor_result[9][578] + xnor_result[9][579] + xnor_result[9][580] + xnor_result[9][581] + xnor_result[9][582] + xnor_result[9][583] + xnor_result[9][584] + xnor_result[9][585] + xnor_result[9][586] + xnor_result[9][587] + xnor_result[9][588] + xnor_result[9][589] + xnor_result[9][590] + xnor_result[9][591] + xnor_result[9][592] + xnor_result[9][593] + xnor_result[9][594] + xnor_result[9][595] + xnor_result[9][596] + xnor_result[9][597] + xnor_result[9][598] + xnor_result[9][599] + xnor_result[9][600] + xnor_result[9][601] + xnor_result[9][602] + xnor_result[9][603] + xnor_result[9][604] + xnor_result[9][605] + xnor_result[9][606] + xnor_result[9][607] + xnor_result[9][608] + xnor_result[9][609] + xnor_result[9][610] + xnor_result[9][611] + xnor_result[9][612] + xnor_result[9][613] + xnor_result[9][614] + xnor_result[9][615] + xnor_result[9][616] + xnor_result[9][617] + xnor_result[9][618] + xnor_result[9][619] + xnor_result[9][620] + xnor_result[9][621] + xnor_result[9][622] + xnor_result[9][623] + xnor_result[9][624] + xnor_result[9][625] + xnor_result[9][626] + xnor_result[9][627] + xnor_result[9][628] + xnor_result[9][629] + xnor_result[9][630] + xnor_result[9][631] + xnor_result[9][632] + xnor_result[9][633] + xnor_result[9][634] + xnor_result[9][635] + xnor_result[9][636] + xnor_result[9][637] + xnor_result[9][638] + xnor_result[9][639] + xnor_result[9][640] + xnor_result[9][641] + xnor_result[9][642] + xnor_result[9][643] + xnor_result[9][644] + xnor_result[9][645] + xnor_result[9][646] + xnor_result[9][647] + xnor_result[9][648] + xnor_result[9][649] + xnor_result[9][650] + xnor_result[9][651] + xnor_result[9][652] + xnor_result[9][653] + xnor_result[9][654] + xnor_result[9][655] + xnor_result[9][656] + xnor_result[9][657] + xnor_result[9][658] + xnor_result[9][659] + xnor_result[9][660] + xnor_result[9][661] + xnor_result[9][662] + xnor_result[9][663] + xnor_result[9][664] + xnor_result[9][665] + xnor_result[9][666] + xnor_result[9][667] + xnor_result[9][668] + xnor_result[9][669] + xnor_result[9][670] + xnor_result[9][671] + xnor_result[9][672] + xnor_result[9][673] + xnor_result[9][674] + xnor_result[9][675] + xnor_result[9][676] + xnor_result[9][677] + xnor_result[9][678] + xnor_result[9][679] + xnor_result[9][680] + xnor_result[9][681] + xnor_result[9][682] + xnor_result[9][683] + xnor_result[9][684] + xnor_result[9][685] + xnor_result[9][686] + xnor_result[9][687] + xnor_result[9][688] + xnor_result[9][689] + xnor_result[9][690] + xnor_result[9][691] + xnor_result[9][692] + xnor_result[9][693] + xnor_result[9][694] + xnor_result[9][695] + xnor_result[9][696] + xnor_result[9][697] + xnor_result[9][698] + xnor_result[9][699] + xnor_result[9][700] + xnor_result[9][701] + xnor_result[9][702] + xnor_result[9][703] + xnor_result[9][704] + xnor_result[9][705] + xnor_result[9][706] + xnor_result[9][707] + xnor_result[9][708] + xnor_result[9][709] + xnor_result[9][710] + xnor_result[9][711] + xnor_result[9][712] + xnor_result[9][713] + xnor_result[9][714] + xnor_result[9][715] + xnor_result[9][716] + xnor_result[9][717] + xnor_result[9][718] + xnor_result[9][719] + xnor_result[9][720] + xnor_result[9][721] + xnor_result[9][722] + xnor_result[9][723] + xnor_result[9][724] + xnor_result[9][725] + xnor_result[9][726] + xnor_result[9][727] + xnor_result[9][728] + xnor_result[9][729] + xnor_result[9][730] + xnor_result[9][731] + xnor_result[9][732] + xnor_result[9][733] + xnor_result[9][734] + xnor_result[9][735] + xnor_result[9][736] + xnor_result[9][737] + xnor_result[9][738] + xnor_result[9][739] + xnor_result[9][740] + xnor_result[9][741] + xnor_result[9][742] + xnor_result[9][743] + xnor_result[9][744] + xnor_result[9][745] + xnor_result[9][746] + xnor_result[9][747] + xnor_result[9][748] + xnor_result[9][749] + xnor_result[9][750] + xnor_result[9][751] + xnor_result[9][752] + xnor_result[9][753] + xnor_result[9][754] + xnor_result[9][755] + xnor_result[9][756] + xnor_result[9][757] + xnor_result[9][758] + xnor_result[9][759] + xnor_result[9][760] + xnor_result[9][761] + xnor_result[9][762] + xnor_result[9][763] + xnor_result[9][764] + xnor_result[9][765] + xnor_result[9][766] + xnor_result[9][767] + xnor_result[9][768] + xnor_result[9][769] + xnor_result[9][770] + xnor_result[9][771] + xnor_result[9][772] + xnor_result[9][773] + xnor_result[9][774] + xnor_result[9][775] + xnor_result[9][776] + xnor_result[9][777] + xnor_result[9][778] + xnor_result[9][779] + xnor_result[9][780] + xnor_result[9][781] + xnor_result[9][782] + xnor_result[9][783] + xnor_result[9][784] + xnor_result[9][785] + xnor_result[9][786] + xnor_result[9][787] + xnor_result[9][788] + xnor_result[9][789] + xnor_result[9][790] + xnor_result[9][791] + xnor_result[9][792] + xnor_result[9][793] + xnor_result[9][794] + xnor_result[9][795] + xnor_result[9][796] + xnor_result[9][797] + xnor_result[9][798] + xnor_result[9][799] + xnor_result[9][800] + xnor_result[9][801] + xnor_result[9][802] + xnor_result[9][803] + xnor_result[9][804] + xnor_result[9][805] + xnor_result[9][806] + xnor_result[9][807] + xnor_result[9][808] + xnor_result[9][809] + xnor_result[9][810] + xnor_result[9][811] + xnor_result[9][812] + xnor_result[9][813] + xnor_result[9][814] + xnor_result[9][815] + xnor_result[9][816] + xnor_result[9][817] + xnor_result[9][818] + xnor_result[9][819] + xnor_result[9][820] + xnor_result[9][821] + xnor_result[9][822] + xnor_result[9][823] + xnor_result[9][824] + xnor_result[9][825] + xnor_result[9][826] + xnor_result[9][827] + xnor_result[9][828] + xnor_result[9][829] + xnor_result[9][830] + xnor_result[9][831] + xnor_result[9][832] + xnor_result[9][833] + xnor_result[9][834] + xnor_result[9][835] + xnor_result[9][836] + xnor_result[9][837] + xnor_result[9][838] + xnor_result[9][839] + xnor_result[9][840] + xnor_result[9][841] + xnor_result[9][842] + xnor_result[9][843] + xnor_result[9][844] + xnor_result[9][845] + xnor_result[9][846] + xnor_result[9][847] + xnor_result[9][848] + xnor_result[9][849] + xnor_result[9][850] + xnor_result[9][851] + xnor_result[9][852] + xnor_result[9][853] + xnor_result[9][854] + xnor_result[9][855] + xnor_result[9][856] + xnor_result[9][857] + xnor_result[9][858] + xnor_result[9][859] + xnor_result[9][860] + xnor_result[9][861] + xnor_result[9][862] + xnor_result[9][863] + xnor_result[9][864] + xnor_result[9][865] + xnor_result[9][866] + xnor_result[9][867] + xnor_result[9][868] + xnor_result[9][869] + xnor_result[9][870] + xnor_result[9][871] + xnor_result[9][872] + xnor_result[9][873] + xnor_result[9][874] + xnor_result[9][875] + xnor_result[9][876] + xnor_result[9][877] + xnor_result[9][878] + xnor_result[9][879] + xnor_result[9][880] + xnor_result[9][881] + xnor_result[9][882] + xnor_result[9][883] + xnor_result[9][884] + xnor_result[9][885] + xnor_result[9][886] + xnor_result[9][887] + xnor_result[9][888] + xnor_result[9][889] + xnor_result[9][890] + xnor_result[9][891] + xnor_result[9][892] + xnor_result[9][893] + xnor_result[9][894] + xnor_result[9][895] + xnor_result[9][896] + xnor_result[9][897] + xnor_result[9][898] + xnor_result[9][899] + xnor_result[9][900] + xnor_result[9][901] + xnor_result[9][902] + xnor_result[9][903] + xnor_result[9][904] + xnor_result[9][905] + xnor_result[9][906] + xnor_result[9][907] + xnor_result[9][908] + xnor_result[9][909] + xnor_result[9][910] + xnor_result[9][911] + xnor_result[9][912] + xnor_result[9][913] + xnor_result[9][914] + xnor_result[9][915] + xnor_result[9][916] + xnor_result[9][917] + xnor_result[9][918] + xnor_result[9][919] + xnor_result[9][920] + xnor_result[9][921] + xnor_result[9][922] + xnor_result[9][923] + xnor_result[9][924] + xnor_result[9][925] + xnor_result[9][926] + xnor_result[9][927] + xnor_result[9][928] + xnor_result[9][929] + xnor_result[9][930] + xnor_result[9][931] + xnor_result[9][932] + xnor_result[9][933] + xnor_result[9][934] + xnor_result[9][935] + xnor_result[9][936] + xnor_result[9][937] + xnor_result[9][938] + xnor_result[9][939] + xnor_result[9][940] + xnor_result[9][941] + xnor_result[9][942] + xnor_result[9][943] + xnor_result[9][944] + xnor_result[9][945] + xnor_result[9][946] + xnor_result[9][947] + xnor_result[9][948] + xnor_result[9][949] + xnor_result[9][950] + xnor_result[9][951] + xnor_result[9][952] + xnor_result[9][953] + xnor_result[9][954] + xnor_result[9][955] + xnor_result[9][956] + xnor_result[9][957] + xnor_result[9][958] + xnor_result[9][959] ;
logic [9:0] acc_store [0:9];

always @(posedge clk) begin
  acc_store <= accumulation_result;
end

assign accumulation_after_bias[0] = acc_store[0] - 9'd480;
assign accumulation_after_bias[1] = acc_store[1] - 9'd480;
assign accumulation_after_bias[2] = acc_store[2] - 9'd480;
assign accumulation_after_bias[3] = acc_store[3] - 9'd480;
assign accumulation_after_bias[4] = acc_store[4] - 9'd480;
assign accumulation_after_bias[5] = acc_store[5] - 9'd480;
assign accumulation_after_bias[6] = acc_store[6] - 9'd480;
assign accumulation_after_bias[7] = acc_store[7] - 9'd480;
assign accumulation_after_bias[8] = acc_store[8] - 9'd480;
assign accumulation_after_bias[9] = acc_store[9] - 9'd480;

logic [16:0] fan_result [0:9];
assign fan_result[0] = accumulation_after_bias[0][9] ? 17'd0 : (accumulation_after_bias[0][8:0] * weights[0]);
assign fan_result[1] = accumulation_after_bias[1][9] ? 17'd0 : (accumulation_after_bias[1][8:0] * weights[1]);
assign fan_result[2] = accumulation_after_bias[2][9] ? 17'd0 : (accumulation_after_bias[2][8:0] * weights[2]);
assign fan_result[3] = accumulation_after_bias[3][9] ? 17'd0 : (accumulation_after_bias[3][8:0] * weights[3]);
assign fan_result[4] = accumulation_after_bias[4][9] ? 17'd0 : (accumulation_after_bias[4][8:0] * weights[4]);
assign fan_result[5] = accumulation_after_bias[5][9] ? 17'd0 : (accumulation_after_bias[5][8:0] * weights[5]);
assign fan_result[6] = accumulation_after_bias[6][9] ? 17'd0 : (accumulation_after_bias[6][8:0] * weights[6]);
assign fan_result[7] = accumulation_after_bias[7][9] ? 17'd0 : (accumulation_after_bias[7][8:0] * weights[7]);
assign fan_result[8] = accumulation_after_bias[8][9] ? 17'd0 : (accumulation_after_bias[8][8:0] * weights[8]);
assign fan_result[9] = accumulation_after_bias[9][9] ? 17'd0 : (accumulation_after_bias[9][8:0] * weights[9]);


always @(posedge clk) begin
  fan_out <= fan_result;
end

endmodule









