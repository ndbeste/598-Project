module conv2
    #( parameter bW = 8 )
    (
    input  logic [0:18*12*12 -1]      image         ,
    input  logic [0:18*60*5*5-1]      kernels       ,
    output logic [0:18*60*8*8*bW-1]   xor_out 
    );

convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[1*5*5:2*5*5-1]), .o_out_fmap(xor_out[1*8*8*bW:2*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[2*5*5:3*5*5-1]), .o_out_fmap(xor_out[2*8*8*bW:3*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[3*5*5:4*5*5-1]), .o_out_fmap(xor_out[3*8*8*bW:4*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[4*5*5:5*5*5-1]), .o_out_fmap(xor_out[4*8*8*bW:5*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[5*5*5:6*5*5-1]), .o_out_fmap(xor_out[5*8*8*bW:6*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[6*5*5:7*5*5-1]), .o_out_fmap(xor_out[6*8*8*bW:7*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[7*5*5:8*5*5-1]), .o_out_fmap(xor_out[7*8*8*bW:8*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[8*5*5:9*5*5-1]), .o_out_fmap(xor_out[8*8*8*bW:9*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[9*5*5:10*5*5-1]), .o_out_fmap(xor_out[9*8*8*bW:10*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[10*5*5:11*5*5-1]), .o_out_fmap(xor_out[10*8*8*bW:11*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[11*5*5:12*5*5-1]), .o_out_fmap(xor_out[11*8*8*bW:12*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[12*5*5:13*5*5-1]), .o_out_fmap(xor_out[12*8*8*bW:13*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[13*5*5:14*5*5-1]), .o_out_fmap(xor_out[13*8*8*bW:14*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[14*5*5:15*5*5-1]), .o_out_fmap(xor_out[14*8*8*bW:15*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[15*5*5:16*5*5-1]), .o_out_fmap(xor_out[15*8*8*bW:16*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[16*5*5:17*5*5-1]), .o_out_fmap(xor_out[16*8*8*bW:17*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[17*5*5:18*5*5-1]), .o_out_fmap(xor_out[17*8*8*bW:18*8*8*bW-1]));
convchan2 c_2_18 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[18*5*5:19*5*5-1]), .o_out_fmap(xor_out[18*8*8*bW:19*8*8*bW-1]));
convchan2 c_2_19 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[19*5*5:20*5*5-1]), .o_out_fmap(xor_out[19*8*8*bW:20*8*8*bW-1]));
convchan2 c_2_20 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[20*5*5:21*5*5-1]), .o_out_fmap(xor_out[20*8*8*bW:21*8*8*bW-1]));
convchan2 c_2_21 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[21*5*5:22*5*5-1]), .o_out_fmap(xor_out[21*8*8*bW:22*8*8*bW-1]));
convchan2 c_2_22 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[22*5*5:23*5*5-1]), .o_out_fmap(xor_out[22*8*8*bW:23*8*8*bW-1]));
convchan2 c_2_23 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[23*5*5:24*5*5-1]), .o_out_fmap(xor_out[23*8*8*bW:24*8*8*bW-1]));
convchan2 c_2_24 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[24*5*5:25*5*5-1]), .o_out_fmap(xor_out[24*8*8*bW:25*8*8*bW-1]));
convchan2 c_2_25 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[25*5*5:26*5*5-1]), .o_out_fmap(xor_out[25*8*8*bW:26*8*8*bW-1]));
convchan2 c_2_26 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[26*5*5:27*5*5-1]), .o_out_fmap(xor_out[26*8*8*bW:27*8*8*bW-1]));
convchan2 c_2_27 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[27*5*5:28*5*5-1]), .o_out_fmap(xor_out[27*8*8*bW:28*8*8*bW-1]));
convchan2 c_2_28 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[28*5*5:29*5*5-1]), .o_out_fmap(xor_out[28*8*8*bW:29*8*8*bW-1]));
convchan2 c_2_29 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[29*5*5:30*5*5-1]), .o_out_fmap(xor_out[29*8*8*bW:30*8*8*bW-1]));
convchan2 c_2_30 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[30*5*5:31*5*5-1]), .o_out_fmap(xor_out[30*8*8*bW:31*8*8*bW-1]));
convchan2 c_2_31 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[31*5*5:32*5*5-1]), .o_out_fmap(xor_out[31*8*8*bW:32*8*8*bW-1]));
convchan2 c_2_32 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[32*5*5:33*5*5-1]), .o_out_fmap(xor_out[32*8*8*bW:33*8*8*bW-1]));
convchan2 c_2_33 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[33*5*5:34*5*5-1]), .o_out_fmap(xor_out[33*8*8*bW:34*8*8*bW-1]));
convchan2 c_2_34 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[34*5*5:35*5*5-1]), .o_out_fmap(xor_out[34*8*8*bW:35*8*8*bW-1]));
convchan2 c_2_35 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[35*5*5:36*5*5-1]), .o_out_fmap(xor_out[35*8*8*bW:36*8*8*bW-1]));
convchan2 c_2_36 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[36*5*5:37*5*5-1]), .o_out_fmap(xor_out[36*8*8*bW:37*8*8*bW-1]));
convchan2 c_2_37 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[37*5*5:38*5*5-1]), .o_out_fmap(xor_out[37*8*8*bW:38*8*8*bW-1]));
convchan2 c_2_38 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[38*5*5:39*5*5-1]), .o_out_fmap(xor_out[38*8*8*bW:39*8*8*bW-1]));
convchan2 c_2_39 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[39*5*5:40*5*5-1]), .o_out_fmap(xor_out[39*8*8*bW:40*8*8*bW-1]));
convchan2 c_2_40 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[40*5*5:41*5*5-1]), .o_out_fmap(xor_out[40*8*8*bW:41*8*8*bW-1]));
convchan2 c_2_41 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[41*5*5:42*5*5-1]), .o_out_fmap(xor_out[41*8*8*bW:42*8*8*bW-1]));
convchan2 c_2_42 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[42*5*5:43*5*5-1]), .o_out_fmap(xor_out[42*8*8*bW:43*8*8*bW-1]));
convchan2 c_2_43 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[43*5*5:44*5*5-1]), .o_out_fmap(xor_out[43*8*8*bW:44*8*8*bW-1]));
convchan2 c_2_44 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[44*5*5:45*5*5-1]), .o_out_fmap(xor_out[44*8*8*bW:45*8*8*bW-1]));
convchan2 c_2_45 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[45*5*5:46*5*5-1]), .o_out_fmap(xor_out[45*8*8*bW:46*8*8*bW-1]));
convchan2 c_2_46 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[46*5*5:47*5*5-1]), .o_out_fmap(xor_out[46*8*8*bW:47*8*8*bW-1]));
convchan2 c_2_47 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[47*5*5:48*5*5-1]), .o_out_fmap(xor_out[47*8*8*bW:48*8*8*bW-1]));
convchan2 c_2_48 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[48*5*5:49*5*5-1]), .o_out_fmap(xor_out[48*8*8*bW:49*8*8*bW-1]));
convchan2 c_2_49 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[49*5*5:50*5*5-1]), .o_out_fmap(xor_out[49*8*8*bW:50*8*8*bW-1]));
convchan2 c_2_50 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[50*5*5:51*5*5-1]), .o_out_fmap(xor_out[50*8*8*bW:51*8*8*bW-1]));
convchan2 c_2_51 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[51*5*5:52*5*5-1]), .o_out_fmap(xor_out[51*8*8*bW:52*8*8*bW-1]));
convchan2 c_2_52 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[52*5*5:53*5*5-1]), .o_out_fmap(xor_out[52*8*8*bW:53*8*8*bW-1]));
convchan2 c_2_53 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[53*5*5:54*5*5-1]), .o_out_fmap(xor_out[53*8*8*bW:54*8*8*bW-1]));
convchan2 c_2_54 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[54*5*5:55*5*5-1]), .o_out_fmap(xor_out[54*8*8*bW:55*8*8*bW-1]));
convchan2 c_2_55 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[55*5*5:56*5*5-1]), .o_out_fmap(xor_out[55*8*8*bW:56*8*8*bW-1]));
convchan2 c_2_56 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[56*5*5:57*5*5-1]), .o_out_fmap(xor_out[56*8*8*bW:57*8*8*bW-1]));
convchan2 c_2_57 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[57*5*5:58*5*5-1]), .o_out_fmap(xor_out[57*8*8*bW:58*8*8*bW-1]));
convchan2 c_2_58 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[58*5*5:59*5*5-1]), .o_out_fmap(xor_out[58*8*8*bW:59*8*8*bW-1]));
convchan2 c_2_59 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[59*5*5:60*5*5-1]), .o_out_fmap(xor_out[59*8*8*bW:60*8*8*bW-1]));
convchan2 c_2_60 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[60*5*5:61*5*5-1]), .o_out_fmap(xor_out[60*8*8*bW:61*8*8*bW-1]));
convchan2 c_2_61 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[61*5*5:62*5*5-1]), .o_out_fmap(xor_out[61*8*8*bW:62*8*8*bW-1]));
convchan2 c_2_62 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[62*5*5:63*5*5-1]), .o_out_fmap(xor_out[62*8*8*bW:63*8*8*bW-1]));
convchan2 c_2_63 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[63*5*5:64*5*5-1]), .o_out_fmap(xor_out[63*8*8*bW:64*8*8*bW-1]));
convchan2 c_2_64 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[64*5*5:65*5*5-1]), .o_out_fmap(xor_out[64*8*8*bW:65*8*8*bW-1]));
convchan2 c_2_65 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[65*5*5:66*5*5-1]), .o_out_fmap(xor_out[65*8*8*bW:66*8*8*bW-1]));
convchan2 c_2_66 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[66*5*5:67*5*5-1]), .o_out_fmap(xor_out[66*8*8*bW:67*8*8*bW-1]));
convchan2 c_2_67 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[67*5*5:68*5*5-1]), .o_out_fmap(xor_out[67*8*8*bW:68*8*8*bW-1]));
convchan2 c_2_68 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[68*5*5:69*5*5-1]), .o_out_fmap(xor_out[68*8*8*bW:69*8*8*bW-1]));
convchan2 c_2_69 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[69*5*5:70*5*5-1]), .o_out_fmap(xor_out[69*8*8*bW:70*8*8*bW-1]));
convchan2 c_2_70 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[70*5*5:71*5*5-1]), .o_out_fmap(xor_out[70*8*8*bW:71*8*8*bW-1]));
convchan2 c_2_71 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[71*5*5:72*5*5-1]), .o_out_fmap(xor_out[71*8*8*bW:72*8*8*bW-1]));
convchan2 c_2_72 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[72*5*5:73*5*5-1]), .o_out_fmap(xor_out[72*8*8*bW:73*8*8*bW-1]));
convchan2 c_2_73 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[73*5*5:74*5*5-1]), .o_out_fmap(xor_out[73*8*8*bW:74*8*8*bW-1]));
convchan2 c_2_74 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[74*5*5:75*5*5-1]), .o_out_fmap(xor_out[74*8*8*bW:75*8*8*bW-1]));
convchan2 c_2_75 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[75*5*5:76*5*5-1]), .o_out_fmap(xor_out[75*8*8*bW:76*8*8*bW-1]));
convchan2 c_2_76 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[76*5*5:77*5*5-1]), .o_out_fmap(xor_out[76*8*8*bW:77*8*8*bW-1]));
convchan2 c_2_77 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[77*5*5:78*5*5-1]), .o_out_fmap(xor_out[77*8*8*bW:78*8*8*bW-1]));
convchan2 c_2_78 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[78*5*5:79*5*5-1]), .o_out_fmap(xor_out[78*8*8*bW:79*8*8*bW-1]));
convchan2 c_2_79 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[79*5*5:80*5*5-1]), .o_out_fmap(xor_out[79*8*8*bW:80*8*8*bW-1]));
convchan2 c_2_80 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[80*5*5:81*5*5-1]), .o_out_fmap(xor_out[80*8*8*bW:81*8*8*bW-1]));
convchan2 c_2_81 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[81*5*5:82*5*5-1]), .o_out_fmap(xor_out[81*8*8*bW:82*8*8*bW-1]));
convchan2 c_2_82 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[82*5*5:83*5*5-1]), .o_out_fmap(xor_out[82*8*8*bW:83*8*8*bW-1]));
convchan2 c_2_83 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[83*5*5:84*5*5-1]), .o_out_fmap(xor_out[83*8*8*bW:84*8*8*bW-1]));
convchan2 c_2_84 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[84*5*5:85*5*5-1]), .o_out_fmap(xor_out[84*8*8*bW:85*8*8*bW-1]));
convchan2 c_2_85 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[85*5*5:86*5*5-1]), .o_out_fmap(xor_out[85*8*8*bW:86*8*8*bW-1]));
convchan2 c_2_86 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[86*5*5:87*5*5-1]), .o_out_fmap(xor_out[86*8*8*bW:87*8*8*bW-1]));
convchan2 c_2_87 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[87*5*5:88*5*5-1]), .o_out_fmap(xor_out[87*8*8*bW:88*8*8*bW-1]));
convchan2 c_2_88 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[88*5*5:89*5*5-1]), .o_out_fmap(xor_out[88*8*8*bW:89*8*8*bW-1]));
convchan2 c_2_89 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[89*5*5:90*5*5-1]), .o_out_fmap(xor_out[89*8*8*bW:90*8*8*bW-1]));
convchan2 c_2_90 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[90*5*5:91*5*5-1]), .o_out_fmap(xor_out[90*8*8*bW:91*8*8*bW-1]));
convchan2 c_2_91 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[91*5*5:92*5*5-1]), .o_out_fmap(xor_out[91*8*8*bW:92*8*8*bW-1]));
convchan2 c_2_92 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[92*5*5:93*5*5-1]), .o_out_fmap(xor_out[92*8*8*bW:93*8*8*bW-1]));
convchan2 c_2_93 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[93*5*5:94*5*5-1]), .o_out_fmap(xor_out[93*8*8*bW:94*8*8*bW-1]));
convchan2 c_2_94 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[94*5*5:95*5*5-1]), .o_out_fmap(xor_out[94*8*8*bW:95*8*8*bW-1]));
convchan2 c_2_95 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[95*5*5:96*5*5-1]), .o_out_fmap(xor_out[95*8*8*bW:96*8*8*bW-1]));
convchan2 c_2_96 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[96*5*5:97*5*5-1]), .o_out_fmap(xor_out[96*8*8*bW:97*8*8*bW-1]));
convchan2 c_2_97 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[97*5*5:98*5*5-1]), .o_out_fmap(xor_out[97*8*8*bW:98*8*8*bW-1]));
convchan2 c_2_98 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[98*5*5:99*5*5-1]), .o_out_fmap(xor_out[98*8*8*bW:99*8*8*bW-1]));
convchan2 c_2_99 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[99*5*5:100*5*5-1]), .o_out_fmap(xor_out[99*8*8*bW:100*8*8*bW-1]));
convchan2 c_2_100 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[100*5*5:101*5*5-1]), .o_out_fmap(xor_out[100*8*8*bW:101*8*8*bW-1]));
convchan2 c_2_101 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[101*5*5:102*5*5-1]), .o_out_fmap(xor_out[101*8*8*bW:102*8*8*bW-1]));
convchan2 c_2_102 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[102*5*5:103*5*5-1]), .o_out_fmap(xor_out[102*8*8*bW:103*8*8*bW-1]));
convchan2 c_2_103 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[103*5*5:104*5*5-1]), .o_out_fmap(xor_out[103*8*8*bW:104*8*8*bW-1]));
convchan2 c_2_104 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[104*5*5:105*5*5-1]), .o_out_fmap(xor_out[104*8*8*bW:105*8*8*bW-1]));
convchan2 c_2_105 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[105*5*5:106*5*5-1]), .o_out_fmap(xor_out[105*8*8*bW:106*8*8*bW-1]));
convchan2 c_2_106 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[106*5*5:107*5*5-1]), .o_out_fmap(xor_out[106*8*8*bW:107*8*8*bW-1]));
convchan2 c_2_107 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[107*5*5:108*5*5-1]), .o_out_fmap(xor_out[107*8*8*bW:108*8*8*bW-1]));
convchan2 c_2_108 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[108*5*5:109*5*5-1]), .o_out_fmap(xor_out[108*8*8*bW:109*8*8*bW-1]));
convchan2 c_2_109 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[109*5*5:110*5*5-1]), .o_out_fmap(xor_out[109*8*8*bW:110*8*8*bW-1]));
convchan2 c_2_110 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[110*5*5:111*5*5-1]), .o_out_fmap(xor_out[110*8*8*bW:111*8*8*bW-1]));
convchan2 c_2_111 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[111*5*5:112*5*5-1]), .o_out_fmap(xor_out[111*8*8*bW:112*8*8*bW-1]));
convchan2 c_2_112 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[112*5*5:113*5*5-1]), .o_out_fmap(xor_out[112*8*8*bW:113*8*8*bW-1]));
convchan2 c_2_113 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[113*5*5:114*5*5-1]), .o_out_fmap(xor_out[113*8*8*bW:114*8*8*bW-1]));
convchan2 c_2_114 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[114*5*5:115*5*5-1]), .o_out_fmap(xor_out[114*8*8*bW:115*8*8*bW-1]));
convchan2 c_2_115 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[115*5*5:116*5*5-1]), .o_out_fmap(xor_out[115*8*8*bW:116*8*8*bW-1]));
convchan2 c_2_116 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[116*5*5:117*5*5-1]), .o_out_fmap(xor_out[116*8*8*bW:117*8*8*bW-1]));
convchan2 c_2_117 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[117*5*5:118*5*5-1]), .o_out_fmap(xor_out[117*8*8*bW:118*8*8*bW-1]));
convchan2 c_2_118 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[118*5*5:119*5*5-1]), .o_out_fmap(xor_out[118*8*8*bW:119*8*8*bW-1]));
convchan2 c_2_119 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[119*5*5:120*5*5-1]), .o_out_fmap(xor_out[119*8*8*bW:120*8*8*bW-1]));
convchan2 c_2_120 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[120*5*5:121*5*5-1]), .o_out_fmap(xor_out[120*8*8*bW:121*8*8*bW-1]));
convchan2 c_2_121 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[121*5*5:122*5*5-1]), .o_out_fmap(xor_out[121*8*8*bW:122*8*8*bW-1]));
convchan2 c_2_122 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[122*5*5:123*5*5-1]), .o_out_fmap(xor_out[122*8*8*bW:123*8*8*bW-1]));
convchan2 c_2_123 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[123*5*5:124*5*5-1]), .o_out_fmap(xor_out[123*8*8*bW:124*8*8*bW-1]));
convchan2 c_2_124 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[124*5*5:125*5*5-1]), .o_out_fmap(xor_out[124*8*8*bW:125*8*8*bW-1]));
convchan2 c_2_125 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[125*5*5:126*5*5-1]), .o_out_fmap(xor_out[125*8*8*bW:126*8*8*bW-1]));
convchan2 c_2_126 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[126*5*5:127*5*5-1]), .o_out_fmap(xor_out[126*8*8*bW:127*8*8*bW-1]));
convchan2 c_2_127 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[127*5*5:128*5*5-1]), .o_out_fmap(xor_out[127*8*8*bW:128*8*8*bW-1]));
convchan2 c_2_128 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[128*5*5:129*5*5-1]), .o_out_fmap(xor_out[128*8*8*bW:129*8*8*bW-1]));
convchan2 c_2_129 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[129*5*5:130*5*5-1]), .o_out_fmap(xor_out[129*8*8*bW:130*8*8*bW-1]));
convchan2 c_2_130 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[130*5*5:131*5*5-1]), .o_out_fmap(xor_out[130*8*8*bW:131*8*8*bW-1]));
convchan2 c_2_131 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[131*5*5:132*5*5-1]), .o_out_fmap(xor_out[131*8*8*bW:132*8*8*bW-1]));
convchan2 c_2_132 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[132*5*5:133*5*5-1]), .o_out_fmap(xor_out[132*8*8*bW:133*8*8*bW-1]));
convchan2 c_2_133 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[133*5*5:134*5*5-1]), .o_out_fmap(xor_out[133*8*8*bW:134*8*8*bW-1]));
convchan2 c_2_134 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[134*5*5:135*5*5-1]), .o_out_fmap(xor_out[134*8*8*bW:135*8*8*bW-1]));
convchan2 c_2_135 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[135*5*5:136*5*5-1]), .o_out_fmap(xor_out[135*8*8*bW:136*8*8*bW-1]));
convchan2 c_2_136 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[136*5*5:137*5*5-1]), .o_out_fmap(xor_out[136*8*8*bW:137*8*8*bW-1]));
convchan2 c_2_137 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[137*5*5:138*5*5-1]), .o_out_fmap(xor_out[137*8*8*bW:138*8*8*bW-1]));
convchan2 c_2_138 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[138*5*5:139*5*5-1]), .o_out_fmap(xor_out[138*8*8*bW:139*8*8*bW-1]));
convchan2 c_2_139 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[139*5*5:140*5*5-1]), .o_out_fmap(xor_out[139*8*8*bW:140*8*8*bW-1]));
convchan2 c_2_140 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[140*5*5:141*5*5-1]), .o_out_fmap(xor_out[140*8*8*bW:141*8*8*bW-1]));
convchan2 c_2_141 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[141*5*5:142*5*5-1]), .o_out_fmap(xor_out[141*8*8*bW:142*8*8*bW-1]));
convchan2 c_2_142 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[142*5*5:143*5*5-1]), .o_out_fmap(xor_out[142*8*8*bW:143*8*8*bW-1]));
convchan2 c_2_143 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[143*5*5:144*5*5-1]), .o_out_fmap(xor_out[143*8*8*bW:144*8*8*bW-1]));
convchan2 c_2_144 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[144*5*5:145*5*5-1]), .o_out_fmap(xor_out[144*8*8*bW:145*8*8*bW-1]));
convchan2 c_2_145 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[145*5*5:146*5*5-1]), .o_out_fmap(xor_out[145*8*8*bW:146*8*8*bW-1]));
convchan2 c_2_146 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[146*5*5:147*5*5-1]), .o_out_fmap(xor_out[146*8*8*bW:147*8*8*bW-1]));
convchan2 c_2_147 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[147*5*5:148*5*5-1]), .o_out_fmap(xor_out[147*8*8*bW:148*8*8*bW-1]));
convchan2 c_2_148 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[148*5*5:149*5*5-1]), .o_out_fmap(xor_out[148*8*8*bW:149*8*8*bW-1]));
convchan2 c_2_149 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[149*5*5:150*5*5-1]), .o_out_fmap(xor_out[149*8*8*bW:150*8*8*bW-1]));
convchan2 c_2_150 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[150*5*5:151*5*5-1]), .o_out_fmap(xor_out[150*8*8*bW:151*8*8*bW-1]));
convchan2 c_2_151 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[151*5*5:152*5*5-1]), .o_out_fmap(xor_out[151*8*8*bW:152*8*8*bW-1]));
convchan2 c_2_152 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[152*5*5:153*5*5-1]), .o_out_fmap(xor_out[152*8*8*bW:153*8*8*bW-1]));
convchan2 c_2_153 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[153*5*5:154*5*5-1]), .o_out_fmap(xor_out[153*8*8*bW:154*8*8*bW-1]));
convchan2 c_2_154 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[154*5*5:155*5*5-1]), .o_out_fmap(xor_out[154*8*8*bW:155*8*8*bW-1]));
convchan2 c_2_155 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[155*5*5:156*5*5-1]), .o_out_fmap(xor_out[155*8*8*bW:156*8*8*bW-1]));
convchan2 c_2_156 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[156*5*5:157*5*5-1]), .o_out_fmap(xor_out[156*8*8*bW:157*8*8*bW-1]));
convchan2 c_2_157 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[157*5*5:158*5*5-1]), .o_out_fmap(xor_out[157*8*8*bW:158*8*8*bW-1]));
convchan2 c_2_158 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[158*5*5:159*5*5-1]), .o_out_fmap(xor_out[158*8*8*bW:159*8*8*bW-1]));
convchan2 c_2_159 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[159*5*5:160*5*5-1]), .o_out_fmap(xor_out[159*8*8*bW:160*8*8*bW-1]));
convchan2 c_2_160 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[160*5*5:161*5*5-1]), .o_out_fmap(xor_out[160*8*8*bW:161*8*8*bW-1]));
convchan2 c_2_161 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[161*5*5:162*5*5-1]), .o_out_fmap(xor_out[161*8*8*bW:162*8*8*bW-1]));
convchan2 c_2_162 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[162*5*5:163*5*5-1]), .o_out_fmap(xor_out[162*8*8*bW:163*8*8*bW-1]));
convchan2 c_2_163 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[163*5*5:164*5*5-1]), .o_out_fmap(xor_out[163*8*8*bW:164*8*8*bW-1]));
convchan2 c_2_164 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[164*5*5:165*5*5-1]), .o_out_fmap(xor_out[164*8*8*bW:165*8*8*bW-1]));
convchan2 c_2_165 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[165*5*5:166*5*5-1]), .o_out_fmap(xor_out[165*8*8*bW:166*8*8*bW-1]));
convchan2 c_2_166 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[166*5*5:167*5*5-1]), .o_out_fmap(xor_out[166*8*8*bW:167*8*8*bW-1]));
convchan2 c_2_167 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[167*5*5:168*5*5-1]), .o_out_fmap(xor_out[167*8*8*bW:168*8*8*bW-1]));
convchan2 c_2_168 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[168*5*5:169*5*5-1]), .o_out_fmap(xor_out[168*8*8*bW:169*8*8*bW-1]));
convchan2 c_2_169 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[169*5*5:170*5*5-1]), .o_out_fmap(xor_out[169*8*8*bW:170*8*8*bW-1]));
convchan2 c_2_170 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[170*5*5:171*5*5-1]), .o_out_fmap(xor_out[170*8*8*bW:171*8*8*bW-1]));
convchan2 c_2_171 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[171*5*5:172*5*5-1]), .o_out_fmap(xor_out[171*8*8*bW:172*8*8*bW-1]));
convchan2 c_2_172 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[172*5*5:173*5*5-1]), .o_out_fmap(xor_out[172*8*8*bW:173*8*8*bW-1]));
convchan2 c_2_173 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[173*5*5:174*5*5-1]), .o_out_fmap(xor_out[173*8*8*bW:174*8*8*bW-1]));
convchan2 c_2_174 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[174*5*5:175*5*5-1]), .o_out_fmap(xor_out[174*8*8*bW:175*8*8*bW-1]));
convchan2 c_2_175 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[175*5*5:176*5*5-1]), .o_out_fmap(xor_out[175*8*8*bW:176*8*8*bW-1]));
convchan2 c_2_176 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[176*5*5:177*5*5-1]), .o_out_fmap(xor_out[176*8*8*bW:177*8*8*bW-1]));
convchan2 c_2_177 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[177*5*5:178*5*5-1]), .o_out_fmap(xor_out[177*8*8*bW:178*8*8*bW-1]));
convchan2 c_2_178 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[178*5*5:179*5*5-1]), .o_out_fmap(xor_out[178*8*8*bW:179*8*8*bW-1]));
convchan2 c_2_179 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[179*5*5:180*5*5-1]), .o_out_fmap(xor_out[179*8*8*bW:180*8*8*bW-1]));
convchan2 c_2_180 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[180*5*5:181*5*5-1]), .o_out_fmap(xor_out[180*8*8*bW:181*8*8*bW-1]));
convchan2 c_2_181 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[181*5*5:182*5*5-1]), .o_out_fmap(xor_out[181*8*8*bW:182*8*8*bW-1]));
convchan2 c_2_182 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[182*5*5:183*5*5-1]), .o_out_fmap(xor_out[182*8*8*bW:183*8*8*bW-1]));
convchan2 c_2_183 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[183*5*5:184*5*5-1]), .o_out_fmap(xor_out[183*8*8*bW:184*8*8*bW-1]));
convchan2 c_2_184 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[184*5*5:185*5*5-1]), .o_out_fmap(xor_out[184*8*8*bW:185*8*8*bW-1]));
convchan2 c_2_185 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[185*5*5:186*5*5-1]), .o_out_fmap(xor_out[185*8*8*bW:186*8*8*bW-1]));
convchan2 c_2_186 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[186*5*5:187*5*5-1]), .o_out_fmap(xor_out[186*8*8*bW:187*8*8*bW-1]));
convchan2 c_2_187 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[187*5*5:188*5*5-1]), .o_out_fmap(xor_out[187*8*8*bW:188*8*8*bW-1]));
convchan2 c_2_188 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[188*5*5:189*5*5-1]), .o_out_fmap(xor_out[188*8*8*bW:189*8*8*bW-1]));
convchan2 c_2_189 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[189*5*5:190*5*5-1]), .o_out_fmap(xor_out[189*8*8*bW:190*8*8*bW-1]));
convchan2 c_2_190 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[190*5*5:191*5*5-1]), .o_out_fmap(xor_out[190*8*8*bW:191*8*8*bW-1]));
convchan2 c_2_191 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[191*5*5:192*5*5-1]), .o_out_fmap(xor_out[191*8*8*bW:192*8*8*bW-1]));
convchan2 c_2_192 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[192*5*5:193*5*5-1]), .o_out_fmap(xor_out[192*8*8*bW:193*8*8*bW-1]));
convchan2 c_2_193 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[193*5*5:194*5*5-1]), .o_out_fmap(xor_out[193*8*8*bW:194*8*8*bW-1]));
convchan2 c_2_194 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[194*5*5:195*5*5-1]), .o_out_fmap(xor_out[194*8*8*bW:195*8*8*bW-1]));
convchan2 c_2_195 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[195*5*5:196*5*5-1]), .o_out_fmap(xor_out[195*8*8*bW:196*8*8*bW-1]));
convchan2 c_2_196 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[196*5*5:197*5*5-1]), .o_out_fmap(xor_out[196*8*8*bW:197*8*8*bW-1]));
convchan2 c_2_197 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[197*5*5:198*5*5-1]), .o_out_fmap(xor_out[197*8*8*bW:198*8*8*bW-1]));
convchan2 c_2_198 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[198*5*5:199*5*5-1]), .o_out_fmap(xor_out[198*8*8*bW:199*8*8*bW-1]));
convchan2 c_2_199 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[199*5*5:200*5*5-1]), .o_out_fmap(xor_out[199*8*8*bW:200*8*8*bW-1]));
convchan2 c_2_200 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[200*5*5:201*5*5-1]), .o_out_fmap(xor_out[200*8*8*bW:201*8*8*bW-1]));
convchan2 c_2_201 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[201*5*5:202*5*5-1]), .o_out_fmap(xor_out[201*8*8*bW:202*8*8*bW-1]));
convchan2 c_2_202 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[202*5*5:203*5*5-1]), .o_out_fmap(xor_out[202*8*8*bW:203*8*8*bW-1]));
convchan2 c_2_203 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[203*5*5:204*5*5-1]), .o_out_fmap(xor_out[203*8*8*bW:204*8*8*bW-1]));
convchan2 c_2_204 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[204*5*5:205*5*5-1]), .o_out_fmap(xor_out[204*8*8*bW:205*8*8*bW-1]));
convchan2 c_2_205 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[205*5*5:206*5*5-1]), .o_out_fmap(xor_out[205*8*8*bW:206*8*8*bW-1]));
convchan2 c_2_206 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[206*5*5:207*5*5-1]), .o_out_fmap(xor_out[206*8*8*bW:207*8*8*bW-1]));
convchan2 c_2_207 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[207*5*5:208*5*5-1]), .o_out_fmap(xor_out[207*8*8*bW:208*8*8*bW-1]));
convchan2 c_2_208 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[208*5*5:209*5*5-1]), .o_out_fmap(xor_out[208*8*8*bW:209*8*8*bW-1]));
convchan2 c_2_209 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[209*5*5:210*5*5-1]), .o_out_fmap(xor_out[209*8*8*bW:210*8*8*bW-1]));
convchan2 c_2_210 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[210*5*5:211*5*5-1]), .o_out_fmap(xor_out[210*8*8*bW:211*8*8*bW-1]));
convchan2 c_2_211 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[211*5*5:212*5*5-1]), .o_out_fmap(xor_out[211*8*8*bW:212*8*8*bW-1]));
convchan2 c_2_212 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[212*5*5:213*5*5-1]), .o_out_fmap(xor_out[212*8*8*bW:213*8*8*bW-1]));
convchan2 c_2_213 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[213*5*5:214*5*5-1]), .o_out_fmap(xor_out[213*8*8*bW:214*8*8*bW-1]));
convchan2 c_2_214 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[214*5*5:215*5*5-1]), .o_out_fmap(xor_out[214*8*8*bW:215*8*8*bW-1]));
convchan2 c_2_215 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[215*5*5:216*5*5-1]), .o_out_fmap(xor_out[215*8*8*bW:216*8*8*bW-1]));
convchan2 c_2_216 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[216*5*5:217*5*5-1]), .o_out_fmap(xor_out[216*8*8*bW:217*8*8*bW-1]));
convchan2 c_2_217 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[217*5*5:218*5*5-1]), .o_out_fmap(xor_out[217*8*8*bW:218*8*8*bW-1]));
convchan2 c_2_218 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[218*5*5:219*5*5-1]), .o_out_fmap(xor_out[218*8*8*bW:219*8*8*bW-1]));
convchan2 c_2_219 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[219*5*5:220*5*5-1]), .o_out_fmap(xor_out[219*8*8*bW:220*8*8*bW-1]));
convchan2 c_2_220 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[220*5*5:221*5*5-1]), .o_out_fmap(xor_out[220*8*8*bW:221*8*8*bW-1]));
convchan2 c_2_221 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[221*5*5:222*5*5-1]), .o_out_fmap(xor_out[221*8*8*bW:222*8*8*bW-1]));
convchan2 c_2_222 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[222*5*5:223*5*5-1]), .o_out_fmap(xor_out[222*8*8*bW:223*8*8*bW-1]));
convchan2 c_2_223 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[223*5*5:224*5*5-1]), .o_out_fmap(xor_out[223*8*8*bW:224*8*8*bW-1]));
convchan2 c_2_224 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[224*5*5:225*5*5-1]), .o_out_fmap(xor_out[224*8*8*bW:225*8*8*bW-1]));
convchan2 c_2_225 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[225*5*5:226*5*5-1]), .o_out_fmap(xor_out[225*8*8*bW:226*8*8*bW-1]));
convchan2 c_2_226 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[226*5*5:227*5*5-1]), .o_out_fmap(xor_out[226*8*8*bW:227*8*8*bW-1]));
convchan2 c_2_227 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[227*5*5:228*5*5-1]), .o_out_fmap(xor_out[227*8*8*bW:228*8*8*bW-1]));
convchan2 c_2_228 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[228*5*5:229*5*5-1]), .o_out_fmap(xor_out[228*8*8*bW:229*8*8*bW-1]));
convchan2 c_2_229 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[229*5*5:230*5*5-1]), .o_out_fmap(xor_out[229*8*8*bW:230*8*8*bW-1]));
convchan2 c_2_230 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[230*5*5:231*5*5-1]), .o_out_fmap(xor_out[230*8*8*bW:231*8*8*bW-1]));
convchan2 c_2_231 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[231*5*5:232*5*5-1]), .o_out_fmap(xor_out[231*8*8*bW:232*8*8*bW-1]));
convchan2 c_2_232 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[232*5*5:233*5*5-1]), .o_out_fmap(xor_out[232*8*8*bW:233*8*8*bW-1]));
convchan2 c_2_233 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[233*5*5:234*5*5-1]), .o_out_fmap(xor_out[233*8*8*bW:234*8*8*bW-1]));
convchan2 c_2_234 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[234*5*5:235*5*5-1]), .o_out_fmap(xor_out[234*8*8*bW:235*8*8*bW-1]));
convchan2 c_2_235 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[235*5*5:236*5*5-1]), .o_out_fmap(xor_out[235*8*8*bW:236*8*8*bW-1]));
convchan2 c_2_236 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[236*5*5:237*5*5-1]), .o_out_fmap(xor_out[236*8*8*bW:237*8*8*bW-1]));
convchan2 c_2_237 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[237*5*5:238*5*5-1]), .o_out_fmap(xor_out[237*8*8*bW:238*8*8*bW-1]));
convchan2 c_2_238 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[238*5*5:239*5*5-1]), .o_out_fmap(xor_out[238*8*8*bW:239*8*8*bW-1]));
convchan2 c_2_239 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[239*5*5:240*5*5-1]), .o_out_fmap(xor_out[239*8*8*bW:240*8*8*bW-1]));
convchan2 c_2_240 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[240*5*5:241*5*5-1]), .o_out_fmap(xor_out[240*8*8*bW:241*8*8*bW-1]));
convchan2 c_2_241 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[241*5*5:242*5*5-1]), .o_out_fmap(xor_out[241*8*8*bW:242*8*8*bW-1]));
convchan2 c_2_242 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[242*5*5:243*5*5-1]), .o_out_fmap(xor_out[242*8*8*bW:243*8*8*bW-1]));
convchan2 c_2_243 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[243*5*5:244*5*5-1]), .o_out_fmap(xor_out[243*8*8*bW:244*8*8*bW-1]));
convchan2 c_2_244 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[244*5*5:245*5*5-1]), .o_out_fmap(xor_out[244*8*8*bW:245*8*8*bW-1]));
convchan2 c_2_245 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[245*5*5:246*5*5-1]), .o_out_fmap(xor_out[245*8*8*bW:246*8*8*bW-1]));
convchan2 c_2_246 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[246*5*5:247*5*5-1]), .o_out_fmap(xor_out[246*8*8*bW:247*8*8*bW-1]));
convchan2 c_2_247 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[247*5*5:248*5*5-1]), .o_out_fmap(xor_out[247*8*8*bW:248*8*8*bW-1]));
convchan2 c_2_248 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[248*5*5:249*5*5-1]), .o_out_fmap(xor_out[248*8*8*bW:249*8*8*bW-1]));
convchan2 c_2_249 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[249*5*5:250*5*5-1]), .o_out_fmap(xor_out[249*8*8*bW:250*8*8*bW-1]));
convchan2 c_2_250 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[250*5*5:251*5*5-1]), .o_out_fmap(xor_out[250*8*8*bW:251*8*8*bW-1]));
convchan2 c_2_251 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[251*5*5:252*5*5-1]), .o_out_fmap(xor_out[251*8*8*bW:252*8*8*bW-1]));
convchan2 c_2_252 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[252*5*5:253*5*5-1]), .o_out_fmap(xor_out[252*8*8*bW:253*8*8*bW-1]));
convchan2 c_2_253 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[253*5*5:254*5*5-1]), .o_out_fmap(xor_out[253*8*8*bW:254*8*8*bW-1]));
convchan2 c_2_254 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[254*5*5:255*5*5-1]), .o_out_fmap(xor_out[254*8*8*bW:255*8*8*bW-1]));
convchan2 c_2_255 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[255*5*5:256*5*5-1]), .o_out_fmap(xor_out[255*8*8*bW:256*8*8*bW-1]));
convchan2 c_2_256 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[256*5*5:257*5*5-1]), .o_out_fmap(xor_out[256*8*8*bW:257*8*8*bW-1]));
convchan2 c_2_257 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[257*5*5:258*5*5-1]), .o_out_fmap(xor_out[257*8*8*bW:258*8*8*bW-1]));
convchan2 c_2_258 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[258*5*5:259*5*5-1]), .o_out_fmap(xor_out[258*8*8*bW:259*8*8*bW-1]));
convchan2 c_2_259 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[259*5*5:260*5*5-1]), .o_out_fmap(xor_out[259*8*8*bW:260*8*8*bW-1]));
convchan2 c_2_260 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[260*5*5:261*5*5-1]), .o_out_fmap(xor_out[260*8*8*bW:261*8*8*bW-1]));
convchan2 c_2_261 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[261*5*5:262*5*5-1]), .o_out_fmap(xor_out[261*8*8*bW:262*8*8*bW-1]));
convchan2 c_2_262 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[262*5*5:263*5*5-1]), .o_out_fmap(xor_out[262*8*8*bW:263*8*8*bW-1]));
convchan2 c_2_263 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[263*5*5:264*5*5-1]), .o_out_fmap(xor_out[263*8*8*bW:264*8*8*bW-1]));
convchan2 c_2_264 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[264*5*5:265*5*5-1]), .o_out_fmap(xor_out[264*8*8*bW:265*8*8*bW-1]));
convchan2 c_2_265 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[265*5*5:266*5*5-1]), .o_out_fmap(xor_out[265*8*8*bW:266*8*8*bW-1]));
convchan2 c_2_266 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[266*5*5:267*5*5-1]), .o_out_fmap(xor_out[266*8*8*bW:267*8*8*bW-1]));
convchan2 c_2_267 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[267*5*5:268*5*5-1]), .o_out_fmap(xor_out[267*8*8*bW:268*8*8*bW-1]));
convchan2 c_2_268 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[268*5*5:269*5*5-1]), .o_out_fmap(xor_out[268*8*8*bW:269*8*8*bW-1]));
convchan2 c_2_269 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[269*5*5:270*5*5-1]), .o_out_fmap(xor_out[269*8*8*bW:270*8*8*bW-1]));
convchan2 c_2_270 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[270*5*5:271*5*5-1]), .o_out_fmap(xor_out[270*8*8*bW:271*8*8*bW-1]));
convchan2 c_2_271 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[271*5*5:272*5*5-1]), .o_out_fmap(xor_out[271*8*8*bW:272*8*8*bW-1]));
convchan2 c_2_272 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[272*5*5:273*5*5-1]), .o_out_fmap(xor_out[272*8*8*bW:273*8*8*bW-1]));
convchan2 c_2_273 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[273*5*5:274*5*5-1]), .o_out_fmap(xor_out[273*8*8*bW:274*8*8*bW-1]));
convchan2 c_2_274 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[274*5*5:275*5*5-1]), .o_out_fmap(xor_out[274*8*8*bW:275*8*8*bW-1]));
convchan2 c_2_275 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[275*5*5:276*5*5-1]), .o_out_fmap(xor_out[275*8*8*bW:276*8*8*bW-1]));
convchan2 c_2_276 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[276*5*5:277*5*5-1]), .o_out_fmap(xor_out[276*8*8*bW:277*8*8*bW-1]));
convchan2 c_2_277 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[277*5*5:278*5*5-1]), .o_out_fmap(xor_out[277*8*8*bW:278*8*8*bW-1]));
convchan2 c_2_278 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[278*5*5:279*5*5-1]), .o_out_fmap(xor_out[278*8*8*bW:279*8*8*bW-1]));
convchan2 c_2_279 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[279*5*5:280*5*5-1]), .o_out_fmap(xor_out[279*8*8*bW:280*8*8*bW-1]));
convchan2 c_2_280 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[280*5*5:281*5*5-1]), .o_out_fmap(xor_out[280*8*8*bW:281*8*8*bW-1]));
convchan2 c_2_281 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[281*5*5:282*5*5-1]), .o_out_fmap(xor_out[281*8*8*bW:282*8*8*bW-1]));
convchan2 c_2_282 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[282*5*5:283*5*5-1]), .o_out_fmap(xor_out[282*8*8*bW:283*8*8*bW-1]));
convchan2 c_2_283 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[283*5*5:284*5*5-1]), .o_out_fmap(xor_out[283*8*8*bW:284*8*8*bW-1]));
convchan2 c_2_284 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[284*5*5:285*5*5-1]), .o_out_fmap(xor_out[284*8*8*bW:285*8*8*bW-1]));
convchan2 c_2_285 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[285*5*5:286*5*5-1]), .o_out_fmap(xor_out[285*8*8*bW:286*8*8*bW-1]));
convchan2 c_2_286 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[286*5*5:287*5*5-1]), .o_out_fmap(xor_out[286*8*8*bW:287*8*8*bW-1]));
convchan2 c_2_287 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[287*5*5:288*5*5-1]), .o_out_fmap(xor_out[287*8*8*bW:288*8*8*bW-1]));
convchan2 c_2_288 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[288*5*5:289*5*5-1]), .o_out_fmap(xor_out[288*8*8*bW:289*8*8*bW-1]));
convchan2 c_2_289 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[289*5*5:290*5*5-1]), .o_out_fmap(xor_out[289*8*8*bW:290*8*8*bW-1]));
convchan2 c_2_290 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[290*5*5:291*5*5-1]), .o_out_fmap(xor_out[290*8*8*bW:291*8*8*bW-1]));
convchan2 c_2_291 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[291*5*5:292*5*5-1]), .o_out_fmap(xor_out[291*8*8*bW:292*8*8*bW-1]));
convchan2 c_2_292 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[292*5*5:293*5*5-1]), .o_out_fmap(xor_out[292*8*8*bW:293*8*8*bW-1]));
convchan2 c_2_293 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[293*5*5:294*5*5-1]), .o_out_fmap(xor_out[293*8*8*bW:294*8*8*bW-1]));
convchan2 c_2_294 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[294*5*5:295*5*5-1]), .o_out_fmap(xor_out[294*8*8*bW:295*8*8*bW-1]));
convchan2 c_2_295 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[295*5*5:296*5*5-1]), .o_out_fmap(xor_out[295*8*8*bW:296*8*8*bW-1]));
convchan2 c_2_296 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[296*5*5:297*5*5-1]), .o_out_fmap(xor_out[296*8*8*bW:297*8*8*bW-1]));
convchan2 c_2_297 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[297*5*5:298*5*5-1]), .o_out_fmap(xor_out[297*8*8*bW:298*8*8*bW-1]));
convchan2 c_2_298 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[298*5*5:299*5*5-1]), .o_out_fmap(xor_out[298*8*8*bW:299*8*8*bW-1]));
convchan2 c_2_299 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[299*5*5:300*5*5-1]), .o_out_fmap(xor_out[299*8*8*bW:300*8*8*bW-1]));
convchan2 c_2_300 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[300*5*5:301*5*5-1]), .o_out_fmap(xor_out[300*8*8*bW:301*8*8*bW-1]));
convchan2 c_2_301 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[301*5*5:302*5*5-1]), .o_out_fmap(xor_out[301*8*8*bW:302*8*8*bW-1]));
convchan2 c_2_302 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[302*5*5:303*5*5-1]), .o_out_fmap(xor_out[302*8*8*bW:303*8*8*bW-1]));
convchan2 c_2_303 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[303*5*5:304*5*5-1]), .o_out_fmap(xor_out[303*8*8*bW:304*8*8*bW-1]));
convchan2 c_2_304 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[304*5*5:305*5*5-1]), .o_out_fmap(xor_out[304*8*8*bW:305*8*8*bW-1]));
convchan2 c_2_305 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[305*5*5:306*5*5-1]), .o_out_fmap(xor_out[305*8*8*bW:306*8*8*bW-1]));
convchan2 c_2_306 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[306*5*5:307*5*5-1]), .o_out_fmap(xor_out[306*8*8*bW:307*8*8*bW-1]));
convchan2 c_2_307 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[307*5*5:308*5*5-1]), .o_out_fmap(xor_out[307*8*8*bW:308*8*8*bW-1]));
convchan2 c_2_308 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[308*5*5:309*5*5-1]), .o_out_fmap(xor_out[308*8*8*bW:309*8*8*bW-1]));
convchan2 c_2_309 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[309*5*5:310*5*5-1]), .o_out_fmap(xor_out[309*8*8*bW:310*8*8*bW-1]));
convchan2 c_2_310 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[310*5*5:311*5*5-1]), .o_out_fmap(xor_out[310*8*8*bW:311*8*8*bW-1]));
convchan2 c_2_311 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[311*5*5:312*5*5-1]), .o_out_fmap(xor_out[311*8*8*bW:312*8*8*bW-1]));
convchan2 c_2_312 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[312*5*5:313*5*5-1]), .o_out_fmap(xor_out[312*8*8*bW:313*8*8*bW-1]));
convchan2 c_2_313 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[313*5*5:314*5*5-1]), .o_out_fmap(xor_out[313*8*8*bW:314*8*8*bW-1]));
convchan2 c_2_314 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[314*5*5:315*5*5-1]), .o_out_fmap(xor_out[314*8*8*bW:315*8*8*bW-1]));
convchan2 c_2_315 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[315*5*5:316*5*5-1]), .o_out_fmap(xor_out[315*8*8*bW:316*8*8*bW-1]));
convchan2 c_2_316 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[316*5*5:317*5*5-1]), .o_out_fmap(xor_out[316*8*8*bW:317*8*8*bW-1]));
convchan2 c_2_317 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[317*5*5:318*5*5-1]), .o_out_fmap(xor_out[317*8*8*bW:318*8*8*bW-1]));
convchan2 c_2_318 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[318*5*5:319*5*5-1]), .o_out_fmap(xor_out[318*8*8*bW:319*8*8*bW-1]));
convchan2 c_2_319 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[319*5*5:320*5*5-1]), .o_out_fmap(xor_out[319*8*8*bW:320*8*8*bW-1]));
convchan2 c_2_320 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[320*5*5:321*5*5-1]), .o_out_fmap(xor_out[320*8*8*bW:321*8*8*bW-1]));
convchan2 c_2_321 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[321*5*5:322*5*5-1]), .o_out_fmap(xor_out[321*8*8*bW:322*8*8*bW-1]));
convchan2 c_2_322 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[322*5*5:323*5*5-1]), .o_out_fmap(xor_out[322*8*8*bW:323*8*8*bW-1]));
convchan2 c_2_323 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[323*5*5:324*5*5-1]), .o_out_fmap(xor_out[323*8*8*bW:324*8*8*bW-1]));
convchan2 c_2_324 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[324*5*5:325*5*5-1]), .o_out_fmap(xor_out[324*8*8*bW:325*8*8*bW-1]));
convchan2 c_2_325 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[325*5*5:326*5*5-1]), .o_out_fmap(xor_out[325*8*8*bW:326*8*8*bW-1]));
convchan2 c_2_326 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[326*5*5:327*5*5-1]), .o_out_fmap(xor_out[326*8*8*bW:327*8*8*bW-1]));
convchan2 c_2_327 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[327*5*5:328*5*5-1]), .o_out_fmap(xor_out[327*8*8*bW:328*8*8*bW-1]));
convchan2 c_2_328 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[328*5*5:329*5*5-1]), .o_out_fmap(xor_out[328*8*8*bW:329*8*8*bW-1]));
convchan2 c_2_329 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[329*5*5:330*5*5-1]), .o_out_fmap(xor_out[329*8*8*bW:330*8*8*bW-1]));
convchan2 c_2_330 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[330*5*5:331*5*5-1]), .o_out_fmap(xor_out[330*8*8*bW:331*8*8*bW-1]));
convchan2 c_2_331 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[331*5*5:332*5*5-1]), .o_out_fmap(xor_out[331*8*8*bW:332*8*8*bW-1]));
convchan2 c_2_332 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[332*5*5:333*5*5-1]), .o_out_fmap(xor_out[332*8*8*bW:333*8*8*bW-1]));
convchan2 c_2_333 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[333*5*5:334*5*5-1]), .o_out_fmap(xor_out[333*8*8*bW:334*8*8*bW-1]));
convchan2 c_2_334 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[334*5*5:335*5*5-1]), .o_out_fmap(xor_out[334*8*8*bW:335*8*8*bW-1]));
convchan2 c_2_335 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[335*5*5:336*5*5-1]), .o_out_fmap(xor_out[335*8*8*bW:336*8*8*bW-1]));
convchan2 c_2_336 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[336*5*5:337*5*5-1]), .o_out_fmap(xor_out[336*8*8*bW:337*8*8*bW-1]));
convchan2 c_2_337 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[337*5*5:338*5*5-1]), .o_out_fmap(xor_out[337*8*8*bW:338*8*8*bW-1]));
convchan2 c_2_338 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[338*5*5:339*5*5-1]), .o_out_fmap(xor_out[338*8*8*bW:339*8*8*bW-1]));
convchan2 c_2_339 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[339*5*5:340*5*5-1]), .o_out_fmap(xor_out[339*8*8*bW:340*8*8*bW-1]));
convchan2 c_2_340 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[340*5*5:341*5*5-1]), .o_out_fmap(xor_out[340*8*8*bW:341*8*8*bW-1]));
convchan2 c_2_341 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[341*5*5:342*5*5-1]), .o_out_fmap(xor_out[341*8*8*bW:342*8*8*bW-1]));
convchan2 c_2_342 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[342*5*5:343*5*5-1]), .o_out_fmap(xor_out[342*8*8*bW:343*8*8*bW-1]));
convchan2 c_2_343 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[343*5*5:344*5*5-1]), .o_out_fmap(xor_out[343*8*8*bW:344*8*8*bW-1]));
convchan2 c_2_344 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[344*5*5:345*5*5-1]), .o_out_fmap(xor_out[344*8*8*bW:345*8*8*bW-1]));
convchan2 c_2_345 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[345*5*5:346*5*5-1]), .o_out_fmap(xor_out[345*8*8*bW:346*8*8*bW-1]));
convchan2 c_2_346 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[346*5*5:347*5*5-1]), .o_out_fmap(xor_out[346*8*8*bW:347*8*8*bW-1]));
convchan2 c_2_347 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[347*5*5:348*5*5-1]), .o_out_fmap(xor_out[347*8*8*bW:348*8*8*bW-1]));
convchan2 c_2_348 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[348*5*5:349*5*5-1]), .o_out_fmap(xor_out[348*8*8*bW:349*8*8*bW-1]));
convchan2 c_2_349 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[349*5*5:350*5*5-1]), .o_out_fmap(xor_out[349*8*8*bW:350*8*8*bW-1]));
convchan2 c_2_350 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[350*5*5:351*5*5-1]), .o_out_fmap(xor_out[350*8*8*bW:351*8*8*bW-1]));
convchan2 c_2_351 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[351*5*5:352*5*5-1]), .o_out_fmap(xor_out[351*8*8*bW:352*8*8*bW-1]));
convchan2 c_2_352 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[352*5*5:353*5*5-1]), .o_out_fmap(xor_out[352*8*8*bW:353*8*8*bW-1]));
convchan2 c_2_353 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[353*5*5:354*5*5-1]), .o_out_fmap(xor_out[353*8*8*bW:354*8*8*bW-1]));
convchan2 c_2_354 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[354*5*5:355*5*5-1]), .o_out_fmap(xor_out[354*8*8*bW:355*8*8*bW-1]));
convchan2 c_2_355 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[355*5*5:356*5*5-1]), .o_out_fmap(xor_out[355*8*8*bW:356*8*8*bW-1]));
convchan2 c_2_356 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[356*5*5:357*5*5-1]), .o_out_fmap(xor_out[356*8*8*bW:357*8*8*bW-1]));
convchan2 c_2_357 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[357*5*5:358*5*5-1]), .o_out_fmap(xor_out[357*8*8*bW:358*8*8*bW-1]));
convchan2 c_2_358 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[358*5*5:359*5*5-1]), .o_out_fmap(xor_out[358*8*8*bW:359*8*8*bW-1]));
convchan2 c_2_359 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[359*5*5:360*5*5-1]), .o_out_fmap(xor_out[359*8*8*bW:360*8*8*bW-1]));
convchan2 c_2_360 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[360*5*5:361*5*5-1]), .o_out_fmap(xor_out[360*8*8*bW:361*8*8*bW-1]));
convchan2 c_2_361 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[361*5*5:362*5*5-1]), .o_out_fmap(xor_out[361*8*8*bW:362*8*8*bW-1]));
convchan2 c_2_362 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[362*5*5:363*5*5-1]), .o_out_fmap(xor_out[362*8*8*bW:363*8*8*bW-1]));
convchan2 c_2_363 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[363*5*5:364*5*5-1]), .o_out_fmap(xor_out[363*8*8*bW:364*8*8*bW-1]));
convchan2 c_2_364 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[364*5*5:365*5*5-1]), .o_out_fmap(xor_out[364*8*8*bW:365*8*8*bW-1]));
convchan2 c_2_365 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[365*5*5:366*5*5-1]), .o_out_fmap(xor_out[365*8*8*bW:366*8*8*bW-1]));
convchan2 c_2_366 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[366*5*5:367*5*5-1]), .o_out_fmap(xor_out[366*8*8*bW:367*8*8*bW-1]));
convchan2 c_2_367 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[367*5*5:368*5*5-1]), .o_out_fmap(xor_out[367*8*8*bW:368*8*8*bW-1]));
convchan2 c_2_368 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[368*5*5:369*5*5-1]), .o_out_fmap(xor_out[368*8*8*bW:369*8*8*bW-1]));
convchan2 c_2_369 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[369*5*5:370*5*5-1]), .o_out_fmap(xor_out[369*8*8*bW:370*8*8*bW-1]));
convchan2 c_2_370 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[370*5*5:371*5*5-1]), .o_out_fmap(xor_out[370*8*8*bW:371*8*8*bW-1]));
convchan2 c_2_371 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[371*5*5:372*5*5-1]), .o_out_fmap(xor_out[371*8*8*bW:372*8*8*bW-1]));
convchan2 c_2_372 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[372*5*5:373*5*5-1]), .o_out_fmap(xor_out[372*8*8*bW:373*8*8*bW-1]));
convchan2 c_2_373 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[373*5*5:374*5*5-1]), .o_out_fmap(xor_out[373*8*8*bW:374*8*8*bW-1]));
convchan2 c_2_374 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[374*5*5:375*5*5-1]), .o_out_fmap(xor_out[374*8*8*bW:375*8*8*bW-1]));
convchan2 c_2_375 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[375*5*5:376*5*5-1]), .o_out_fmap(xor_out[375*8*8*bW:376*8*8*bW-1]));
convchan2 c_2_376 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[376*5*5:377*5*5-1]), .o_out_fmap(xor_out[376*8*8*bW:377*8*8*bW-1]));
convchan2 c_2_377 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[377*5*5:378*5*5-1]), .o_out_fmap(xor_out[377*8*8*bW:378*8*8*bW-1]));
convchan2 c_2_378 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[378*5*5:379*5*5-1]), .o_out_fmap(xor_out[378*8*8*bW:379*8*8*bW-1]));
convchan2 c_2_379 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[379*5*5:380*5*5-1]), .o_out_fmap(xor_out[379*8*8*bW:380*8*8*bW-1]));
convchan2 c_2_380 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[380*5*5:381*5*5-1]), .o_out_fmap(xor_out[380*8*8*bW:381*8*8*bW-1]));
convchan2 c_2_381 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[381*5*5:382*5*5-1]), .o_out_fmap(xor_out[381*8*8*bW:382*8*8*bW-1]));
convchan2 c_2_382 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[382*5*5:383*5*5-1]), .o_out_fmap(xor_out[382*8*8*bW:383*8*8*bW-1]));
convchan2 c_2_383 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[383*5*5:384*5*5-1]), .o_out_fmap(xor_out[383*8*8*bW:384*8*8*bW-1]));
convchan2 c_2_384 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[384*5*5:385*5*5-1]), .o_out_fmap(xor_out[384*8*8*bW:385*8*8*bW-1]));
convchan2 c_2_385 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[385*5*5:386*5*5-1]), .o_out_fmap(xor_out[385*8*8*bW:386*8*8*bW-1]));
convchan2 c_2_386 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[386*5*5:387*5*5-1]), .o_out_fmap(xor_out[386*8*8*bW:387*8*8*bW-1]));
convchan2 c_2_387 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[387*5*5:388*5*5-1]), .o_out_fmap(xor_out[387*8*8*bW:388*8*8*bW-1]));
convchan2 c_2_388 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[388*5*5:389*5*5-1]), .o_out_fmap(xor_out[388*8*8*bW:389*8*8*bW-1]));
convchan2 c_2_389 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[389*5*5:390*5*5-1]), .o_out_fmap(xor_out[389*8*8*bW:390*8*8*bW-1]));
convchan2 c_2_390 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[390*5*5:391*5*5-1]), .o_out_fmap(xor_out[390*8*8*bW:391*8*8*bW-1]));
convchan2 c_2_391 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[391*5*5:392*5*5-1]), .o_out_fmap(xor_out[391*8*8*bW:392*8*8*bW-1]));
convchan2 c_2_392 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[392*5*5:393*5*5-1]), .o_out_fmap(xor_out[392*8*8*bW:393*8*8*bW-1]));
convchan2 c_2_393 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[393*5*5:394*5*5-1]), .o_out_fmap(xor_out[393*8*8*bW:394*8*8*bW-1]));
convchan2 c_2_394 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[394*5*5:395*5*5-1]), .o_out_fmap(xor_out[394*8*8*bW:395*8*8*bW-1]));
convchan2 c_2_395 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[395*5*5:396*5*5-1]), .o_out_fmap(xor_out[395*8*8*bW:396*8*8*bW-1]));
convchan2 c_2_396 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[396*5*5:397*5*5-1]), .o_out_fmap(xor_out[396*8*8*bW:397*8*8*bW-1]));
convchan2 c_2_397 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[397*5*5:398*5*5-1]), .o_out_fmap(xor_out[397*8*8*bW:398*8*8*bW-1]));
convchan2 c_2_398 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[398*5*5:399*5*5-1]), .o_out_fmap(xor_out[398*8*8*bW:399*8*8*bW-1]));
convchan2 c_2_399 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[399*5*5:400*5*5-1]), .o_out_fmap(xor_out[399*8*8*bW:400*8*8*bW-1]));
convchan2 c_2_400 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[400*5*5:401*5*5-1]), .o_out_fmap(xor_out[400*8*8*bW:401*8*8*bW-1]));
convchan2 c_2_401 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[401*5*5:402*5*5-1]), .o_out_fmap(xor_out[401*8*8*bW:402*8*8*bW-1]));
convchan2 c_2_402 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[402*5*5:403*5*5-1]), .o_out_fmap(xor_out[402*8*8*bW:403*8*8*bW-1]));
convchan2 c_2_403 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[403*5*5:404*5*5-1]), .o_out_fmap(xor_out[403*8*8*bW:404*8*8*bW-1]));
convchan2 c_2_404 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[404*5*5:405*5*5-1]), .o_out_fmap(xor_out[404*8*8*bW:405*8*8*bW-1]));
convchan2 c_2_405 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[405*5*5:406*5*5-1]), .o_out_fmap(xor_out[405*8*8*bW:406*8*8*bW-1]));
convchan2 c_2_406 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[406*5*5:407*5*5-1]), .o_out_fmap(xor_out[406*8*8*bW:407*8*8*bW-1]));
convchan2 c_2_407 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[407*5*5:408*5*5-1]), .o_out_fmap(xor_out[407*8*8*bW:408*8*8*bW-1]));
convchan2 c_2_408 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[408*5*5:409*5*5-1]), .o_out_fmap(xor_out[408*8*8*bW:409*8*8*bW-1]));
convchan2 c_2_409 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[409*5*5:410*5*5-1]), .o_out_fmap(xor_out[409*8*8*bW:410*8*8*bW-1]));
convchan2 c_2_410 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[410*5*5:411*5*5-1]), .o_out_fmap(xor_out[410*8*8*bW:411*8*8*bW-1]));
convchan2 c_2_411 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[411*5*5:412*5*5-1]), .o_out_fmap(xor_out[411*8*8*bW:412*8*8*bW-1]));
convchan2 c_2_412 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[412*5*5:413*5*5-1]), .o_out_fmap(xor_out[412*8*8*bW:413*8*8*bW-1]));
convchan2 c_2_413 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[413*5*5:414*5*5-1]), .o_out_fmap(xor_out[413*8*8*bW:414*8*8*bW-1]));
convchan2 c_2_414 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[414*5*5:415*5*5-1]), .o_out_fmap(xor_out[414*8*8*bW:415*8*8*bW-1]));
convchan2 c_2_415 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[415*5*5:416*5*5-1]), .o_out_fmap(xor_out[415*8*8*bW:416*8*8*bW-1]));
convchan2 c_2_416 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[416*5*5:417*5*5-1]), .o_out_fmap(xor_out[416*8*8*bW:417*8*8*bW-1]));
convchan2 c_2_417 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[417*5*5:418*5*5-1]), .o_out_fmap(xor_out[417*8*8*bW:418*8*8*bW-1]));
convchan2 c_2_418 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[418*5*5:419*5*5-1]), .o_out_fmap(xor_out[418*8*8*bW:419*8*8*bW-1]));
convchan2 c_2_419 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[419*5*5:420*5*5-1]), .o_out_fmap(xor_out[419*8*8*bW:420*8*8*bW-1]));
convchan2 c_2_420 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[420*5*5:421*5*5-1]), .o_out_fmap(xor_out[420*8*8*bW:421*8*8*bW-1]));
convchan2 c_2_421 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[421*5*5:422*5*5-1]), .o_out_fmap(xor_out[421*8*8*bW:422*8*8*bW-1]));
convchan2 c_2_422 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[422*5*5:423*5*5-1]), .o_out_fmap(xor_out[422*8*8*bW:423*8*8*bW-1]));
convchan2 c_2_423 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[423*5*5:424*5*5-1]), .o_out_fmap(xor_out[423*8*8*bW:424*8*8*bW-1]));
convchan2 c_2_424 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[424*5*5:425*5*5-1]), .o_out_fmap(xor_out[424*8*8*bW:425*8*8*bW-1]));
convchan2 c_2_425 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[425*5*5:426*5*5-1]), .o_out_fmap(xor_out[425*8*8*bW:426*8*8*bW-1]));
convchan2 c_2_426 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[426*5*5:427*5*5-1]), .o_out_fmap(xor_out[426*8*8*bW:427*8*8*bW-1]));
convchan2 c_2_427 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[427*5*5:428*5*5-1]), .o_out_fmap(xor_out[427*8*8*bW:428*8*8*bW-1]));
convchan2 c_2_428 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[428*5*5:429*5*5-1]), .o_out_fmap(xor_out[428*8*8*bW:429*8*8*bW-1]));
convchan2 c_2_429 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[429*5*5:430*5*5-1]), .o_out_fmap(xor_out[429*8*8*bW:430*8*8*bW-1]));
convchan2 c_2_430 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[430*5*5:431*5*5-1]), .o_out_fmap(xor_out[430*8*8*bW:431*8*8*bW-1]));
convchan2 c_2_431 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[431*5*5:432*5*5-1]), .o_out_fmap(xor_out[431*8*8*bW:432*8*8*bW-1]));
convchan2 c_2_432 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[432*5*5:433*5*5-1]), .o_out_fmap(xor_out[432*8*8*bW:433*8*8*bW-1]));
convchan2 c_2_433 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[433*5*5:434*5*5-1]), .o_out_fmap(xor_out[433*8*8*bW:434*8*8*bW-1]));
convchan2 c_2_434 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[434*5*5:435*5*5-1]), .o_out_fmap(xor_out[434*8*8*bW:435*8*8*bW-1]));
convchan2 c_2_435 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[435*5*5:436*5*5-1]), .o_out_fmap(xor_out[435*8*8*bW:436*8*8*bW-1]));
convchan2 c_2_436 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[436*5*5:437*5*5-1]), .o_out_fmap(xor_out[436*8*8*bW:437*8*8*bW-1]));
convchan2 c_2_437 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[437*5*5:438*5*5-1]), .o_out_fmap(xor_out[437*8*8*bW:438*8*8*bW-1]));
convchan2 c_2_438 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[438*5*5:439*5*5-1]), .o_out_fmap(xor_out[438*8*8*bW:439*8*8*bW-1]));
convchan2 c_2_439 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[439*5*5:440*5*5-1]), .o_out_fmap(xor_out[439*8*8*bW:440*8*8*bW-1]));
convchan2 c_2_440 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[440*5*5:441*5*5-1]), .o_out_fmap(xor_out[440*8*8*bW:441*8*8*bW-1]));
convchan2 c_2_441 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[441*5*5:442*5*5-1]), .o_out_fmap(xor_out[441*8*8*bW:442*8*8*bW-1]));
convchan2 c_2_442 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[442*5*5:443*5*5-1]), .o_out_fmap(xor_out[442*8*8*bW:443*8*8*bW-1]));
convchan2 c_2_443 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[443*5*5:444*5*5-1]), .o_out_fmap(xor_out[443*8*8*bW:444*8*8*bW-1]));
convchan2 c_2_444 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[444*5*5:445*5*5-1]), .o_out_fmap(xor_out[444*8*8*bW:445*8*8*bW-1]));
convchan2 c_2_445 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[445*5*5:446*5*5-1]), .o_out_fmap(xor_out[445*8*8*bW:446*8*8*bW-1]));
convchan2 c_2_446 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[446*5*5:447*5*5-1]), .o_out_fmap(xor_out[446*8*8*bW:447*8*8*bW-1]));
convchan2 c_2_447 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[447*5*5:448*5*5-1]), .o_out_fmap(xor_out[447*8*8*bW:448*8*8*bW-1]));
convchan2 c_2_448 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[448*5*5:449*5*5-1]), .o_out_fmap(xor_out[448*8*8*bW:449*8*8*bW-1]));
convchan2 c_2_449 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[449*5*5:450*5*5-1]), .o_out_fmap(xor_out[449*8*8*bW:450*8*8*bW-1]));
convchan2 c_2_450 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[450*5*5:451*5*5-1]), .o_out_fmap(xor_out[450*8*8*bW:451*8*8*bW-1]));
convchan2 c_2_451 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[451*5*5:452*5*5-1]), .o_out_fmap(xor_out[451*8*8*bW:452*8*8*bW-1]));
convchan2 c_2_452 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[452*5*5:453*5*5-1]), .o_out_fmap(xor_out[452*8*8*bW:453*8*8*bW-1]));
convchan2 c_2_453 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[453*5*5:454*5*5-1]), .o_out_fmap(xor_out[453*8*8*bW:454*8*8*bW-1]));
convchan2 c_2_454 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[454*5*5:455*5*5-1]), .o_out_fmap(xor_out[454*8*8*bW:455*8*8*bW-1]));
convchan2 c_2_455 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[455*5*5:456*5*5-1]), .o_out_fmap(xor_out[455*8*8*bW:456*8*8*bW-1]));
convchan2 c_2_456 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[456*5*5:457*5*5-1]), .o_out_fmap(xor_out[456*8*8*bW:457*8*8*bW-1]));
convchan2 c_2_457 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[457*5*5:458*5*5-1]), .o_out_fmap(xor_out[457*8*8*bW:458*8*8*bW-1]));
convchan2 c_2_458 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[458*5*5:459*5*5-1]), .o_out_fmap(xor_out[458*8*8*bW:459*8*8*bW-1]));
convchan2 c_2_459 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[459*5*5:460*5*5-1]), .o_out_fmap(xor_out[459*8*8*bW:460*8*8*bW-1]));
convchan2 c_2_460 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[460*5*5:461*5*5-1]), .o_out_fmap(xor_out[460*8*8*bW:461*8*8*bW-1]));
convchan2 c_2_461 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[461*5*5:462*5*5-1]), .o_out_fmap(xor_out[461*8*8*bW:462*8*8*bW-1]));
convchan2 c_2_462 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[462*5*5:463*5*5-1]), .o_out_fmap(xor_out[462*8*8*bW:463*8*8*bW-1]));
convchan2 c_2_463 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[463*5*5:464*5*5-1]), .o_out_fmap(xor_out[463*8*8*bW:464*8*8*bW-1]));
convchan2 c_2_464 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[464*5*5:465*5*5-1]), .o_out_fmap(xor_out[464*8*8*bW:465*8*8*bW-1]));
convchan2 c_2_465 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[465*5*5:466*5*5-1]), .o_out_fmap(xor_out[465*8*8*bW:466*8*8*bW-1]));
convchan2 c_2_466 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[466*5*5:467*5*5-1]), .o_out_fmap(xor_out[466*8*8*bW:467*8*8*bW-1]));
convchan2 c_2_467 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[467*5*5:468*5*5-1]), .o_out_fmap(xor_out[467*8*8*bW:468*8*8*bW-1]));
convchan2 c_2_468 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[468*5*5:469*5*5-1]), .o_out_fmap(xor_out[468*8*8*bW:469*8*8*bW-1]));
convchan2 c_2_469 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[469*5*5:470*5*5-1]), .o_out_fmap(xor_out[469*8*8*bW:470*8*8*bW-1]));
convchan2 c_2_470 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[470*5*5:471*5*5-1]), .o_out_fmap(xor_out[470*8*8*bW:471*8*8*bW-1]));
convchan2 c_2_471 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[471*5*5:472*5*5-1]), .o_out_fmap(xor_out[471*8*8*bW:472*8*8*bW-1]));
convchan2 c_2_472 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[472*5*5:473*5*5-1]), .o_out_fmap(xor_out[472*8*8*bW:473*8*8*bW-1]));
convchan2 c_2_473 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[473*5*5:474*5*5-1]), .o_out_fmap(xor_out[473*8*8*bW:474*8*8*bW-1]));
convchan2 c_2_474 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[474*5*5:475*5*5-1]), .o_out_fmap(xor_out[474*8*8*bW:475*8*8*bW-1]));
convchan2 c_2_475 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[475*5*5:476*5*5-1]), .o_out_fmap(xor_out[475*8*8*bW:476*8*8*bW-1]));
convchan2 c_2_476 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[476*5*5:477*5*5-1]), .o_out_fmap(xor_out[476*8*8*bW:477*8*8*bW-1]));
convchan2 c_2_477 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[477*5*5:478*5*5-1]), .o_out_fmap(xor_out[477*8*8*bW:478*8*8*bW-1]));
convchan2 c_2_478 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[478*5*5:479*5*5-1]), .o_out_fmap(xor_out[478*8*8*bW:479*8*8*bW-1]));
convchan2 c_2_479 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[479*5*5:480*5*5-1]), .o_out_fmap(xor_out[479*8*8*bW:480*8*8*bW-1]));
convchan2 c_2_480 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[480*5*5:481*5*5-1]), .o_out_fmap(xor_out[480*8*8*bW:481*8*8*bW-1]));
convchan2 c_2_481 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[481*5*5:482*5*5-1]), .o_out_fmap(xor_out[481*8*8*bW:482*8*8*bW-1]));
convchan2 c_2_482 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[482*5*5:483*5*5-1]), .o_out_fmap(xor_out[482*8*8*bW:483*8*8*bW-1]));
convchan2 c_2_483 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[483*5*5:484*5*5-1]), .o_out_fmap(xor_out[483*8*8*bW:484*8*8*bW-1]));
convchan2 c_2_484 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[484*5*5:485*5*5-1]), .o_out_fmap(xor_out[484*8*8*bW:485*8*8*bW-1]));
convchan2 c_2_485 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[485*5*5:486*5*5-1]), .o_out_fmap(xor_out[485*8*8*bW:486*8*8*bW-1]));
convchan2 c_2_486 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[486*5*5:487*5*5-1]), .o_out_fmap(xor_out[486*8*8*bW:487*8*8*bW-1]));
convchan2 c_2_487 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[487*5*5:488*5*5-1]), .o_out_fmap(xor_out[487*8*8*bW:488*8*8*bW-1]));
convchan2 c_2_488 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[488*5*5:489*5*5-1]), .o_out_fmap(xor_out[488*8*8*bW:489*8*8*bW-1]));
convchan2 c_2_489 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[489*5*5:490*5*5-1]), .o_out_fmap(xor_out[489*8*8*bW:490*8*8*bW-1]));
convchan2 c_2_490 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[490*5*5:491*5*5-1]), .o_out_fmap(xor_out[490*8*8*bW:491*8*8*bW-1]));
convchan2 c_2_491 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[491*5*5:492*5*5-1]), .o_out_fmap(xor_out[491*8*8*bW:492*8*8*bW-1]));
convchan2 c_2_492 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[492*5*5:493*5*5-1]), .o_out_fmap(xor_out[492*8*8*bW:493*8*8*bW-1]));
convchan2 c_2_493 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[493*5*5:494*5*5-1]), .o_out_fmap(xor_out[493*8*8*bW:494*8*8*bW-1]));
convchan2 c_2_494 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[494*5*5:495*5*5-1]), .o_out_fmap(xor_out[494*8*8*bW:495*8*8*bW-1]));
convchan2 c_2_495 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[495*5*5:496*5*5-1]), .o_out_fmap(xor_out[495*8*8*bW:496*8*8*bW-1]));
convchan2 c_2_496 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[496*5*5:497*5*5-1]), .o_out_fmap(xor_out[496*8*8*bW:497*8*8*bW-1]));
convchan2 c_2_497 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[497*5*5:498*5*5-1]), .o_out_fmap(xor_out[497*8*8*bW:498*8*8*bW-1]));
convchan2 c_2_498 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[498*5*5:499*5*5-1]), .o_out_fmap(xor_out[498*8*8*bW:499*8*8*bW-1]));
convchan2 c_2_499 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[499*5*5:500*5*5-1]), .o_out_fmap(xor_out[499*8*8*bW:500*8*8*bW-1]));
convchan2 c_2_500 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[500*5*5:501*5*5-1]), .o_out_fmap(xor_out[500*8*8*bW:501*8*8*bW-1]));
convchan2 c_2_501 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[501*5*5:502*5*5-1]), .o_out_fmap(xor_out[501*8*8*bW:502*8*8*bW-1]));
convchan2 c_2_502 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[502*5*5:503*5*5-1]), .o_out_fmap(xor_out[502*8*8*bW:503*8*8*bW-1]));
convchan2 c_2_503 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[503*5*5:504*5*5-1]), .o_out_fmap(xor_out[503*8*8*bW:504*8*8*bW-1]));
convchan2 c_2_504 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[504*5*5:505*5*5-1]), .o_out_fmap(xor_out[504*8*8*bW:505*8*8*bW-1]));
convchan2 c_2_505 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[505*5*5:506*5*5-1]), .o_out_fmap(xor_out[505*8*8*bW:506*8*8*bW-1]));
convchan2 c_2_506 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[506*5*5:507*5*5-1]), .o_out_fmap(xor_out[506*8*8*bW:507*8*8*bW-1]));
convchan2 c_2_507 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[507*5*5:508*5*5-1]), .o_out_fmap(xor_out[507*8*8*bW:508*8*8*bW-1]));
convchan2 c_2_508 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[508*5*5:509*5*5-1]), .o_out_fmap(xor_out[508*8*8*bW:509*8*8*bW-1]));
convchan2 c_2_509 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[509*5*5:510*5*5-1]), .o_out_fmap(xor_out[509*8*8*bW:510*8*8*bW-1]));
convchan2 c_2_510 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[510*5*5:511*5*5-1]), .o_out_fmap(xor_out[510*8*8*bW:511*8*8*bW-1]));
convchan2 c_2_511 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[511*5*5:512*5*5-1]), .o_out_fmap(xor_out[511*8*8*bW:512*8*8*bW-1]));
convchan2 c_2_512 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[512*5*5:513*5*5-1]), .o_out_fmap(xor_out[512*8*8*bW:513*8*8*bW-1]));
convchan2 c_2_513 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[513*5*5:514*5*5-1]), .o_out_fmap(xor_out[513*8*8*bW:514*8*8*bW-1]));
convchan2 c_2_514 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[514*5*5:515*5*5-1]), .o_out_fmap(xor_out[514*8*8*bW:515*8*8*bW-1]));
convchan2 c_2_515 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[515*5*5:516*5*5-1]), .o_out_fmap(xor_out[515*8*8*bW:516*8*8*bW-1]));
convchan2 c_2_516 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[516*5*5:517*5*5-1]), .o_out_fmap(xor_out[516*8*8*bW:517*8*8*bW-1]));
convchan2 c_2_517 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[517*5*5:518*5*5-1]), .o_out_fmap(xor_out[517*8*8*bW:518*8*8*bW-1]));
convchan2 c_2_518 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[518*5*5:519*5*5-1]), .o_out_fmap(xor_out[518*8*8*bW:519*8*8*bW-1]));
convchan2 c_2_519 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[519*5*5:520*5*5-1]), .o_out_fmap(xor_out[519*8*8*bW:520*8*8*bW-1]));
convchan2 c_2_520 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[520*5*5:521*5*5-1]), .o_out_fmap(xor_out[520*8*8*bW:521*8*8*bW-1]));
convchan2 c_2_521 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[521*5*5:522*5*5-1]), .o_out_fmap(xor_out[521*8*8*bW:522*8*8*bW-1]));
convchan2 c_2_522 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[522*5*5:523*5*5-1]), .o_out_fmap(xor_out[522*8*8*bW:523*8*8*bW-1]));
convchan2 c_2_523 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[523*5*5:524*5*5-1]), .o_out_fmap(xor_out[523*8*8*bW:524*8*8*bW-1]));
convchan2 c_2_524 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[524*5*5:525*5*5-1]), .o_out_fmap(xor_out[524*8*8*bW:525*8*8*bW-1]));
convchan2 c_2_525 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[525*5*5:526*5*5-1]), .o_out_fmap(xor_out[525*8*8*bW:526*8*8*bW-1]));
convchan2 c_2_526 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[526*5*5:527*5*5-1]), .o_out_fmap(xor_out[526*8*8*bW:527*8*8*bW-1]));
convchan2 c_2_527 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[527*5*5:528*5*5-1]), .o_out_fmap(xor_out[527*8*8*bW:528*8*8*bW-1]));
convchan2 c_2_528 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[528*5*5:529*5*5-1]), .o_out_fmap(xor_out[528*8*8*bW:529*8*8*bW-1]));
convchan2 c_2_529 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[529*5*5:530*5*5-1]), .o_out_fmap(xor_out[529*8*8*bW:530*8*8*bW-1]));
convchan2 c_2_530 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[530*5*5:531*5*5-1]), .o_out_fmap(xor_out[530*8*8*bW:531*8*8*bW-1]));
convchan2 c_2_531 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[531*5*5:532*5*5-1]), .o_out_fmap(xor_out[531*8*8*bW:532*8*8*bW-1]));
convchan2 c_2_532 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[532*5*5:533*5*5-1]), .o_out_fmap(xor_out[532*8*8*bW:533*8*8*bW-1]));
convchan2 c_2_533 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[533*5*5:534*5*5-1]), .o_out_fmap(xor_out[533*8*8*bW:534*8*8*bW-1]));
convchan2 c_2_534 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[534*5*5:535*5*5-1]), .o_out_fmap(xor_out[534*8*8*bW:535*8*8*bW-1]));
convchan2 c_2_535 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[535*5*5:536*5*5-1]), .o_out_fmap(xor_out[535*8*8*bW:536*8*8*bW-1]));
convchan2 c_2_536 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[536*5*5:537*5*5-1]), .o_out_fmap(xor_out[536*8*8*bW:537*8*8*bW-1]));
convchan2 c_2_537 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[537*5*5:538*5*5-1]), .o_out_fmap(xor_out[537*8*8*bW:538*8*8*bW-1]));
convchan2 c_2_538 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[538*5*5:539*5*5-1]), .o_out_fmap(xor_out[538*8*8*bW:539*8*8*bW-1]));
convchan2 c_2_539 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[539*5*5:540*5*5-1]), .o_out_fmap(xor_out[539*8*8*bW:540*8*8*bW-1]));
convchan2 c_2_540 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[540*5*5:541*5*5-1]), .o_out_fmap(xor_out[540*8*8*bW:541*8*8*bW-1]));
convchan2 c_2_541 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[541*5*5:542*5*5-1]), .o_out_fmap(xor_out[541*8*8*bW:542*8*8*bW-1]));
convchan2 c_2_542 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[542*5*5:543*5*5-1]), .o_out_fmap(xor_out[542*8*8*bW:543*8*8*bW-1]));
convchan2 c_2_543 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[543*5*5:544*5*5-1]), .o_out_fmap(xor_out[543*8*8*bW:544*8*8*bW-1]));
convchan2 c_2_544 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[544*5*5:545*5*5-1]), .o_out_fmap(xor_out[544*8*8*bW:545*8*8*bW-1]));
convchan2 c_2_545 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[545*5*5:546*5*5-1]), .o_out_fmap(xor_out[545*8*8*bW:546*8*8*bW-1]));
convchan2 c_2_546 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[546*5*5:547*5*5-1]), .o_out_fmap(xor_out[546*8*8*bW:547*8*8*bW-1]));
convchan2 c_2_547 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[547*5*5:548*5*5-1]), .o_out_fmap(xor_out[547*8*8*bW:548*8*8*bW-1]));
convchan2 c_2_548 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[548*5*5:549*5*5-1]), .o_out_fmap(xor_out[548*8*8*bW:549*8*8*bW-1]));
convchan2 c_2_549 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[549*5*5:550*5*5-1]), .o_out_fmap(xor_out[549*8*8*bW:550*8*8*bW-1]));
convchan2 c_2_550 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[550*5*5:551*5*5-1]), .o_out_fmap(xor_out[550*8*8*bW:551*8*8*bW-1]));
convchan2 c_2_551 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[551*5*5:552*5*5-1]), .o_out_fmap(xor_out[551*8*8*bW:552*8*8*bW-1]));
convchan2 c_2_552 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[552*5*5:553*5*5-1]), .o_out_fmap(xor_out[552*8*8*bW:553*8*8*bW-1]));
convchan2 c_2_553 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[553*5*5:554*5*5-1]), .o_out_fmap(xor_out[553*8*8*bW:554*8*8*bW-1]));
convchan2 c_2_554 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[554*5*5:555*5*5-1]), .o_out_fmap(xor_out[554*8*8*bW:555*8*8*bW-1]));
convchan2 c_2_555 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[555*5*5:556*5*5-1]), .o_out_fmap(xor_out[555*8*8*bW:556*8*8*bW-1]));
convchan2 c_2_556 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[556*5*5:557*5*5-1]), .o_out_fmap(xor_out[556*8*8*bW:557*8*8*bW-1]));
convchan2 c_2_557 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[557*5*5:558*5*5-1]), .o_out_fmap(xor_out[557*8*8*bW:558*8*8*bW-1]));
convchan2 c_2_558 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[558*5*5:559*5*5-1]), .o_out_fmap(xor_out[558*8*8*bW:559*8*8*bW-1]));
convchan2 c_2_559 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[559*5*5:560*5*5-1]), .o_out_fmap(xor_out[559*8*8*bW:560*8*8*bW-1]));
convchan2 c_2_560 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[560*5*5:561*5*5-1]), .o_out_fmap(xor_out[560*8*8*bW:561*8*8*bW-1]));
convchan2 c_2_561 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[561*5*5:562*5*5-1]), .o_out_fmap(xor_out[561*8*8*bW:562*8*8*bW-1]));
convchan2 c_2_562 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[562*5*5:563*5*5-1]), .o_out_fmap(xor_out[562*8*8*bW:563*8*8*bW-1]));
convchan2 c_2_563 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[563*5*5:564*5*5-1]), .o_out_fmap(xor_out[563*8*8*bW:564*8*8*bW-1]));
convchan2 c_2_564 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[564*5*5:565*5*5-1]), .o_out_fmap(xor_out[564*8*8*bW:565*8*8*bW-1]));
convchan2 c_2_565 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[565*5*5:566*5*5-1]), .o_out_fmap(xor_out[565*8*8*bW:566*8*8*bW-1]));
convchan2 c_2_566 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[566*5*5:567*5*5-1]), .o_out_fmap(xor_out[566*8*8*bW:567*8*8*bW-1]));
convchan2 c_2_567 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[567*5*5:568*5*5-1]), .o_out_fmap(xor_out[567*8*8*bW:568*8*8*bW-1]));
convchan2 c_2_568 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[568*5*5:569*5*5-1]), .o_out_fmap(xor_out[568*8*8*bW:569*8*8*bW-1]));
convchan2 c_2_569 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[569*5*5:570*5*5-1]), .o_out_fmap(xor_out[569*8*8*bW:570*8*8*bW-1]));
convchan2 c_2_570 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[570*5*5:571*5*5-1]), .o_out_fmap(xor_out[570*8*8*bW:571*8*8*bW-1]));
convchan2 c_2_571 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[571*5*5:572*5*5-1]), .o_out_fmap(xor_out[571*8*8*bW:572*8*8*bW-1]));
convchan2 c_2_572 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[572*5*5:573*5*5-1]), .o_out_fmap(xor_out[572*8*8*bW:573*8*8*bW-1]));
convchan2 c_2_573 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[573*5*5:574*5*5-1]), .o_out_fmap(xor_out[573*8*8*bW:574*8*8*bW-1]));
convchan2 c_2_574 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[574*5*5:575*5*5-1]), .o_out_fmap(xor_out[574*8*8*bW:575*8*8*bW-1]));
convchan2 c_2_575 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[575*5*5:576*5*5-1]), .o_out_fmap(xor_out[575*8*8*bW:576*8*8*bW-1]));
convchan2 c_2_576 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[576*5*5:577*5*5-1]), .o_out_fmap(xor_out[576*8*8*bW:577*8*8*bW-1]));
convchan2 c_2_577 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[577*5*5:578*5*5-1]), .o_out_fmap(xor_out[577*8*8*bW:578*8*8*bW-1]));
convchan2 c_2_578 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[578*5*5:579*5*5-1]), .o_out_fmap(xor_out[578*8*8*bW:579*8*8*bW-1]));
convchan2 c_2_579 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[579*5*5:580*5*5-1]), .o_out_fmap(xor_out[579*8*8*bW:580*8*8*bW-1]));
convchan2 c_2_580 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[580*5*5:581*5*5-1]), .o_out_fmap(xor_out[580*8*8*bW:581*8*8*bW-1]));
convchan2 c_2_581 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[581*5*5:582*5*5-1]), .o_out_fmap(xor_out[581*8*8*bW:582*8*8*bW-1]));
convchan2 c_2_582 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[582*5*5:583*5*5-1]), .o_out_fmap(xor_out[582*8*8*bW:583*8*8*bW-1]));
convchan2 c_2_583 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[583*5*5:584*5*5-1]), .o_out_fmap(xor_out[583*8*8*bW:584*8*8*bW-1]));
convchan2 c_2_584 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[584*5*5:585*5*5-1]), .o_out_fmap(xor_out[584*8*8*bW:585*8*8*bW-1]));
convchan2 c_2_585 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[585*5*5:586*5*5-1]), .o_out_fmap(xor_out[585*8*8*bW:586*8*8*bW-1]));
convchan2 c_2_586 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[586*5*5:587*5*5-1]), .o_out_fmap(xor_out[586*8*8*bW:587*8*8*bW-1]));
convchan2 c_2_587 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[587*5*5:588*5*5-1]), .o_out_fmap(xor_out[587*8*8*bW:588*8*8*bW-1]));
convchan2 c_2_588 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[588*5*5:589*5*5-1]), .o_out_fmap(xor_out[588*8*8*bW:589*8*8*bW-1]));
convchan2 c_2_589 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[589*5*5:590*5*5-1]), .o_out_fmap(xor_out[589*8*8*bW:590*8*8*bW-1]));
convchan2 c_2_590 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[590*5*5:591*5*5-1]), .o_out_fmap(xor_out[590*8*8*bW:591*8*8*bW-1]));
convchan2 c_2_591 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[591*5*5:592*5*5-1]), .o_out_fmap(xor_out[591*8*8*bW:592*8*8*bW-1]));
convchan2 c_2_592 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[592*5*5:593*5*5-1]), .o_out_fmap(xor_out[592*8*8*bW:593*8*8*bW-1]));
convchan2 c_2_593 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[593*5*5:594*5*5-1]), .o_out_fmap(xor_out[593*8*8*bW:594*8*8*bW-1]));
convchan2 c_2_594 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[594*5*5:595*5*5-1]), .o_out_fmap(xor_out[594*8*8*bW:595*8*8*bW-1]));
convchan2 c_2_595 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[595*5*5:596*5*5-1]), .o_out_fmap(xor_out[595*8*8*bW:596*8*8*bW-1]));
convchan2 c_2_596 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[596*5*5:597*5*5-1]), .o_out_fmap(xor_out[596*8*8*bW:597*8*8*bW-1]));
convchan2 c_2_597 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[597*5*5:598*5*5-1]), .o_out_fmap(xor_out[597*8*8*bW:598*8*8*bW-1]));
convchan2 c_2_598 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[598*5*5:599*5*5-1]), .o_out_fmap(xor_out[598*8*8*bW:599*8*8*bW-1]));
convchan2 c_2_599 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[599*5*5:600*5*5-1]), .o_out_fmap(xor_out[599*8*8*bW:600*8*8*bW-1]));
convchan2 c_2_600 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[600*5*5:601*5*5-1]), .o_out_fmap(xor_out[600*8*8*bW:601*8*8*bW-1]));
convchan2 c_2_601 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[601*5*5:602*5*5-1]), .o_out_fmap(xor_out[601*8*8*bW:602*8*8*bW-1]));
convchan2 c_2_602 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[602*5*5:603*5*5-1]), .o_out_fmap(xor_out[602*8*8*bW:603*8*8*bW-1]));
convchan2 c_2_603 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[603*5*5:604*5*5-1]), .o_out_fmap(xor_out[603*8*8*bW:604*8*8*bW-1]));
convchan2 c_2_604 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[604*5*5:605*5*5-1]), .o_out_fmap(xor_out[604*8*8*bW:605*8*8*bW-1]));
convchan2 c_2_605 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[605*5*5:606*5*5-1]), .o_out_fmap(xor_out[605*8*8*bW:606*8*8*bW-1]));
convchan2 c_2_606 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[606*5*5:607*5*5-1]), .o_out_fmap(xor_out[606*8*8*bW:607*8*8*bW-1]));
convchan2 c_2_607 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[607*5*5:608*5*5-1]), .o_out_fmap(xor_out[607*8*8*bW:608*8*8*bW-1]));
convchan2 c_2_608 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[608*5*5:609*5*5-1]), .o_out_fmap(xor_out[608*8*8*bW:609*8*8*bW-1]));
convchan2 c_2_609 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[609*5*5:610*5*5-1]), .o_out_fmap(xor_out[609*8*8*bW:610*8*8*bW-1]));
convchan2 c_2_610 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[610*5*5:611*5*5-1]), .o_out_fmap(xor_out[610*8*8*bW:611*8*8*bW-1]));
convchan2 c_2_611 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[611*5*5:612*5*5-1]), .o_out_fmap(xor_out[611*8*8*bW:612*8*8*bW-1]));
convchan2 c_2_612 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[612*5*5:613*5*5-1]), .o_out_fmap(xor_out[612*8*8*bW:613*8*8*bW-1]));
convchan2 c_2_613 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[613*5*5:614*5*5-1]), .o_out_fmap(xor_out[613*8*8*bW:614*8*8*bW-1]));
convchan2 c_2_614 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[614*5*5:615*5*5-1]), .o_out_fmap(xor_out[614*8*8*bW:615*8*8*bW-1]));
convchan2 c_2_615 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[615*5*5:616*5*5-1]), .o_out_fmap(xor_out[615*8*8*bW:616*8*8*bW-1]));
convchan2 c_2_616 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[616*5*5:617*5*5-1]), .o_out_fmap(xor_out[616*8*8*bW:617*8*8*bW-1]));
convchan2 c_2_617 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[617*5*5:618*5*5-1]), .o_out_fmap(xor_out[617*8*8*bW:618*8*8*bW-1]));
convchan2 c_2_618 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[618*5*5:619*5*5-1]), .o_out_fmap(xor_out[618*8*8*bW:619*8*8*bW-1]));
convchan2 c_2_619 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[619*5*5:620*5*5-1]), .o_out_fmap(xor_out[619*8*8*bW:620*8*8*bW-1]));
convchan2 c_2_620 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[620*5*5:621*5*5-1]), .o_out_fmap(xor_out[620*8*8*bW:621*8*8*bW-1]));
convchan2 c_2_621 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[621*5*5:622*5*5-1]), .o_out_fmap(xor_out[621*8*8*bW:622*8*8*bW-1]));
convchan2 c_2_622 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[622*5*5:623*5*5-1]), .o_out_fmap(xor_out[622*8*8*bW:623*8*8*bW-1]));
convchan2 c_2_623 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[623*5*5:624*5*5-1]), .o_out_fmap(xor_out[623*8*8*bW:624*8*8*bW-1]));
convchan2 c_2_624 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[624*5*5:625*5*5-1]), .o_out_fmap(xor_out[624*8*8*bW:625*8*8*bW-1]));
convchan2 c_2_625 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[625*5*5:626*5*5-1]), .o_out_fmap(xor_out[625*8*8*bW:626*8*8*bW-1]));
convchan2 c_2_626 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[626*5*5:627*5*5-1]), .o_out_fmap(xor_out[626*8*8*bW:627*8*8*bW-1]));
convchan2 c_2_627 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[627*5*5:628*5*5-1]), .o_out_fmap(xor_out[627*8*8*bW:628*8*8*bW-1]));
convchan2 c_2_628 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[628*5*5:629*5*5-1]), .o_out_fmap(xor_out[628*8*8*bW:629*8*8*bW-1]));
convchan2 c_2_629 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[629*5*5:630*5*5-1]), .o_out_fmap(xor_out[629*8*8*bW:630*8*8*bW-1]));
convchan2 c_2_630 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[630*5*5:631*5*5-1]), .o_out_fmap(xor_out[630*8*8*bW:631*8*8*bW-1]));
convchan2 c_2_631 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[631*5*5:632*5*5-1]), .o_out_fmap(xor_out[631*8*8*bW:632*8*8*bW-1]));
convchan2 c_2_632 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[632*5*5:633*5*5-1]), .o_out_fmap(xor_out[632*8*8*bW:633*8*8*bW-1]));
convchan2 c_2_633 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[633*5*5:634*5*5-1]), .o_out_fmap(xor_out[633*8*8*bW:634*8*8*bW-1]));
convchan2 c_2_634 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[634*5*5:635*5*5-1]), .o_out_fmap(xor_out[634*8*8*bW:635*8*8*bW-1]));
convchan2 c_2_635 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[635*5*5:636*5*5-1]), .o_out_fmap(xor_out[635*8*8*bW:636*8*8*bW-1]));
convchan2 c_2_636 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[636*5*5:637*5*5-1]), .o_out_fmap(xor_out[636*8*8*bW:637*8*8*bW-1]));
convchan2 c_2_637 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[637*5*5:638*5*5-1]), .o_out_fmap(xor_out[637*8*8*bW:638*8*8*bW-1]));
convchan2 c_2_638 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[638*5*5:639*5*5-1]), .o_out_fmap(xor_out[638*8*8*bW:639*8*8*bW-1]));
convchan2 c_2_639 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[639*5*5:640*5*5-1]), .o_out_fmap(xor_out[639*8*8*bW:640*8*8*bW-1]));
convchan2 c_2_640 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[640*5*5:641*5*5-1]), .o_out_fmap(xor_out[640*8*8*bW:641*8*8*bW-1]));
convchan2 c_2_641 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[641*5*5:642*5*5-1]), .o_out_fmap(xor_out[641*8*8*bW:642*8*8*bW-1]));
convchan2 c_2_642 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[642*5*5:643*5*5-1]), .o_out_fmap(xor_out[642*8*8*bW:643*8*8*bW-1]));
convchan2 c_2_643 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[643*5*5:644*5*5-1]), .o_out_fmap(xor_out[643*8*8*bW:644*8*8*bW-1]));
convchan2 c_2_644 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[644*5*5:645*5*5-1]), .o_out_fmap(xor_out[644*8*8*bW:645*8*8*bW-1]));
convchan2 c_2_645 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[645*5*5:646*5*5-1]), .o_out_fmap(xor_out[645*8*8*bW:646*8*8*bW-1]));
convchan2 c_2_646 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[646*5*5:647*5*5-1]), .o_out_fmap(xor_out[646*8*8*bW:647*8*8*bW-1]));
convchan2 c_2_647 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[647*5*5:648*5*5-1]), .o_out_fmap(xor_out[647*8*8*bW:648*8*8*bW-1]));
convchan2 c_2_648 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[648*5*5:649*5*5-1]), .o_out_fmap(xor_out[648*8*8*bW:649*8*8*bW-1]));
convchan2 c_2_649 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[649*5*5:650*5*5-1]), .o_out_fmap(xor_out[649*8*8*bW:650*8*8*bW-1]));
convchan2 c_2_650 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[650*5*5:651*5*5-1]), .o_out_fmap(xor_out[650*8*8*bW:651*8*8*bW-1]));
convchan2 c_2_651 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[651*5*5:652*5*5-1]), .o_out_fmap(xor_out[651*8*8*bW:652*8*8*bW-1]));
convchan2 c_2_652 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[652*5*5:653*5*5-1]), .o_out_fmap(xor_out[652*8*8*bW:653*8*8*bW-1]));
convchan2 c_2_653 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[653*5*5:654*5*5-1]), .o_out_fmap(xor_out[653*8*8*bW:654*8*8*bW-1]));
convchan2 c_2_654 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[654*5*5:655*5*5-1]), .o_out_fmap(xor_out[654*8*8*bW:655*8*8*bW-1]));
convchan2 c_2_655 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[655*5*5:656*5*5-1]), .o_out_fmap(xor_out[655*8*8*bW:656*8*8*bW-1]));
convchan2 c_2_656 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[656*5*5:657*5*5-1]), .o_out_fmap(xor_out[656*8*8*bW:657*8*8*bW-1]));
convchan2 c_2_657 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[657*5*5:658*5*5-1]), .o_out_fmap(xor_out[657*8*8*bW:658*8*8*bW-1]));
convchan2 c_2_658 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[658*5*5:659*5*5-1]), .o_out_fmap(xor_out[658*8*8*bW:659*8*8*bW-1]));
convchan2 c_2_659 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[659*5*5:660*5*5-1]), .o_out_fmap(xor_out[659*8*8*bW:660*8*8*bW-1]));
convchan2 c_2_660 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[660*5*5:661*5*5-1]), .o_out_fmap(xor_out[660*8*8*bW:661*8*8*bW-1]));
convchan2 c_2_661 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[661*5*5:662*5*5-1]), .o_out_fmap(xor_out[661*8*8*bW:662*8*8*bW-1]));
convchan2 c_2_662 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[662*5*5:663*5*5-1]), .o_out_fmap(xor_out[662*8*8*bW:663*8*8*bW-1]));
convchan2 c_2_663 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[663*5*5:664*5*5-1]), .o_out_fmap(xor_out[663*8*8*bW:664*8*8*bW-1]));
convchan2 c_2_664 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[664*5*5:665*5*5-1]), .o_out_fmap(xor_out[664*8*8*bW:665*8*8*bW-1]));
convchan2 c_2_665 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[665*5*5:666*5*5-1]), .o_out_fmap(xor_out[665*8*8*bW:666*8*8*bW-1]));
convchan2 c_2_666 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[666*5*5:667*5*5-1]), .o_out_fmap(xor_out[666*8*8*bW:667*8*8*bW-1]));
convchan2 c_2_667 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[667*5*5:668*5*5-1]), .o_out_fmap(xor_out[667*8*8*bW:668*8*8*bW-1]));
convchan2 c_2_668 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[668*5*5:669*5*5-1]), .o_out_fmap(xor_out[668*8*8*bW:669*8*8*bW-1]));
convchan2 c_2_669 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[669*5*5:670*5*5-1]), .o_out_fmap(xor_out[669*8*8*bW:670*8*8*bW-1]));
convchan2 c_2_670 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[670*5*5:671*5*5-1]), .o_out_fmap(xor_out[670*8*8*bW:671*8*8*bW-1]));
convchan2 c_2_671 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[671*5*5:672*5*5-1]), .o_out_fmap(xor_out[671*8*8*bW:672*8*8*bW-1]));
convchan2 c_2_672 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[672*5*5:673*5*5-1]), .o_out_fmap(xor_out[672*8*8*bW:673*8*8*bW-1]));
convchan2 c_2_673 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[673*5*5:674*5*5-1]), .o_out_fmap(xor_out[673*8*8*bW:674*8*8*bW-1]));
convchan2 c_2_674 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[674*5*5:675*5*5-1]), .o_out_fmap(xor_out[674*8*8*bW:675*8*8*bW-1]));
convchan2 c_2_675 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[675*5*5:676*5*5-1]), .o_out_fmap(xor_out[675*8*8*bW:676*8*8*bW-1]));
convchan2 c_2_676 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[676*5*5:677*5*5-1]), .o_out_fmap(xor_out[676*8*8*bW:677*8*8*bW-1]));
convchan2 c_2_677 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[677*5*5:678*5*5-1]), .o_out_fmap(xor_out[677*8*8*bW:678*8*8*bW-1]));
convchan2 c_2_678 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[678*5*5:679*5*5-1]), .o_out_fmap(xor_out[678*8*8*bW:679*8*8*bW-1]));
convchan2 c_2_679 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[679*5*5:680*5*5-1]), .o_out_fmap(xor_out[679*8*8*bW:680*8*8*bW-1]));
convchan2 c_2_680 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[680*5*5:681*5*5-1]), .o_out_fmap(xor_out[680*8*8*bW:681*8*8*bW-1]));
convchan2 c_2_681 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[681*5*5:682*5*5-1]), .o_out_fmap(xor_out[681*8*8*bW:682*8*8*bW-1]));
convchan2 c_2_682 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[682*5*5:683*5*5-1]), .o_out_fmap(xor_out[682*8*8*bW:683*8*8*bW-1]));
convchan2 c_2_683 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[683*5*5:684*5*5-1]), .o_out_fmap(xor_out[683*8*8*bW:684*8*8*bW-1]));
convchan2 c_2_684 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[684*5*5:685*5*5-1]), .o_out_fmap(xor_out[684*8*8*bW:685*8*8*bW-1]));
convchan2 c_2_685 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[685*5*5:686*5*5-1]), .o_out_fmap(xor_out[685*8*8*bW:686*8*8*bW-1]));
convchan2 c_2_686 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[686*5*5:687*5*5-1]), .o_out_fmap(xor_out[686*8*8*bW:687*8*8*bW-1]));
convchan2 c_2_687 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[687*5*5:688*5*5-1]), .o_out_fmap(xor_out[687*8*8*bW:688*8*8*bW-1]));
convchan2 c_2_688 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[688*5*5:689*5*5-1]), .o_out_fmap(xor_out[688*8*8*bW:689*8*8*bW-1]));
convchan2 c_2_689 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[689*5*5:690*5*5-1]), .o_out_fmap(xor_out[689*8*8*bW:690*8*8*bW-1]));
convchan2 c_2_690 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[690*5*5:691*5*5-1]), .o_out_fmap(xor_out[690*8*8*bW:691*8*8*bW-1]));
convchan2 c_2_691 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[691*5*5:692*5*5-1]), .o_out_fmap(xor_out[691*8*8*bW:692*8*8*bW-1]));
convchan2 c_2_692 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[692*5*5:693*5*5-1]), .o_out_fmap(xor_out[692*8*8*bW:693*8*8*bW-1]));
convchan2 c_2_693 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[693*5*5:694*5*5-1]), .o_out_fmap(xor_out[693*8*8*bW:694*8*8*bW-1]));
convchan2 c_2_694 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[694*5*5:695*5*5-1]), .o_out_fmap(xor_out[694*8*8*bW:695*8*8*bW-1]));
convchan2 c_2_695 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[695*5*5:696*5*5-1]), .o_out_fmap(xor_out[695*8*8*bW:696*8*8*bW-1]));
convchan2 c_2_696 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[696*5*5:697*5*5-1]), .o_out_fmap(xor_out[696*8*8*bW:697*8*8*bW-1]));
convchan2 c_2_697 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[697*5*5:698*5*5-1]), .o_out_fmap(xor_out[697*8*8*bW:698*8*8*bW-1]));
convchan2 c_2_698 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[698*5*5:699*5*5-1]), .o_out_fmap(xor_out[698*8*8*bW:699*8*8*bW-1]));
convchan2 c_2_699 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[699*5*5:700*5*5-1]), .o_out_fmap(xor_out[699*8*8*bW:700*8*8*bW-1]));
convchan2 c_2_700 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[700*5*5:701*5*5-1]), .o_out_fmap(xor_out[700*8*8*bW:701*8*8*bW-1]));
convchan2 c_2_701 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[701*5*5:702*5*5-1]), .o_out_fmap(xor_out[701*8*8*bW:702*8*8*bW-1]));
convchan2 c_2_702 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[702*5*5:703*5*5-1]), .o_out_fmap(xor_out[702*8*8*bW:703*8*8*bW-1]));
convchan2 c_2_703 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[703*5*5:704*5*5-1]), .o_out_fmap(xor_out[703*8*8*bW:704*8*8*bW-1]));
convchan2 c_2_704 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[704*5*5:705*5*5-1]), .o_out_fmap(xor_out[704*8*8*bW:705*8*8*bW-1]));
convchan2 c_2_705 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[705*5*5:706*5*5-1]), .o_out_fmap(xor_out[705*8*8*bW:706*8*8*bW-1]));
convchan2 c_2_706 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[706*5*5:707*5*5-1]), .o_out_fmap(xor_out[706*8*8*bW:707*8*8*bW-1]));
convchan2 c_2_707 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[707*5*5:708*5*5-1]), .o_out_fmap(xor_out[707*8*8*bW:708*8*8*bW-1]));
convchan2 c_2_708 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[708*5*5:709*5*5-1]), .o_out_fmap(xor_out[708*8*8*bW:709*8*8*bW-1]));
convchan2 c_2_709 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[709*5*5:710*5*5-1]), .o_out_fmap(xor_out[709*8*8*bW:710*8*8*bW-1]));
convchan2 c_2_710 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[710*5*5:711*5*5-1]), .o_out_fmap(xor_out[710*8*8*bW:711*8*8*bW-1]));
convchan2 c_2_711 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[711*5*5:712*5*5-1]), .o_out_fmap(xor_out[711*8*8*bW:712*8*8*bW-1]));
convchan2 c_2_712 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[712*5*5:713*5*5-1]), .o_out_fmap(xor_out[712*8*8*bW:713*8*8*bW-1]));
convchan2 c_2_713 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[713*5*5:714*5*5-1]), .o_out_fmap(xor_out[713*8*8*bW:714*8*8*bW-1]));
convchan2 c_2_714 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[714*5*5:715*5*5-1]), .o_out_fmap(xor_out[714*8*8*bW:715*8*8*bW-1]));
convchan2 c_2_715 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[715*5*5:716*5*5-1]), .o_out_fmap(xor_out[715*8*8*bW:716*8*8*bW-1]));
convchan2 c_2_716 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[716*5*5:717*5*5-1]), .o_out_fmap(xor_out[716*8*8*bW:717*8*8*bW-1]));
convchan2 c_2_717 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[717*5*5:718*5*5-1]), .o_out_fmap(xor_out[717*8*8*bW:718*8*8*bW-1]));
convchan2 c_2_718 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[718*5*5:719*5*5-1]), .o_out_fmap(xor_out[718*8*8*bW:719*8*8*bW-1]));
convchan2 c_2_719 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[719*5*5:720*5*5-1]), .o_out_fmap(xor_out[719*8*8*bW:720*8*8*bW-1]));
convchan2 c_2_720 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[720*5*5:721*5*5-1]), .o_out_fmap(xor_out[720*8*8*bW:721*8*8*bW-1]));
convchan2 c_2_721 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[721*5*5:722*5*5-1]), .o_out_fmap(xor_out[721*8*8*bW:722*8*8*bW-1]));
convchan2 c_2_722 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[722*5*5:723*5*5-1]), .o_out_fmap(xor_out[722*8*8*bW:723*8*8*bW-1]));
convchan2 c_2_723 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[723*5*5:724*5*5-1]), .o_out_fmap(xor_out[723*8*8*bW:724*8*8*bW-1]));
convchan2 c_2_724 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[724*5*5:725*5*5-1]), .o_out_fmap(xor_out[724*8*8*bW:725*8*8*bW-1]));
convchan2 c_2_725 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[725*5*5:726*5*5-1]), .o_out_fmap(xor_out[725*8*8*bW:726*8*8*bW-1]));
convchan2 c_2_726 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[726*5*5:727*5*5-1]), .o_out_fmap(xor_out[726*8*8*bW:727*8*8*bW-1]));
convchan2 c_2_727 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[727*5*5:728*5*5-1]), .o_out_fmap(xor_out[727*8*8*bW:728*8*8*bW-1]));
convchan2 c_2_728 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[728*5*5:729*5*5-1]), .o_out_fmap(xor_out[728*8*8*bW:729*8*8*bW-1]));
convchan2 c_2_729 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[729*5*5:730*5*5-1]), .o_out_fmap(xor_out[729*8*8*bW:730*8*8*bW-1]));
convchan2 c_2_730 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[730*5*5:731*5*5-1]), .o_out_fmap(xor_out[730*8*8*bW:731*8*8*bW-1]));
convchan2 c_2_731 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[731*5*5:732*5*5-1]), .o_out_fmap(xor_out[731*8*8*bW:732*8*8*bW-1]));
convchan2 c_2_732 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[732*5*5:733*5*5-1]), .o_out_fmap(xor_out[732*8*8*bW:733*8*8*bW-1]));
convchan2 c_2_733 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[733*5*5:734*5*5-1]), .o_out_fmap(xor_out[733*8*8*bW:734*8*8*bW-1]));
convchan2 c_2_734 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[734*5*5:735*5*5-1]), .o_out_fmap(xor_out[734*8*8*bW:735*8*8*bW-1]));
convchan2 c_2_735 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[735*5*5:736*5*5-1]), .o_out_fmap(xor_out[735*8*8*bW:736*8*8*bW-1]));
convchan2 c_2_736 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[736*5*5:737*5*5-1]), .o_out_fmap(xor_out[736*8*8*bW:737*8*8*bW-1]));
convchan2 c_2_737 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[737*5*5:738*5*5-1]), .o_out_fmap(xor_out[737*8*8*bW:738*8*8*bW-1]));
convchan2 c_2_738 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[738*5*5:739*5*5-1]), .o_out_fmap(xor_out[738*8*8*bW:739*8*8*bW-1]));
convchan2 c_2_739 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[739*5*5:740*5*5-1]), .o_out_fmap(xor_out[739*8*8*bW:740*8*8*bW-1]));
convchan2 c_2_740 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[740*5*5:741*5*5-1]), .o_out_fmap(xor_out[740*8*8*bW:741*8*8*bW-1]));
convchan2 c_2_741 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[741*5*5:742*5*5-1]), .o_out_fmap(xor_out[741*8*8*bW:742*8*8*bW-1]));
convchan2 c_2_742 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[742*5*5:743*5*5-1]), .o_out_fmap(xor_out[742*8*8*bW:743*8*8*bW-1]));
convchan2 c_2_743 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[743*5*5:744*5*5-1]), .o_out_fmap(xor_out[743*8*8*bW:744*8*8*bW-1]));
convchan2 c_2_744 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[744*5*5:745*5*5-1]), .o_out_fmap(xor_out[744*8*8*bW:745*8*8*bW-1]));
convchan2 c_2_745 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[745*5*5:746*5*5-1]), .o_out_fmap(xor_out[745*8*8*bW:746*8*8*bW-1]));
convchan2 c_2_746 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[746*5*5:747*5*5-1]), .o_out_fmap(xor_out[746*8*8*bW:747*8*8*bW-1]));
convchan2 c_2_747 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[747*5*5:748*5*5-1]), .o_out_fmap(xor_out[747*8*8*bW:748*8*8*bW-1]));
convchan2 c_2_748 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[748*5*5:749*5*5-1]), .o_out_fmap(xor_out[748*8*8*bW:749*8*8*bW-1]));
convchan2 c_2_749 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[749*5*5:750*5*5-1]), .o_out_fmap(xor_out[749*8*8*bW:750*8*8*bW-1]));
convchan2 c_2_750 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[750*5*5:751*5*5-1]), .o_out_fmap(xor_out[750*8*8*bW:751*8*8*bW-1]));
convchan2 c_2_751 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[751*5*5:752*5*5-1]), .o_out_fmap(xor_out[751*8*8*bW:752*8*8*bW-1]));
convchan2 c_2_752 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[752*5*5:753*5*5-1]), .o_out_fmap(xor_out[752*8*8*bW:753*8*8*bW-1]));
convchan2 c_2_753 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[753*5*5:754*5*5-1]), .o_out_fmap(xor_out[753*8*8*bW:754*8*8*bW-1]));
convchan2 c_2_754 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[754*5*5:755*5*5-1]), .o_out_fmap(xor_out[754*8*8*bW:755*8*8*bW-1]));
convchan2 c_2_755 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[755*5*5:756*5*5-1]), .o_out_fmap(xor_out[755*8*8*bW:756*8*8*bW-1]));
convchan2 c_2_756 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[756*5*5:757*5*5-1]), .o_out_fmap(xor_out[756*8*8*bW:757*8*8*bW-1]));
convchan2 c_2_757 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[757*5*5:758*5*5-1]), .o_out_fmap(xor_out[757*8*8*bW:758*8*8*bW-1]));
convchan2 c_2_758 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[758*5*5:759*5*5-1]), .o_out_fmap(xor_out[758*8*8*bW:759*8*8*bW-1]));
convchan2 c_2_759 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[759*5*5:760*5*5-1]), .o_out_fmap(xor_out[759*8*8*bW:760*8*8*bW-1]));
convchan2 c_2_760 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[760*5*5:761*5*5-1]), .o_out_fmap(xor_out[760*8*8*bW:761*8*8*bW-1]));
convchan2 c_2_761 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[761*5*5:762*5*5-1]), .o_out_fmap(xor_out[761*8*8*bW:762*8*8*bW-1]));
convchan2 c_2_762 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[762*5*5:763*5*5-1]), .o_out_fmap(xor_out[762*8*8*bW:763*8*8*bW-1]));
convchan2 c_2_763 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[763*5*5:764*5*5-1]), .o_out_fmap(xor_out[763*8*8*bW:764*8*8*bW-1]));
convchan2 c_2_764 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[764*5*5:765*5*5-1]), .o_out_fmap(xor_out[764*8*8*bW:765*8*8*bW-1]));
convchan2 c_2_765 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[765*5*5:766*5*5-1]), .o_out_fmap(xor_out[765*8*8*bW:766*8*8*bW-1]));
convchan2 c_2_766 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[766*5*5:767*5*5-1]), .o_out_fmap(xor_out[766*8*8*bW:767*8*8*bW-1]));
convchan2 c_2_767 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[767*5*5:768*5*5-1]), .o_out_fmap(xor_out[767*8*8*bW:768*8*8*bW-1]));
convchan2 c_2_768 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[768*5*5:769*5*5-1]), .o_out_fmap(xor_out[768*8*8*bW:769*8*8*bW-1]));
convchan2 c_2_769 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[769*5*5:770*5*5-1]), .o_out_fmap(xor_out[769*8*8*bW:770*8*8*bW-1]));
convchan2 c_2_770 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[770*5*5:771*5*5-1]), .o_out_fmap(xor_out[770*8*8*bW:771*8*8*bW-1]));
convchan2 c_2_771 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[771*5*5:772*5*5-1]), .o_out_fmap(xor_out[771*8*8*bW:772*8*8*bW-1]));
convchan2 c_2_772 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[772*5*5:773*5*5-1]), .o_out_fmap(xor_out[772*8*8*bW:773*8*8*bW-1]));
convchan2 c_2_773 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[773*5*5:774*5*5-1]), .o_out_fmap(xor_out[773*8*8*bW:774*8*8*bW-1]));
convchan2 c_2_774 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[774*5*5:775*5*5-1]), .o_out_fmap(xor_out[774*8*8*bW:775*8*8*bW-1]));
convchan2 c_2_775 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[775*5*5:776*5*5-1]), .o_out_fmap(xor_out[775*8*8*bW:776*8*8*bW-1]));
convchan2 c_2_776 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[776*5*5:777*5*5-1]), .o_out_fmap(xor_out[776*8*8*bW:777*8*8*bW-1]));
convchan2 c_2_777 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[777*5*5:778*5*5-1]), .o_out_fmap(xor_out[777*8*8*bW:778*8*8*bW-1]));
convchan2 c_2_778 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[778*5*5:779*5*5-1]), .o_out_fmap(xor_out[778*8*8*bW:779*8*8*bW-1]));
convchan2 c_2_779 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[779*5*5:780*5*5-1]), .o_out_fmap(xor_out[779*8*8*bW:780*8*8*bW-1]));
convchan2 c_2_780 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[780*5*5:781*5*5-1]), .o_out_fmap(xor_out[780*8*8*bW:781*8*8*bW-1]));
convchan2 c_2_781 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[781*5*5:782*5*5-1]), .o_out_fmap(xor_out[781*8*8*bW:782*8*8*bW-1]));
convchan2 c_2_782 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[782*5*5:783*5*5-1]), .o_out_fmap(xor_out[782*8*8*bW:783*8*8*bW-1]));
convchan2 c_2_783 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[783*5*5:784*5*5-1]), .o_out_fmap(xor_out[783*8*8*bW:784*8*8*bW-1]));
convchan2 c_2_784 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[784*5*5:785*5*5-1]), .o_out_fmap(xor_out[784*8*8*bW:785*8*8*bW-1]));
convchan2 c_2_785 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[785*5*5:786*5*5-1]), .o_out_fmap(xor_out[785*8*8*bW:786*8*8*bW-1]));
convchan2 c_2_786 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[786*5*5:787*5*5-1]), .o_out_fmap(xor_out[786*8*8*bW:787*8*8*bW-1]));
convchan2 c_2_787 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[787*5*5:788*5*5-1]), .o_out_fmap(xor_out[787*8*8*bW:788*8*8*bW-1]));
convchan2 c_2_788 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[788*5*5:789*5*5-1]), .o_out_fmap(xor_out[788*8*8*bW:789*8*8*bW-1]));
convchan2 c_2_789 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[789*5*5:790*5*5-1]), .o_out_fmap(xor_out[789*8*8*bW:790*8*8*bW-1]));
convchan2 c_2_790 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[790*5*5:791*5*5-1]), .o_out_fmap(xor_out[790*8*8*bW:791*8*8*bW-1]));
convchan2 c_2_791 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[791*5*5:792*5*5-1]), .o_out_fmap(xor_out[791*8*8*bW:792*8*8*bW-1]));
convchan2 c_2_792 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[792*5*5:793*5*5-1]), .o_out_fmap(xor_out[792*8*8*bW:793*8*8*bW-1]));
convchan2 c_2_793 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[793*5*5:794*5*5-1]), .o_out_fmap(xor_out[793*8*8*bW:794*8*8*bW-1]));
convchan2 c_2_794 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[794*5*5:795*5*5-1]), .o_out_fmap(xor_out[794*8*8*bW:795*8*8*bW-1]));
convchan2 c_2_795 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[795*5*5:796*5*5-1]), .o_out_fmap(xor_out[795*8*8*bW:796*8*8*bW-1]));
convchan2 c_2_796 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[796*5*5:797*5*5-1]), .o_out_fmap(xor_out[796*8*8*bW:797*8*8*bW-1]));
convchan2 c_2_797 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[797*5*5:798*5*5-1]), .o_out_fmap(xor_out[797*8*8*bW:798*8*8*bW-1]));
convchan2 c_2_798 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[798*5*5:799*5*5-1]), .o_out_fmap(xor_out[798*8*8*bW:799*8*8*bW-1]));
convchan2 c_2_799 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[799*5*5:800*5*5-1]), .o_out_fmap(xor_out[799*8*8*bW:800*8*8*bW-1]));
convchan2 c_2_800 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[800*5*5:801*5*5-1]), .o_out_fmap(xor_out[800*8*8*bW:801*8*8*bW-1]));
convchan2 c_2_801 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[801*5*5:802*5*5-1]), .o_out_fmap(xor_out[801*8*8*bW:802*8*8*bW-1]));
convchan2 c_2_802 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[802*5*5:803*5*5-1]), .o_out_fmap(xor_out[802*8*8*bW:803*8*8*bW-1]));
convchan2 c_2_803 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[803*5*5:804*5*5-1]), .o_out_fmap(xor_out[803*8*8*bW:804*8*8*bW-1]));
convchan2 c_2_804 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[804*5*5:805*5*5-1]), .o_out_fmap(xor_out[804*8*8*bW:805*8*8*bW-1]));
convchan2 c_2_805 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[805*5*5:806*5*5-1]), .o_out_fmap(xor_out[805*8*8*bW:806*8*8*bW-1]));
convchan2 c_2_806 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[806*5*5:807*5*5-1]), .o_out_fmap(xor_out[806*8*8*bW:807*8*8*bW-1]));
convchan2 c_2_807 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[807*5*5:808*5*5-1]), .o_out_fmap(xor_out[807*8*8*bW:808*8*8*bW-1]));
convchan2 c_2_808 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[808*5*5:809*5*5-1]), .o_out_fmap(xor_out[808*8*8*bW:809*8*8*bW-1]));
convchan2 c_2_809 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[809*5*5:810*5*5-1]), .o_out_fmap(xor_out[809*8*8*bW:810*8*8*bW-1]));
convchan2 c_2_810 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[810*5*5:811*5*5-1]), .o_out_fmap(xor_out[810*8*8*bW:811*8*8*bW-1]));
convchan2 c_2_811 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[811*5*5:812*5*5-1]), .o_out_fmap(xor_out[811*8*8*bW:812*8*8*bW-1]));
convchan2 c_2_812 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[812*5*5:813*5*5-1]), .o_out_fmap(xor_out[812*8*8*bW:813*8*8*bW-1]));
convchan2 c_2_813 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[813*5*5:814*5*5-1]), .o_out_fmap(xor_out[813*8*8*bW:814*8*8*bW-1]));
convchan2 c_2_814 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[814*5*5:815*5*5-1]), .o_out_fmap(xor_out[814*8*8*bW:815*8*8*bW-1]));
convchan2 c_2_815 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[815*5*5:816*5*5-1]), .o_out_fmap(xor_out[815*8*8*bW:816*8*8*bW-1]));
convchan2 c_2_816 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[816*5*5:817*5*5-1]), .o_out_fmap(xor_out[816*8*8*bW:817*8*8*bW-1]));
convchan2 c_2_817 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[817*5*5:818*5*5-1]), .o_out_fmap(xor_out[817*8*8*bW:818*8*8*bW-1]));
convchan2 c_2_818 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[818*5*5:819*5*5-1]), .o_out_fmap(xor_out[818*8*8*bW:819*8*8*bW-1]));
convchan2 c_2_819 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[819*5*5:820*5*5-1]), .o_out_fmap(xor_out[819*8*8*bW:820*8*8*bW-1]));
convchan2 c_2_820 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[820*5*5:821*5*5-1]), .o_out_fmap(xor_out[820*8*8*bW:821*8*8*bW-1]));
convchan2 c_2_821 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[821*5*5:822*5*5-1]), .o_out_fmap(xor_out[821*8*8*bW:822*8*8*bW-1]));
convchan2 c_2_822 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[822*5*5:823*5*5-1]), .o_out_fmap(xor_out[822*8*8*bW:823*8*8*bW-1]));
convchan2 c_2_823 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[823*5*5:824*5*5-1]), .o_out_fmap(xor_out[823*8*8*bW:824*8*8*bW-1]));
convchan2 c_2_824 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[824*5*5:825*5*5-1]), .o_out_fmap(xor_out[824*8*8*bW:825*8*8*bW-1]));
convchan2 c_2_825 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[825*5*5:826*5*5-1]), .o_out_fmap(xor_out[825*8*8*bW:826*8*8*bW-1]));
convchan2 c_2_826 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[826*5*5:827*5*5-1]), .o_out_fmap(xor_out[826*8*8*bW:827*8*8*bW-1]));
convchan2 c_2_827 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[827*5*5:828*5*5-1]), .o_out_fmap(xor_out[827*8*8*bW:828*8*8*bW-1]));
convchan2 c_2_828 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[828*5*5:829*5*5-1]), .o_out_fmap(xor_out[828*8*8*bW:829*8*8*bW-1]));
convchan2 c_2_829 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[829*5*5:830*5*5-1]), .o_out_fmap(xor_out[829*8*8*bW:830*8*8*bW-1]));
convchan2 c_2_830 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[830*5*5:831*5*5-1]), .o_out_fmap(xor_out[830*8*8*bW:831*8*8*bW-1]));
convchan2 c_2_831 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[831*5*5:832*5*5-1]), .o_out_fmap(xor_out[831*8*8*bW:832*8*8*bW-1]));
convchan2 c_2_832 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[832*5*5:833*5*5-1]), .o_out_fmap(xor_out[832*8*8*bW:833*8*8*bW-1]));
convchan2 c_2_833 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[833*5*5:834*5*5-1]), .o_out_fmap(xor_out[833*8*8*bW:834*8*8*bW-1]));
convchan2 c_2_834 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[834*5*5:835*5*5-1]), .o_out_fmap(xor_out[834*8*8*bW:835*8*8*bW-1]));
convchan2 c_2_835 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[835*5*5:836*5*5-1]), .o_out_fmap(xor_out[835*8*8*bW:836*8*8*bW-1]));
convchan2 c_2_836 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[836*5*5:837*5*5-1]), .o_out_fmap(xor_out[836*8*8*bW:837*8*8*bW-1]));
convchan2 c_2_837 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[837*5*5:838*5*5-1]), .o_out_fmap(xor_out[837*8*8*bW:838*8*8*bW-1]));
convchan2 c_2_838 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[838*5*5:839*5*5-1]), .o_out_fmap(xor_out[838*8*8*bW:839*8*8*bW-1]));
convchan2 c_2_839 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[839*5*5:840*5*5-1]), .o_out_fmap(xor_out[839*8*8*bW:840*8*8*bW-1]));
convchan2 c_2_840 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[840*5*5:841*5*5-1]), .o_out_fmap(xor_out[840*8*8*bW:841*8*8*bW-1]));
convchan2 c_2_841 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[841*5*5:842*5*5-1]), .o_out_fmap(xor_out[841*8*8*bW:842*8*8*bW-1]));
convchan2 c_2_842 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[842*5*5:843*5*5-1]), .o_out_fmap(xor_out[842*8*8*bW:843*8*8*bW-1]));
convchan2 c_2_843 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[843*5*5:844*5*5-1]), .o_out_fmap(xor_out[843*8*8*bW:844*8*8*bW-1]));
convchan2 c_2_844 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[844*5*5:845*5*5-1]), .o_out_fmap(xor_out[844*8*8*bW:845*8*8*bW-1]));
convchan2 c_2_845 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[845*5*5:846*5*5-1]), .o_out_fmap(xor_out[845*8*8*bW:846*8*8*bW-1]));
convchan2 c_2_846 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[846*5*5:847*5*5-1]), .o_out_fmap(xor_out[846*8*8*bW:847*8*8*bW-1]));
convchan2 c_2_847 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[847*5*5:848*5*5-1]), .o_out_fmap(xor_out[847*8*8*bW:848*8*8*bW-1]));
convchan2 c_2_848 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[848*5*5:849*5*5-1]), .o_out_fmap(xor_out[848*8*8*bW:849*8*8*bW-1]));
convchan2 c_2_849 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[849*5*5:850*5*5-1]), .o_out_fmap(xor_out[849*8*8*bW:850*8*8*bW-1]));
convchan2 c_2_850 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[850*5*5:851*5*5-1]), .o_out_fmap(xor_out[850*8*8*bW:851*8*8*bW-1]));
convchan2 c_2_851 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[851*5*5:852*5*5-1]), .o_out_fmap(xor_out[851*8*8*bW:852*8*8*bW-1]));
convchan2 c_2_852 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[852*5*5:853*5*5-1]), .o_out_fmap(xor_out[852*8*8*bW:853*8*8*bW-1]));
convchan2 c_2_853 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[853*5*5:854*5*5-1]), .o_out_fmap(xor_out[853*8*8*bW:854*8*8*bW-1]));
convchan2 c_2_854 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[854*5*5:855*5*5-1]), .o_out_fmap(xor_out[854*8*8*bW:855*8*8*bW-1]));
convchan2 c_2_855 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[855*5*5:856*5*5-1]), .o_out_fmap(xor_out[855*8*8*bW:856*8*8*bW-1]));
convchan2 c_2_856 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[856*5*5:857*5*5-1]), .o_out_fmap(xor_out[856*8*8*bW:857*8*8*bW-1]));
convchan2 c_2_857 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[857*5*5:858*5*5-1]), .o_out_fmap(xor_out[857*8*8*bW:858*8*8*bW-1]));
convchan2 c_2_858 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[858*5*5:859*5*5-1]), .o_out_fmap(xor_out[858*8*8*bW:859*8*8*bW-1]));
convchan2 c_2_859 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[859*5*5:860*5*5-1]), .o_out_fmap(xor_out[859*8*8*bW:860*8*8*bW-1]));
convchan2 c_2_860 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[860*5*5:861*5*5-1]), .o_out_fmap(xor_out[860*8*8*bW:861*8*8*bW-1]));
convchan2 c_2_861 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[861*5*5:862*5*5-1]), .o_out_fmap(xor_out[861*8*8*bW:862*8*8*bW-1]));
convchan2 c_2_862 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[862*5*5:863*5*5-1]), .o_out_fmap(xor_out[862*8*8*bW:863*8*8*bW-1]));
convchan2 c_2_863 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[863*5*5:864*5*5-1]), .o_out_fmap(xor_out[863*8*8*bW:864*8*8*bW-1]));
convchan2 c_2_864 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[864*5*5:865*5*5-1]), .o_out_fmap(xor_out[864*8*8*bW:865*8*8*bW-1]));
convchan2 c_2_865 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[865*5*5:866*5*5-1]), .o_out_fmap(xor_out[865*8*8*bW:866*8*8*bW-1]));
convchan2 c_2_866 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[866*5*5:867*5*5-1]), .o_out_fmap(xor_out[866*8*8*bW:867*8*8*bW-1]));
convchan2 c_2_867 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[867*5*5:868*5*5-1]), .o_out_fmap(xor_out[867*8*8*bW:868*8*8*bW-1]));
convchan2 c_2_868 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[868*5*5:869*5*5-1]), .o_out_fmap(xor_out[868*8*8*bW:869*8*8*bW-1]));
convchan2 c_2_869 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[869*5*5:870*5*5-1]), .o_out_fmap(xor_out[869*8*8*bW:870*8*8*bW-1]));
convchan2 c_2_870 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[870*5*5:871*5*5-1]), .o_out_fmap(xor_out[870*8*8*bW:871*8*8*bW-1]));
convchan2 c_2_871 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[871*5*5:872*5*5-1]), .o_out_fmap(xor_out[871*8*8*bW:872*8*8*bW-1]));
convchan2 c_2_872 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[872*5*5:873*5*5-1]), .o_out_fmap(xor_out[872*8*8*bW:873*8*8*bW-1]));
convchan2 c_2_873 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[873*5*5:874*5*5-1]), .o_out_fmap(xor_out[873*8*8*bW:874*8*8*bW-1]));
convchan2 c_2_874 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[874*5*5:875*5*5-1]), .o_out_fmap(xor_out[874*8*8*bW:875*8*8*bW-1]));
convchan2 c_2_875 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[875*5*5:876*5*5-1]), .o_out_fmap(xor_out[875*8*8*bW:876*8*8*bW-1]));
convchan2 c_2_876 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[876*5*5:877*5*5-1]), .o_out_fmap(xor_out[876*8*8*bW:877*8*8*bW-1]));
convchan2 c_2_877 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[877*5*5:878*5*5-1]), .o_out_fmap(xor_out[877*8*8*bW:878*8*8*bW-1]));
convchan2 c_2_878 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[878*5*5:879*5*5-1]), .o_out_fmap(xor_out[878*8*8*bW:879*8*8*bW-1]));
convchan2 c_2_879 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[879*5*5:880*5*5-1]), .o_out_fmap(xor_out[879*8*8*bW:880*8*8*bW-1]));
convchan2 c_2_880 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[880*5*5:881*5*5-1]), .o_out_fmap(xor_out[880*8*8*bW:881*8*8*bW-1]));
convchan2 c_2_881 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[881*5*5:882*5*5-1]), .o_out_fmap(xor_out[881*8*8*bW:882*8*8*bW-1]));
convchan2 c_2_882 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[882*5*5:883*5*5-1]), .o_out_fmap(xor_out[882*8*8*bW:883*8*8*bW-1]));
convchan2 c_2_883 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[883*5*5:884*5*5-1]), .o_out_fmap(xor_out[883*8*8*bW:884*8*8*bW-1]));
convchan2 c_2_884 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[884*5*5:885*5*5-1]), .o_out_fmap(xor_out[884*8*8*bW:885*8*8*bW-1]));
convchan2 c_2_885 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[885*5*5:886*5*5-1]), .o_out_fmap(xor_out[885*8*8*bW:886*8*8*bW-1]));
convchan2 c_2_886 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[886*5*5:887*5*5-1]), .o_out_fmap(xor_out[886*8*8*bW:887*8*8*bW-1]));
convchan2 c_2_887 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[887*5*5:888*5*5-1]), .o_out_fmap(xor_out[887*8*8*bW:888*8*8*bW-1]));
convchan2 c_2_888 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[888*5*5:889*5*5-1]), .o_out_fmap(xor_out[888*8*8*bW:889*8*8*bW-1]));
convchan2 c_2_889 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[889*5*5:890*5*5-1]), .o_out_fmap(xor_out[889*8*8*bW:890*8*8*bW-1]));
convchan2 c_2_890 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[890*5*5:891*5*5-1]), .o_out_fmap(xor_out[890*8*8*bW:891*8*8*bW-1]));
convchan2 c_2_891 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[891*5*5:892*5*5-1]), .o_out_fmap(xor_out[891*8*8*bW:892*8*8*bW-1]));
convchan2 c_2_892 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[892*5*5:893*5*5-1]), .o_out_fmap(xor_out[892*8*8*bW:893*8*8*bW-1]));
convchan2 c_2_893 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[893*5*5:894*5*5-1]), .o_out_fmap(xor_out[893*8*8*bW:894*8*8*bW-1]));
convchan2 c_2_894 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[894*5*5:895*5*5-1]), .o_out_fmap(xor_out[894*8*8*bW:895*8*8*bW-1]));
convchan2 c_2_895 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[895*5*5:896*5*5-1]), .o_out_fmap(xor_out[895*8*8*bW:896*8*8*bW-1]));
convchan2 c_2_896 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[896*5*5:897*5*5-1]), .o_out_fmap(xor_out[896*8*8*bW:897*8*8*bW-1]));
convchan2 c_2_897 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[897*5*5:898*5*5-1]), .o_out_fmap(xor_out[897*8*8*bW:898*8*8*bW-1]));
convchan2 c_2_898 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[898*5*5:899*5*5-1]), .o_out_fmap(xor_out[898*8*8*bW:899*8*8*bW-1]));
convchan2 c_2_899 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[899*5*5:900*5*5-1]), .o_out_fmap(xor_out[899*8*8*bW:900*8*8*bW-1]));
convchan2 c_2_900 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[900*5*5:901*5*5-1]), .o_out_fmap(xor_out[900*8*8*bW:901*8*8*bW-1]));
convchan2 c_2_901 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[901*5*5:902*5*5-1]), .o_out_fmap(xor_out[901*8*8*bW:902*8*8*bW-1]));
convchan2 c_2_902 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[902*5*5:903*5*5-1]), .o_out_fmap(xor_out[902*8*8*bW:903*8*8*bW-1]));
convchan2 c_2_903 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[903*5*5:904*5*5-1]), .o_out_fmap(xor_out[903*8*8*bW:904*8*8*bW-1]));
convchan2 c_2_904 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[904*5*5:905*5*5-1]), .o_out_fmap(xor_out[904*8*8*bW:905*8*8*bW-1]));
convchan2 c_2_905 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[905*5*5:906*5*5-1]), .o_out_fmap(xor_out[905*8*8*bW:906*8*8*bW-1]));
convchan2 c_2_906 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[906*5*5:907*5*5-1]), .o_out_fmap(xor_out[906*8*8*bW:907*8*8*bW-1]));
convchan2 c_2_907 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[907*5*5:908*5*5-1]), .o_out_fmap(xor_out[907*8*8*bW:908*8*8*bW-1]));
convchan2 c_2_908 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[908*5*5:909*5*5-1]), .o_out_fmap(xor_out[908*8*8*bW:909*8*8*bW-1]));
convchan2 c_2_909 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[909*5*5:910*5*5-1]), .o_out_fmap(xor_out[909*8*8*bW:910*8*8*bW-1]));
convchan2 c_2_910 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[910*5*5:911*5*5-1]), .o_out_fmap(xor_out[910*8*8*bW:911*8*8*bW-1]));
convchan2 c_2_911 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[911*5*5:912*5*5-1]), .o_out_fmap(xor_out[911*8*8*bW:912*8*8*bW-1]));
convchan2 c_2_912 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[912*5*5:913*5*5-1]), .o_out_fmap(xor_out[912*8*8*bW:913*8*8*bW-1]));
convchan2 c_2_913 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[913*5*5:914*5*5-1]), .o_out_fmap(xor_out[913*8*8*bW:914*8*8*bW-1]));
convchan2 c_2_914 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[914*5*5:915*5*5-1]), .o_out_fmap(xor_out[914*8*8*bW:915*8*8*bW-1]));
convchan2 c_2_915 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[915*5*5:916*5*5-1]), .o_out_fmap(xor_out[915*8*8*bW:916*8*8*bW-1]));
convchan2 c_2_916 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[916*5*5:917*5*5-1]), .o_out_fmap(xor_out[916*8*8*bW:917*8*8*bW-1]));
convchan2 c_2_917 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[917*5*5:918*5*5-1]), .o_out_fmap(xor_out[917*8*8*bW:918*8*8*bW-1]));
convchan2 c_2_918 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[918*5*5:919*5*5-1]), .o_out_fmap(xor_out[918*8*8*bW:919*8*8*bW-1]));
convchan2 c_2_919 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[919*5*5:920*5*5-1]), .o_out_fmap(xor_out[919*8*8*bW:920*8*8*bW-1]));
convchan2 c_2_920 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[920*5*5:921*5*5-1]), .o_out_fmap(xor_out[920*8*8*bW:921*8*8*bW-1]));
convchan2 c_2_921 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[921*5*5:922*5*5-1]), .o_out_fmap(xor_out[921*8*8*bW:922*8*8*bW-1]));
convchan2 c_2_922 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[922*5*5:923*5*5-1]), .o_out_fmap(xor_out[922*8*8*bW:923*8*8*bW-1]));
convchan2 c_2_923 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[923*5*5:924*5*5-1]), .o_out_fmap(xor_out[923*8*8*bW:924*8*8*bW-1]));
convchan2 c_2_924 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[924*5*5:925*5*5-1]), .o_out_fmap(xor_out[924*8*8*bW:925*8*8*bW-1]));
convchan2 c_2_925 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[925*5*5:926*5*5-1]), .o_out_fmap(xor_out[925*8*8*bW:926*8*8*bW-1]));
convchan2 c_2_926 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[926*5*5:927*5*5-1]), .o_out_fmap(xor_out[926*8*8*bW:927*8*8*bW-1]));
convchan2 c_2_927 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[927*5*5:928*5*5-1]), .o_out_fmap(xor_out[927*8*8*bW:928*8*8*bW-1]));
convchan2 c_2_928 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[928*5*5:929*5*5-1]), .o_out_fmap(xor_out[928*8*8*bW:929*8*8*bW-1]));
convchan2 c_2_929 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[929*5*5:930*5*5-1]), .o_out_fmap(xor_out[929*8*8*bW:930*8*8*bW-1]));
convchan2 c_2_930 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[930*5*5:931*5*5-1]), .o_out_fmap(xor_out[930*8*8*bW:931*8*8*bW-1]));
convchan2 c_2_931 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[931*5*5:932*5*5-1]), .o_out_fmap(xor_out[931*8*8*bW:932*8*8*bW-1]));
convchan2 c_2_932 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[932*5*5:933*5*5-1]), .o_out_fmap(xor_out[932*8*8*bW:933*8*8*bW-1]));
convchan2 c_2_933 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[933*5*5:934*5*5-1]), .o_out_fmap(xor_out[933*8*8*bW:934*8*8*bW-1]));
convchan2 c_2_934 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[934*5*5:935*5*5-1]), .o_out_fmap(xor_out[934*8*8*bW:935*8*8*bW-1]));
convchan2 c_2_935 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[935*5*5:936*5*5-1]), .o_out_fmap(xor_out[935*8*8*bW:936*8*8*bW-1]));
convchan2 c_2_936 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[936*5*5:937*5*5-1]), .o_out_fmap(xor_out[936*8*8*bW:937*8*8*bW-1]));
convchan2 c_2_937 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[937*5*5:938*5*5-1]), .o_out_fmap(xor_out[937*8*8*bW:938*8*8*bW-1]));
convchan2 c_2_938 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[938*5*5:939*5*5-1]), .o_out_fmap(xor_out[938*8*8*bW:939*8*8*bW-1]));
convchan2 c_2_939 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[939*5*5:940*5*5-1]), .o_out_fmap(xor_out[939*8*8*bW:940*8*8*bW-1]));
convchan2 c_2_940 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[940*5*5:941*5*5-1]), .o_out_fmap(xor_out[940*8*8*bW:941*8*8*bW-1]));
convchan2 c_2_941 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[941*5*5:942*5*5-1]), .o_out_fmap(xor_out[941*8*8*bW:942*8*8*bW-1]));
convchan2 c_2_942 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[942*5*5:943*5*5-1]), .o_out_fmap(xor_out[942*8*8*bW:943*8*8*bW-1]));
convchan2 c_2_943 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[943*5*5:944*5*5-1]), .o_out_fmap(xor_out[943*8*8*bW:944*8*8*bW-1]));
convchan2 c_2_944 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[944*5*5:945*5*5-1]), .o_out_fmap(xor_out[944*8*8*bW:945*8*8*bW-1]));
convchan2 c_2_945 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[945*5*5:946*5*5-1]), .o_out_fmap(xor_out[945*8*8*bW:946*8*8*bW-1]));
convchan2 c_2_946 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[946*5*5:947*5*5-1]), .o_out_fmap(xor_out[946*8*8*bW:947*8*8*bW-1]));
convchan2 c_2_947 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[947*5*5:948*5*5-1]), .o_out_fmap(xor_out[947*8*8*bW:948*8*8*bW-1]));
convchan2 c_2_948 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[948*5*5:949*5*5-1]), .o_out_fmap(xor_out[948*8*8*bW:949*8*8*bW-1]));
convchan2 c_2_949 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[949*5*5:950*5*5-1]), .o_out_fmap(xor_out[949*8*8*bW:950*8*8*bW-1]));
convchan2 c_2_950 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[950*5*5:951*5*5-1]), .o_out_fmap(xor_out[950*8*8*bW:951*8*8*bW-1]));
convchan2 c_2_951 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[951*5*5:952*5*5-1]), .o_out_fmap(xor_out[951*8*8*bW:952*8*8*bW-1]));
convchan2 c_2_952 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[952*5*5:953*5*5-1]), .o_out_fmap(xor_out[952*8*8*bW:953*8*8*bW-1]));
convchan2 c_2_953 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[953*5*5:954*5*5-1]), .o_out_fmap(xor_out[953*8*8*bW:954*8*8*bW-1]));
convchan2 c_2_954 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[954*5*5:955*5*5-1]), .o_out_fmap(xor_out[954*8*8*bW:955*8*8*bW-1]));
convchan2 c_2_955 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[955*5*5:956*5*5-1]), .o_out_fmap(xor_out[955*8*8*bW:956*8*8*bW-1]));
convchan2 c_2_956 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[956*5*5:957*5*5-1]), .o_out_fmap(xor_out[956*8*8*bW:957*8*8*bW-1]));
convchan2 c_2_957 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[957*5*5:958*5*5-1]), .o_out_fmap(xor_out[957*8*8*bW:958*8*8*bW-1]));
convchan2 c_2_958 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[958*5*5:959*5*5-1]), .o_out_fmap(xor_out[958*8*8*bW:959*8*8*bW-1]));
convchan2 c_2_959 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[959*5*5:960*5*5-1]), .o_out_fmap(xor_out[959*8*8*bW:960*8*8*bW-1]));
convchan2 c_2_960 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[960*5*5:961*5*5-1]), .o_out_fmap(xor_out[960*8*8*bW:961*8*8*bW-1]));
convchan2 c_2_961 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[961*5*5:962*5*5-1]), .o_out_fmap(xor_out[961*8*8*bW:962*8*8*bW-1]));
convchan2 c_2_962 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[962*5*5:963*5*5-1]), .o_out_fmap(xor_out[962*8*8*bW:963*8*8*bW-1]));
convchan2 c_2_963 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[963*5*5:964*5*5-1]), .o_out_fmap(xor_out[963*8*8*bW:964*8*8*bW-1]));
convchan2 c_2_964 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[964*5*5:965*5*5-1]), .o_out_fmap(xor_out[964*8*8*bW:965*8*8*bW-1]));
convchan2 c_2_965 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[965*5*5:966*5*5-1]), .o_out_fmap(xor_out[965*8*8*bW:966*8*8*bW-1]));
convchan2 c_2_966 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[966*5*5:967*5*5-1]), .o_out_fmap(xor_out[966*8*8*bW:967*8*8*bW-1]));
convchan2 c_2_967 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[967*5*5:968*5*5-1]), .o_out_fmap(xor_out[967*8*8*bW:968*8*8*bW-1]));
convchan2 c_2_968 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[968*5*5:969*5*5-1]), .o_out_fmap(xor_out[968*8*8*bW:969*8*8*bW-1]));
convchan2 c_2_969 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[969*5*5:970*5*5-1]), .o_out_fmap(xor_out[969*8*8*bW:970*8*8*bW-1]));
convchan2 c_2_970 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[970*5*5:971*5*5-1]), .o_out_fmap(xor_out[970*8*8*bW:971*8*8*bW-1]));
convchan2 c_2_971 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[971*5*5:972*5*5-1]), .o_out_fmap(xor_out[971*8*8*bW:972*8*8*bW-1]));
convchan2 c_2_972 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[972*5*5:973*5*5-1]), .o_out_fmap(xor_out[972*8*8*bW:973*8*8*bW-1]));
convchan2 c_2_973 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[973*5*5:974*5*5-1]), .o_out_fmap(xor_out[973*8*8*bW:974*8*8*bW-1]));
convchan2 c_2_974 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[974*5*5:975*5*5-1]), .o_out_fmap(xor_out[974*8*8*bW:975*8*8*bW-1]));
convchan2 c_2_975 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[975*5*5:976*5*5-1]), .o_out_fmap(xor_out[975*8*8*bW:976*8*8*bW-1]));
convchan2 c_2_976 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[976*5*5:977*5*5-1]), .o_out_fmap(xor_out[976*8*8*bW:977*8*8*bW-1]));
convchan2 c_2_977 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[977*5*5:978*5*5-1]), .o_out_fmap(xor_out[977*8*8*bW:978*8*8*bW-1]));
convchan2 c_2_978 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[978*5*5:979*5*5-1]), .o_out_fmap(xor_out[978*8*8*bW:979*8*8*bW-1]));
convchan2 c_2_979 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[979*5*5:980*5*5-1]), .o_out_fmap(xor_out[979*8*8*bW:980*8*8*bW-1]));
convchan2 c_2_980 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[980*5*5:981*5*5-1]), .o_out_fmap(xor_out[980*8*8*bW:981*8*8*bW-1]));
convchan2 c_2_981 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[981*5*5:982*5*5-1]), .o_out_fmap(xor_out[981*8*8*bW:982*8*8*bW-1]));
convchan2 c_2_982 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[982*5*5:983*5*5-1]), .o_out_fmap(xor_out[982*8*8*bW:983*8*8*bW-1]));
convchan2 c_2_983 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[983*5*5:984*5*5-1]), .o_out_fmap(xor_out[983*8*8*bW:984*8*8*bW-1]));
convchan2 c_2_984 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[984*5*5:985*5*5-1]), .o_out_fmap(xor_out[984*8*8*bW:985*8*8*bW-1]));
convchan2 c_2_985 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[985*5*5:986*5*5-1]), .o_out_fmap(xor_out[985*8*8*bW:986*8*8*bW-1]));
convchan2 c_2_986 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[986*5*5:987*5*5-1]), .o_out_fmap(xor_out[986*8*8*bW:987*8*8*bW-1]));
convchan2 c_2_987 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[987*5*5:988*5*5-1]), .o_out_fmap(xor_out[987*8*8*bW:988*8*8*bW-1]));
convchan2 c_2_988 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[988*5*5:989*5*5-1]), .o_out_fmap(xor_out[988*8*8*bW:989*8*8*bW-1]));
convchan2 c_2_989 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[989*5*5:990*5*5-1]), .o_out_fmap(xor_out[989*8*8*bW:990*8*8*bW-1]));
convchan2 c_2_990 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[990*5*5:991*5*5-1]), .o_out_fmap(xor_out[990*8*8*bW:991*8*8*bW-1]));
convchan2 c_2_991 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[991*5*5:992*5*5-1]), .o_out_fmap(xor_out[991*8*8*bW:992*8*8*bW-1]));
convchan2 c_2_992 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[992*5*5:993*5*5-1]), .o_out_fmap(xor_out[992*8*8*bW:993*8*8*bW-1]));
convchan2 c_2_993 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[993*5*5:994*5*5-1]), .o_out_fmap(xor_out[993*8*8*bW:994*8*8*bW-1]));
convchan2 c_2_994 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[994*5*5:995*5*5-1]), .o_out_fmap(xor_out[994*8*8*bW:995*8*8*bW-1]));
convchan2 c_2_995 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[995*5*5:996*5*5-1]), .o_out_fmap(xor_out[995*8*8*bW:996*8*8*bW-1]));
convchan2 c_2_996 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[996*5*5:997*5*5-1]), .o_out_fmap(xor_out[996*8*8*bW:997*8*8*bW-1]));
convchan2 c_2_997 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[997*5*5:998*5*5-1]), .o_out_fmap(xor_out[997*8*8*bW:998*8*8*bW-1]));
convchan2 c_2_998 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[998*5*5:999*5*5-1]), .o_out_fmap(xor_out[998*8*8*bW:999*8*8*bW-1]));
convchan2 c_2_999 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[999*5*5:1000*5*5-1]), .o_out_fmap(xor_out[999*8*8*bW:1000*8*8*bW-1]));
convchan2 c_2_1000 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[1000*5*5:1001*5*5-1]), .o_out_fmap(xor_out[1000*8*8*bW:1001*8*8*bW-1]));
convchan2 c_2_1001 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[1001*5*5:1002*5*5-1]), .o_out_fmap(xor_out[1001*8*8*bW:1002*8*8*bW-1]));
convchan2 c_2_1002 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[1002*5*5:1003*5*5-1]), .o_out_fmap(xor_out[1002*8*8*bW:1003*8*8*bW-1]));
convchan2 c_2_1003 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[1003*5*5:1004*5*5-1]), .o_out_fmap(xor_out[1003*8*8*bW:1004*8*8*bW-1]));
convchan2 c_2_1004 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[1004*5*5:1005*5*5-1]), .o_out_fmap(xor_out[1004*8*8*bW:1005*8*8*bW-1]));
convchan2 c_2_1005 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[1005*5*5:1006*5*5-1]), .o_out_fmap(xor_out[1005*8*8*bW:1006*8*8*bW-1]));
convchan2 c_2_1006 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[1006*5*5:1007*5*5-1]), .o_out_fmap(xor_out[1006*8*8*bW:1007*8*8*bW-1]));
convchan2 c_2_1007 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[1007*5*5:1008*5*5-1]), .o_out_fmap(xor_out[1007*8*8*bW:1008*8*8*bW-1]));
convchan2 c_2_1008 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[1008*5*5:1009*5*5-1]), .o_out_fmap(xor_out[1008*8*8*bW:1009*8*8*bW-1]));
convchan2 c_2_1009 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[1009*5*5:1010*5*5-1]), .o_out_fmap(xor_out[1009*8*8*bW:1010*8*8*bW-1]));
convchan2 c_2_1010 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[1010*5*5:1011*5*5-1]), .o_out_fmap(xor_out[1010*8*8*bW:1011*8*8*bW-1]));
convchan2 c_2_1011 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[1011*5*5:1012*5*5-1]), .o_out_fmap(xor_out[1011*8*8*bW:1012*8*8*bW-1]));
convchan2 c_2_1012 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[1012*5*5:1013*5*5-1]), .o_out_fmap(xor_out[1012*8*8*bW:1013*8*8*bW-1]));
convchan2 c_2_1013 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[1013*5*5:1014*5*5-1]), .o_out_fmap(xor_out[1013*8*8*bW:1014*8*8*bW-1]));
convchan2 c_2_1014 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[1014*5*5:1015*5*5-1]), .o_out_fmap(xor_out[1014*8*8*bW:1015*8*8*bW-1]));
convchan2 c_2_1015 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[1015*5*5:1016*5*5-1]), .o_out_fmap(xor_out[1015*8*8*bW:1016*8*8*bW-1]));
convchan2 c_2_1016 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[1016*5*5:1017*5*5-1]), .o_out_fmap(xor_out[1016*8*8*bW:1017*8*8*bW-1]));
convchan2 c_2_1017 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[1017*5*5:1018*5*5-1]), .o_out_fmap(xor_out[1017*8*8*bW:1018*8*8*bW-1]));
convchan2 c_2_1018 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[1018*5*5:1019*5*5-1]), .o_out_fmap(xor_out[1018*8*8*bW:1019*8*8*bW-1]));
convchan2 c_2_1019 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[1019*5*5:1020*5*5-1]), .o_out_fmap(xor_out[1019*8*8*bW:1020*8*8*bW-1]));
convchan2 c_2_1020 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1020*5*5:1021*5*5-1]), .o_out_fmap(xor_out[1020*8*8*bW:1021*8*8*bW-1]));
convchan2 c_2_1021 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1021*5*5:1022*5*5-1]), .o_out_fmap(xor_out[1021*8*8*bW:1022*8*8*bW-1]));
convchan2 c_2_1022 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1022*5*5:1023*5*5-1]), .o_out_fmap(xor_out[1022*8*8*bW:1023*8*8*bW-1]));
convchan2 c_2_1023 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1023*5*5:1024*5*5-1]), .o_out_fmap(xor_out[1023*8*8*bW:1024*8*8*bW-1]));
convchan2 c_2_1024 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1024*5*5:1025*5*5-1]), .o_out_fmap(xor_out[1024*8*8*bW:1025*8*8*bW-1]));
convchan2 c_2_1025 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1025*5*5:1026*5*5-1]), .o_out_fmap(xor_out[1025*8*8*bW:1026*8*8*bW-1]));
convchan2 c_2_1026 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1026*5*5:1027*5*5-1]), .o_out_fmap(xor_out[1026*8*8*bW:1027*8*8*bW-1]));
convchan2 c_2_1027 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1027*5*5:1028*5*5-1]), .o_out_fmap(xor_out[1027*8*8*bW:1028*8*8*bW-1]));
convchan2 c_2_1028 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1028*5*5:1029*5*5-1]), .o_out_fmap(xor_out[1028*8*8*bW:1029*8*8*bW-1]));
convchan2 c_2_1029 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1029*5*5:1030*5*5-1]), .o_out_fmap(xor_out[1029*8*8*bW:1030*8*8*bW-1]));
convchan2 c_2_1030 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1030*5*5:1031*5*5-1]), .o_out_fmap(xor_out[1030*8*8*bW:1031*8*8*bW-1]));
convchan2 c_2_1031 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1031*5*5:1032*5*5-1]), .o_out_fmap(xor_out[1031*8*8*bW:1032*8*8*bW-1]));
convchan2 c_2_1032 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1032*5*5:1033*5*5-1]), .o_out_fmap(xor_out[1032*8*8*bW:1033*8*8*bW-1]));
convchan2 c_2_1033 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1033*5*5:1034*5*5-1]), .o_out_fmap(xor_out[1033*8*8*bW:1034*8*8*bW-1]));
convchan2 c_2_1034 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1034*5*5:1035*5*5-1]), .o_out_fmap(xor_out[1034*8*8*bW:1035*8*8*bW-1]));
convchan2 c_2_1035 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1035*5*5:1036*5*5-1]), .o_out_fmap(xor_out[1035*8*8*bW:1036*8*8*bW-1]));
convchan2 c_2_1036 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1036*5*5:1037*5*5-1]), .o_out_fmap(xor_out[1036*8*8*bW:1037*8*8*bW-1]));
convchan2 c_2_1037 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1037*5*5:1038*5*5-1]), .o_out_fmap(xor_out[1037*8*8*bW:1038*8*8*bW-1]));
convchan2 c_2_1038 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1038*5*5:1039*5*5-1]), .o_out_fmap(xor_out[1038*8*8*bW:1039*8*8*bW-1]));
convchan2 c_2_1039 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1039*5*5:1040*5*5-1]), .o_out_fmap(xor_out[1039*8*8*bW:1040*8*8*bW-1]));
convchan2 c_2_1040 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1040*5*5:1041*5*5-1]), .o_out_fmap(xor_out[1040*8*8*bW:1041*8*8*bW-1]));
convchan2 c_2_1041 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1041*5*5:1042*5*5-1]), .o_out_fmap(xor_out[1041*8*8*bW:1042*8*8*bW-1]));
convchan2 c_2_1042 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1042*5*5:1043*5*5-1]), .o_out_fmap(xor_out[1042*8*8*bW:1043*8*8*bW-1]));
convchan2 c_2_1043 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1043*5*5:1044*5*5-1]), .o_out_fmap(xor_out[1043*8*8*bW:1044*8*8*bW-1]));
convchan2 c_2_1044 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1044*5*5:1045*5*5-1]), .o_out_fmap(xor_out[1044*8*8*bW:1045*8*8*bW-1]));
convchan2 c_2_1045 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1045*5*5:1046*5*5-1]), .o_out_fmap(xor_out[1045*8*8*bW:1046*8*8*bW-1]));
convchan2 c_2_1046 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1046*5*5:1047*5*5-1]), .o_out_fmap(xor_out[1046*8*8*bW:1047*8*8*bW-1]));
convchan2 c_2_1047 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1047*5*5:1048*5*5-1]), .o_out_fmap(xor_out[1047*8*8*bW:1048*8*8*bW-1]));
convchan2 c_2_1048 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1048*5*5:1049*5*5-1]), .o_out_fmap(xor_out[1048*8*8*bW:1049*8*8*bW-1]));
convchan2 c_2_1049 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1049*5*5:1050*5*5-1]), .o_out_fmap(xor_out[1049*8*8*bW:1050*8*8*bW-1]));
convchan2 c_2_1050 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1050*5*5:1051*5*5-1]), .o_out_fmap(xor_out[1050*8*8*bW:1051*8*8*bW-1]));
convchan2 c_2_1051 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1051*5*5:1052*5*5-1]), .o_out_fmap(xor_out[1051*8*8*bW:1052*8*8*bW-1]));
convchan2 c_2_1052 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1052*5*5:1053*5*5-1]), .o_out_fmap(xor_out[1052*8*8*bW:1053*8*8*bW-1]));
convchan2 c_2_1053 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1053*5*5:1054*5*5-1]), .o_out_fmap(xor_out[1053*8*8*bW:1054*8*8*bW-1]));
convchan2 c_2_1054 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1054*5*5:1055*5*5-1]), .o_out_fmap(xor_out[1054*8*8*bW:1055*8*8*bW-1]));
convchan2 c_2_1055 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1055*5*5:1056*5*5-1]), .o_out_fmap(xor_out[1055*8*8*bW:1056*8*8*bW-1]));
convchan2 c_2_1056 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1056*5*5:1057*5*5-1]), .o_out_fmap(xor_out[1056*8*8*bW:1057*8*8*bW-1]));
convchan2 c_2_1057 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1057*5*5:1058*5*5-1]), .o_out_fmap(xor_out[1057*8*8*bW:1058*8*8*bW-1]));
convchan2 c_2_1058 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1058*5*5:1059*5*5-1]), .o_out_fmap(xor_out[1058*8*8*bW:1059*8*8*bW-1]));
convchan2 c_2_1059 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1059*5*5:1060*5*5-1]), .o_out_fmap(xor_out[1059*8*8*bW:1060*8*8*bW-1]));
convchan2 c_2_1060 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1060*5*5:1061*5*5-1]), .o_out_fmap(xor_out[1060*8*8*bW:1061*8*8*bW-1]));
convchan2 c_2_1061 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1061*5*5:1062*5*5-1]), .o_out_fmap(xor_out[1061*8*8*bW:1062*8*8*bW-1]));
convchan2 c_2_1062 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1062*5*5:1063*5*5-1]), .o_out_fmap(xor_out[1062*8*8*bW:1063*8*8*bW-1]));
convchan2 c_2_1063 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1063*5*5:1064*5*5-1]), .o_out_fmap(xor_out[1063*8*8*bW:1064*8*8*bW-1]));
convchan2 c_2_1064 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1064*5*5:1065*5*5-1]), .o_out_fmap(xor_out[1064*8*8*bW:1065*8*8*bW-1]));
convchan2 c_2_1065 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1065*5*5:1066*5*5-1]), .o_out_fmap(xor_out[1065*8*8*bW:1066*8*8*bW-1]));
convchan2 c_2_1066 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1066*5*5:1067*5*5-1]), .o_out_fmap(xor_out[1066*8*8*bW:1067*8*8*bW-1]));
convchan2 c_2_1067 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1067*5*5:1068*5*5-1]), .o_out_fmap(xor_out[1067*8*8*bW:1068*8*8*bW-1]));
convchan2 c_2_1068 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1068*5*5:1069*5*5-1]), .o_out_fmap(xor_out[1068*8*8*bW:1069*8*8*bW-1]));
convchan2 c_2_1069 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1069*5*5:1070*5*5-1]), .o_out_fmap(xor_out[1069*8*8*bW:1070*8*8*bW-1]));
convchan2 c_2_1070 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1070*5*5:1071*5*5-1]), .o_out_fmap(xor_out[1070*8*8*bW:1071*8*8*bW-1]));
convchan2 c_2_1071 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1071*5*5:1072*5*5-1]), .o_out_fmap(xor_out[1071*8*8*bW:1072*8*8*bW-1]));
convchan2 c_2_1072 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1072*5*5:1073*5*5-1]), .o_out_fmap(xor_out[1072*8*8*bW:1073*8*8*bW-1]));
convchan2 c_2_1073 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1073*5*5:1074*5*5-1]), .o_out_fmap(xor_out[1073*8*8*bW:1074*8*8*bW-1]));
convchan2 c_2_1074 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1074*5*5:1075*5*5-1]), .o_out_fmap(xor_out[1074*8*8*bW:1075*8*8*bW-1]));
convchan2 c_2_1075 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1075*5*5:1076*5*5-1]), .o_out_fmap(xor_out[1075*8*8*bW:1076*8*8*bW-1]));
convchan2 c_2_1076 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1076*5*5:1077*5*5-1]), .o_out_fmap(xor_out[1076*8*8*bW:1077*8*8*bW-1]));
convchan2 c_2_1077 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1077*5*5:1078*5*5-1]), .o_out_fmap(xor_out[1077*8*8*bW:1078*8*8*bW-1]));
convchan2 c_2_1078 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1078*5*5:1079*5*5-1]), .o_out_fmap(xor_out[1078*8*8*bW:1079*8*8*bW-1]));
convchan2 c_2_1079 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1079*5*5:1080*5*5-1]), .o_out_fmap(xor_out[1079*8*8*bW:1080*8*8*bW-1]));

endmodule