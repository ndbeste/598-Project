module conv_pool_pixel450
#(parameter chan = 18,
parameter bW = 9)
(
input logic image[0:chan-1][0:5][0:5],
input logic kernels[0:chan-1][0:5-1][0:5-1],
input logic [bW-1:0] offset,
output logic pixel);


logic [chan*5*5-1:0] image_slice1;
assign image_slice1 = {image[0][0][0],image[0][0][1],image[0][0][2],image[0][0][3],image[0][0][4],image[0][1][0],image[0][1][1],image[0][1][2],image[0][1][3],image[0][1][4],image[0][2][0],image[0][2][1],image[0][2][2],image[0][2][3],image[0][2][4],image[0][3][0],image[0][3][1],image[0][3][2],image[0][3][3],image[0][3][4],image[0][4][0],image[0][4][1],image[0][4][2],image[0][4][3],image[0][4][4],image[1][0][0],image[1][0][1],image[1][0][2],image[1][0][3],image[1][0][4],image[1][1][0],image[1][1][1],image[1][1][2],image[1][1][3],image[1][1][4],image[1][2][0],image[1][2][1],image[1][2][2],image[1][2][3],image[1][2][4],image[1][3][0],image[1][3][1],image[1][3][2],image[1][3][3],image[1][3][4],image[1][4][0],image[1][4][1],image[1][4][2],image[1][4][3],image[1][4][4],image[2][0][0],image[2][0][1],image[2][0][2],image[2][0][3],image[2][0][4],image[2][1][0],image[2][1][1],image[2][1][2],image[2][1][3],image[2][1][4],image[2][2][0],image[2][2][1],image[2][2][2],image[2][2][3],image[2][2][4],image[2][3][0],image[2][3][1],image[2][3][2],image[2][3][3],image[2][3][4],image[2][4][0],image[2][4][1],image[2][4][2],image[2][4][3],image[2][4][4],image[3][0][0],image[3][0][1],image[3][0][2],image[3][0][3],image[3][0][4],image[3][1][0],image[3][1][1],image[3][1][2],image[3][1][3],image[3][1][4],image[3][2][0],image[3][2][1],image[3][2][2],image[3][2][3],image[3][2][4],image[3][3][0],image[3][3][1],image[3][3][2],image[3][3][3],image[3][3][4],image[3][4][0],image[3][4][1],image[3][4][2],image[3][4][3],image[3][4][4],image[4][0][0],image[4][0][1],image[4][0][2],image[4][0][3],image[4][0][4],image[4][1][0],image[4][1][1],image[4][1][2],image[4][1][3],image[4][1][4],image[4][2][0],image[4][2][1],image[4][2][2],image[4][2][3],image[4][2][4],image[4][3][0],image[4][3][1],image[4][3][2],image[4][3][3],image[4][3][4],image[4][4][0],image[4][4][1],image[4][4][2],image[4][4][3],image[4][4][4],image[5][0][0],image[5][0][1],image[5][0][2],image[5][0][3],image[5][0][4],image[5][1][0],image[5][1][1],image[5][1][2],image[5][1][3],image[5][1][4],image[5][2][0],image[5][2][1],image[5][2][2],image[5][2][3],image[5][2][4],image[5][3][0],image[5][3][1],image[5][3][2],image[5][3][3],image[5][3][4],image[5][4][0],image[5][4][1],image[5][4][2],image[5][4][3],image[5][4][4],image[6][0][0],image[6][0][1],image[6][0][2],image[6][0][3],image[6][0][4],image[6][1][0],image[6][1][1],image[6][1][2],image[6][1][3],image[6][1][4],image[6][2][0],image[6][2][1],image[6][2][2],image[6][2][3],image[6][2][4],image[6][3][0],image[6][3][1],image[6][3][2],image[6][3][3],image[6][3][4],image[6][4][0],image[6][4][1],image[6][4][2],image[6][4][3],image[6][4][4],image[7][0][0],image[7][0][1],image[7][0][2],image[7][0][3],image[7][0][4],image[7][1][0],image[7][1][1],image[7][1][2],image[7][1][3],image[7][1][4],image[7][2][0],image[7][2][1],image[7][2][2],image[7][2][3],image[7][2][4],image[7][3][0],image[7][3][1],image[7][3][2],image[7][3][3],image[7][3][4],image[7][4][0],image[7][4][1],image[7][4][2],image[7][4][3],image[7][4][4],image[8][0][0],image[8][0][1],image[8][0][2],image[8][0][3],image[8][0][4],image[8][1][0],image[8][1][1],image[8][1][2],image[8][1][3],image[8][1][4],image[8][2][0],image[8][2][1],image[8][2][2],image[8][2][3],image[8][2][4],image[8][3][0],image[8][3][1],image[8][3][2],image[8][3][3],image[8][3][4],image[8][4][0],image[8][4][1],image[8][4][2],image[8][4][3],image[8][4][4],image[9][0][0],image[9][0][1],image[9][0][2],image[9][0][3],image[9][0][4],image[9][1][0],image[9][1][1],image[9][1][2],image[9][1][3],image[9][1][4],image[9][2][0],image[9][2][1],image[9][2][2],image[9][2][3],image[9][2][4],image[9][3][0],image[9][3][1],image[9][3][2],image[9][3][3],image[9][3][4],image[9][4][0],image[9][4][1],image[9][4][2],image[9][4][3],image[9][4][4],image[10][0][0],image[10][0][1],image[10][0][2],image[10][0][3],image[10][0][4],image[10][1][0],image[10][1][1],image[10][1][2],image[10][1][3],image[10][1][4],image[10][2][0],image[10][2][1],image[10][2][2],image[10][2][3],image[10][2][4],image[10][3][0],image[10][3][1],image[10][3][2],image[10][3][3],image[10][3][4],image[10][4][0],image[10][4][1],image[10][4][2],image[10][4][3],image[10][4][4],image[11][0][0],image[11][0][1],image[11][0][2],image[11][0][3],image[11][0][4],image[11][1][0],image[11][1][1],image[11][1][2],image[11][1][3],image[11][1][4],image[11][2][0],image[11][2][1],image[11][2][2],image[11][2][3],image[11][2][4],image[11][3][0],image[11][3][1],image[11][3][2],image[11][3][3],image[11][3][4],image[11][4][0],image[11][4][1],image[11][4][2],image[11][4][3],image[11][4][4],image[12][0][0],image[12][0][1],image[12][0][2],image[12][0][3],image[12][0][4],image[12][1][0],image[12][1][1],image[12][1][2],image[12][1][3],image[12][1][4],image[12][2][0],image[12][2][1],image[12][2][2],image[12][2][3],image[12][2][4],image[12][3][0],image[12][3][1],image[12][3][2],image[12][3][3],image[12][3][4],image[12][4][0],image[12][4][1],image[12][4][2],image[12][4][3],image[12][4][4],image[13][0][0],image[13][0][1],image[13][0][2],image[13][0][3],image[13][0][4],image[13][1][0],image[13][1][1],image[13][1][2],image[13][1][3],image[13][1][4],image[13][2][0],image[13][2][1],image[13][2][2],image[13][2][3],image[13][2][4],image[13][3][0],image[13][3][1],image[13][3][2],image[13][3][3],image[13][3][4],image[13][4][0],image[13][4][1],image[13][4][2],image[13][4][3],image[13][4][4],image[14][0][0],image[14][0][1],image[14][0][2],image[14][0][3],image[14][0][4],image[14][1][0],image[14][1][1],image[14][1][2],image[14][1][3],image[14][1][4],image[14][2][0],image[14][2][1],image[14][2][2],image[14][2][3],image[14][2][4],image[14][3][0],image[14][3][1],image[14][3][2],image[14][3][3],image[14][3][4],image[14][4][0],image[14][4][1],image[14][4][2],image[14][4][3],image[14][4][4],image[15][0][0],image[15][0][1],image[15][0][2],image[15][0][3],image[15][0][4],image[15][1][0],image[15][1][1],image[15][1][2],image[15][1][3],image[15][1][4],image[15][2][0],image[15][2][1],image[15][2][2],image[15][2][3],image[15][2][4],image[15][3][0],image[15][3][1],image[15][3][2],image[15][3][3],image[15][3][4],image[15][4][0],image[15][4][1],image[15][4][2],image[15][4][3],image[15][4][4],image[16][0][0],image[16][0][1],image[16][0][2],image[16][0][3],image[16][0][4],image[16][1][0],image[16][1][1],image[16][1][2],image[16][1][3],image[16][1][4],image[16][2][0],image[16][2][1],image[16][2][2],image[16][2][3],image[16][2][4],image[16][3][0],image[16][3][1],image[16][3][2],image[16][3][3],image[16][3][4],image[16][4][0],image[16][4][1],image[16][4][2],image[16][4][3],image[16][4][4],image[17][0][0],image[17][0][1],image[17][0][2],image[17][0][3],image[17][0][4],image[17][1][0],image[17][1][1],image[17][1][2],image[17][1][3],image[17][1][4],image[17][2][0],image[17][2][1],image[17][2][2],image[17][2][3],image[17][2][4],image[17][3][0],image[17][3][1],image[17][3][2],image[17][3][3],image[17][3][4],image[17][4][0],image[17][4][1],image[17][4][2],image[17][4][3],image[17][4][4]};
logic [chan*5*5-1:0] image_slice2;
assign image_slice2 = {image[0][1][0],image[0][1][1],image[0][1][2],image[0][1][3],image[0][1][4],image[0][2][0],image[0][2][1],image[0][2][2],image[0][2][3],image[0][2][4],image[0][3][0],image[0][3][1],image[0][3][2],image[0][3][3],image[0][3][4],image[0][4][0],image[0][4][1],image[0][4][2],image[0][4][3],image[0][4][4],image[0][5][0],image[0][5][1],image[0][5][2],image[0][5][3],image[0][5][4],image[1][1][0],image[1][1][1],image[1][1][2],image[1][1][3],image[1][1][4],image[1][2][0],image[1][2][1],image[1][2][2],image[1][2][3],image[1][2][4],image[1][3][0],image[1][3][1],image[1][3][2],image[1][3][3],image[1][3][4],image[1][4][0],image[1][4][1],image[1][4][2],image[1][4][3],image[1][4][4],image[1][5][0],image[1][5][1],image[1][5][2],image[1][5][3],image[1][5][4],image[2][1][0],image[2][1][1],image[2][1][2],image[2][1][3],image[2][1][4],image[2][2][0],image[2][2][1],image[2][2][2],image[2][2][3],image[2][2][4],image[2][3][0],image[2][3][1],image[2][3][2],image[2][3][3],image[2][3][4],image[2][4][0],image[2][4][1],image[2][4][2],image[2][4][3],image[2][4][4],image[2][5][0],image[2][5][1],image[2][5][2],image[2][5][3],image[2][5][4],image[3][1][0],image[3][1][1],image[3][1][2],image[3][1][3],image[3][1][4],image[3][2][0],image[3][2][1],image[3][2][2],image[3][2][3],image[3][2][4],image[3][3][0],image[3][3][1],image[3][3][2],image[3][3][3],image[3][3][4],image[3][4][0],image[3][4][1],image[3][4][2],image[3][4][3],image[3][4][4],image[3][5][0],image[3][5][1],image[3][5][2],image[3][5][3],image[3][5][4],image[4][1][0],image[4][1][1],image[4][1][2],image[4][1][3],image[4][1][4],image[4][2][0],image[4][2][1],image[4][2][2],image[4][2][3],image[4][2][4],image[4][3][0],image[4][3][1],image[4][3][2],image[4][3][3],image[4][3][4],image[4][4][0],image[4][4][1],image[4][4][2],image[4][4][3],image[4][4][4],image[4][5][0],image[4][5][1],image[4][5][2],image[4][5][3],image[4][5][4],image[5][1][0],image[5][1][1],image[5][1][2],image[5][1][3],image[5][1][4],image[5][2][0],image[5][2][1],image[5][2][2],image[5][2][3],image[5][2][4],image[5][3][0],image[5][3][1],image[5][3][2],image[5][3][3],image[5][3][4],image[5][4][0],image[5][4][1],image[5][4][2],image[5][4][3],image[5][4][4],image[5][5][0],image[5][5][1],image[5][5][2],image[5][5][3],image[5][5][4],image[6][1][0],image[6][1][1],image[6][1][2],image[6][1][3],image[6][1][4],image[6][2][0],image[6][2][1],image[6][2][2],image[6][2][3],image[6][2][4],image[6][3][0],image[6][3][1],image[6][3][2],image[6][3][3],image[6][3][4],image[6][4][0],image[6][4][1],image[6][4][2],image[6][4][3],image[6][4][4],image[6][5][0],image[6][5][1],image[6][5][2],image[6][5][3],image[6][5][4],image[7][1][0],image[7][1][1],image[7][1][2],image[7][1][3],image[7][1][4],image[7][2][0],image[7][2][1],image[7][2][2],image[7][2][3],image[7][2][4],image[7][3][0],image[7][3][1],image[7][3][2],image[7][3][3],image[7][3][4],image[7][4][0],image[7][4][1],image[7][4][2],image[7][4][3],image[7][4][4],image[7][5][0],image[7][5][1],image[7][5][2],image[7][5][3],image[7][5][4],image[8][1][0],image[8][1][1],image[8][1][2],image[8][1][3],image[8][1][4],image[8][2][0],image[8][2][1],image[8][2][2],image[8][2][3],image[8][2][4],image[8][3][0],image[8][3][1],image[8][3][2],image[8][3][3],image[8][3][4],image[8][4][0],image[8][4][1],image[8][4][2],image[8][4][3],image[8][4][4],image[8][5][0],image[8][5][1],image[8][5][2],image[8][5][3],image[8][5][4],image[9][1][0],image[9][1][1],image[9][1][2],image[9][1][3],image[9][1][4],image[9][2][0],image[9][2][1],image[9][2][2],image[9][2][3],image[9][2][4],image[9][3][0],image[9][3][1],image[9][3][2],image[9][3][3],image[9][3][4],image[9][4][0],image[9][4][1],image[9][4][2],image[9][4][3],image[9][4][4],image[9][5][0],image[9][5][1],image[9][5][2],image[9][5][3],image[9][5][4],image[10][1][0],image[10][1][1],image[10][1][2],image[10][1][3],image[10][1][4],image[10][2][0],image[10][2][1],image[10][2][2],image[10][2][3],image[10][2][4],image[10][3][0],image[10][3][1],image[10][3][2],image[10][3][3],image[10][3][4],image[10][4][0],image[10][4][1],image[10][4][2],image[10][4][3],image[10][4][4],image[10][5][0],image[10][5][1],image[10][5][2],image[10][5][3],image[10][5][4],image[11][1][0],image[11][1][1],image[11][1][2],image[11][1][3],image[11][1][4],image[11][2][0],image[11][2][1],image[11][2][2],image[11][2][3],image[11][2][4],image[11][3][0],image[11][3][1],image[11][3][2],image[11][3][3],image[11][3][4],image[11][4][0],image[11][4][1],image[11][4][2],image[11][4][3],image[11][4][4],image[11][5][0],image[11][5][1],image[11][5][2],image[11][5][3],image[11][5][4],image[12][1][0],image[12][1][1],image[12][1][2],image[12][1][3],image[12][1][4],image[12][2][0],image[12][2][1],image[12][2][2],image[12][2][3],image[12][2][4],image[12][3][0],image[12][3][1],image[12][3][2],image[12][3][3],image[12][3][4],image[12][4][0],image[12][4][1],image[12][4][2],image[12][4][3],image[12][4][4],image[12][5][0],image[12][5][1],image[12][5][2],image[12][5][3],image[12][5][4],image[13][1][0],image[13][1][1],image[13][1][2],image[13][1][3],image[13][1][4],image[13][2][0],image[13][2][1],image[13][2][2],image[13][2][3],image[13][2][4],image[13][3][0],image[13][3][1],image[13][3][2],image[13][3][3],image[13][3][4],image[13][4][0],image[13][4][1],image[13][4][2],image[13][4][3],image[13][4][4],image[13][5][0],image[13][5][1],image[13][5][2],image[13][5][3],image[13][5][4],image[14][1][0],image[14][1][1],image[14][1][2],image[14][1][3],image[14][1][4],image[14][2][0],image[14][2][1],image[14][2][2],image[14][2][3],image[14][2][4],image[14][3][0],image[14][3][1],image[14][3][2],image[14][3][3],image[14][3][4],image[14][4][0],image[14][4][1],image[14][4][2],image[14][4][3],image[14][4][4],image[14][5][0],image[14][5][1],image[14][5][2],image[14][5][3],image[14][5][4],image[15][1][0],image[15][1][1],image[15][1][2],image[15][1][3],image[15][1][4],image[15][2][0],image[15][2][1],image[15][2][2],image[15][2][3],image[15][2][4],image[15][3][0],image[15][3][1],image[15][3][2],image[15][3][3],image[15][3][4],image[15][4][0],image[15][4][1],image[15][4][2],image[15][4][3],image[15][4][4],image[15][5][0],image[15][5][1],image[15][5][2],image[15][5][3],image[15][5][4],image[16][1][0],image[16][1][1],image[16][1][2],image[16][1][3],image[16][1][4],image[16][2][0],image[16][2][1],image[16][2][2],image[16][2][3],image[16][2][4],image[16][3][0],image[16][3][1],image[16][3][2],image[16][3][3],image[16][3][4],image[16][4][0],image[16][4][1],image[16][4][2],image[16][4][3],image[16][4][4],image[16][5][0],image[16][5][1],image[16][5][2],image[16][5][3],image[16][5][4],image[17][1][0],image[17][1][1],image[17][1][2],image[17][1][3],image[17][1][4],image[17][2][0],image[17][2][1],image[17][2][2],image[17][2][3],image[17][2][4],image[17][3][0],image[17][3][1],image[17][3][2],image[17][3][3],image[17][3][4],image[17][4][0],image[17][4][1],image[17][4][2],image[17][4][3],image[17][4][4],image[17][5][0],image[17][5][1],image[17][5][2],image[17][5][3],image[17][5][4]};
logic [chan*5*5-1:0] image_slice3;
assign image_slice3 = {image[0][0][1],image[0][0][2],image[0][0][3],image[0][0][4],image[0][0][5],image[0][1][1],image[0][1][2],image[0][1][3],image[0][1][4],image[0][1][5],image[0][2][1],image[0][2][2],image[0][2][3],image[0][2][4],image[0][2][5],image[0][3][1],image[0][3][2],image[0][3][3],image[0][3][4],image[0][3][5],image[0][4][1],image[0][4][2],image[0][4][3],image[0][4][4],image[0][4][5],image[1][0][1],image[1][0][2],image[1][0][3],image[1][0][4],image[1][0][5],image[1][1][1],image[1][1][2],image[1][1][3],image[1][1][4],image[1][1][5],image[1][2][1],image[1][2][2],image[1][2][3],image[1][2][4],image[1][2][5],image[1][3][1],image[1][3][2],image[1][3][3],image[1][3][4],image[1][3][5],image[1][4][1],image[1][4][2],image[1][4][3],image[1][4][4],image[1][4][5],image[2][0][1],image[2][0][2],image[2][0][3],image[2][0][4],image[2][0][5],image[2][1][1],image[2][1][2],image[2][1][3],image[2][1][4],image[2][1][5],image[2][2][1],image[2][2][2],image[2][2][3],image[2][2][4],image[2][2][5],image[2][3][1],image[2][3][2],image[2][3][3],image[2][3][4],image[2][3][5],image[2][4][1],image[2][4][2],image[2][4][3],image[2][4][4],image[2][4][5],image[3][0][1],image[3][0][2],image[3][0][3],image[3][0][4],image[3][0][5],image[3][1][1],image[3][1][2],image[3][1][3],image[3][1][4],image[3][1][5],image[3][2][1],image[3][2][2],image[3][2][3],image[3][2][4],image[3][2][5],image[3][3][1],image[3][3][2],image[3][3][3],image[3][3][4],image[3][3][5],image[3][4][1],image[3][4][2],image[3][4][3],image[3][4][4],image[3][4][5],image[4][0][1],image[4][0][2],image[4][0][3],image[4][0][4],image[4][0][5],image[4][1][1],image[4][1][2],image[4][1][3],image[4][1][4],image[4][1][5],image[4][2][1],image[4][2][2],image[4][2][3],image[4][2][4],image[4][2][5],image[4][3][1],image[4][3][2],image[4][3][3],image[4][3][4],image[4][3][5],image[4][4][1],image[4][4][2],image[4][4][3],image[4][4][4],image[4][4][5],image[5][0][1],image[5][0][2],image[5][0][3],image[5][0][4],image[5][0][5],image[5][1][1],image[5][1][2],image[5][1][3],image[5][1][4],image[5][1][5],image[5][2][1],image[5][2][2],image[5][2][3],image[5][2][4],image[5][2][5],image[5][3][1],image[5][3][2],image[5][3][3],image[5][3][4],image[5][3][5],image[5][4][1],image[5][4][2],image[5][4][3],image[5][4][4],image[5][4][5],image[6][0][1],image[6][0][2],image[6][0][3],image[6][0][4],image[6][0][5],image[6][1][1],image[6][1][2],image[6][1][3],image[6][1][4],image[6][1][5],image[6][2][1],image[6][2][2],image[6][2][3],image[6][2][4],image[6][2][5],image[6][3][1],image[6][3][2],image[6][3][3],image[6][3][4],image[6][3][5],image[6][4][1],image[6][4][2],image[6][4][3],image[6][4][4],image[6][4][5],image[7][0][1],image[7][0][2],image[7][0][3],image[7][0][4],image[7][0][5],image[7][1][1],image[7][1][2],image[7][1][3],image[7][1][4],image[7][1][5],image[7][2][1],image[7][2][2],image[7][2][3],image[7][2][4],image[7][2][5],image[7][3][1],image[7][3][2],image[7][3][3],image[7][3][4],image[7][3][5],image[7][4][1],image[7][4][2],image[7][4][3],image[7][4][4],image[7][4][5],image[8][0][1],image[8][0][2],image[8][0][3],image[8][0][4],image[8][0][5],image[8][1][1],image[8][1][2],image[8][1][3],image[8][1][4],image[8][1][5],image[8][2][1],image[8][2][2],image[8][2][3],image[8][2][4],image[8][2][5],image[8][3][1],image[8][3][2],image[8][3][3],image[8][3][4],image[8][3][5],image[8][4][1],image[8][4][2],image[8][4][3],image[8][4][4],image[8][4][5],image[9][0][1],image[9][0][2],image[9][0][3],image[9][0][4],image[9][0][5],image[9][1][1],image[9][1][2],image[9][1][3],image[9][1][4],image[9][1][5],image[9][2][1],image[9][2][2],image[9][2][3],image[9][2][4],image[9][2][5],image[9][3][1],image[9][3][2],image[9][3][3],image[9][3][4],image[9][3][5],image[9][4][1],image[9][4][2],image[9][4][3],image[9][4][4],image[9][4][5],image[10][0][1],image[10][0][2],image[10][0][3],image[10][0][4],image[10][0][5],image[10][1][1],image[10][1][2],image[10][1][3],image[10][1][4],image[10][1][5],image[10][2][1],image[10][2][2],image[10][2][3],image[10][2][4],image[10][2][5],image[10][3][1],image[10][3][2],image[10][3][3],image[10][3][4],image[10][3][5],image[10][4][1],image[10][4][2],image[10][4][3],image[10][4][4],image[10][4][5],image[11][0][1],image[11][0][2],image[11][0][3],image[11][0][4],image[11][0][5],image[11][1][1],image[11][1][2],image[11][1][3],image[11][1][4],image[11][1][5],image[11][2][1],image[11][2][2],image[11][2][3],image[11][2][4],image[11][2][5],image[11][3][1],image[11][3][2],image[11][3][3],image[11][3][4],image[11][3][5],image[11][4][1],image[11][4][2],image[11][4][3],image[11][4][4],image[11][4][5],image[12][0][1],image[12][0][2],image[12][0][3],image[12][0][4],image[12][0][5],image[12][1][1],image[12][1][2],image[12][1][3],image[12][1][4],image[12][1][5],image[12][2][1],image[12][2][2],image[12][2][3],image[12][2][4],image[12][2][5],image[12][3][1],image[12][3][2],image[12][3][3],image[12][3][4],image[12][3][5],image[12][4][1],image[12][4][2],image[12][4][3],image[12][4][4],image[12][4][5],image[13][0][1],image[13][0][2],image[13][0][3],image[13][0][4],image[13][0][5],image[13][1][1],image[13][1][2],image[13][1][3],image[13][1][4],image[13][1][5],image[13][2][1],image[13][2][2],image[13][2][3],image[13][2][4],image[13][2][5],image[13][3][1],image[13][3][2],image[13][3][3],image[13][3][4],image[13][3][5],image[13][4][1],image[13][4][2],image[13][4][3],image[13][4][4],image[13][4][5],image[14][0][1],image[14][0][2],image[14][0][3],image[14][0][4],image[14][0][5],image[14][1][1],image[14][1][2],image[14][1][3],image[14][1][4],image[14][1][5],image[14][2][1],image[14][2][2],image[14][2][3],image[14][2][4],image[14][2][5],image[14][3][1],image[14][3][2],image[14][3][3],image[14][3][4],image[14][3][5],image[14][4][1],image[14][4][2],image[14][4][3],image[14][4][4],image[14][4][5],image[15][0][1],image[15][0][2],image[15][0][3],image[15][0][4],image[15][0][5],image[15][1][1],image[15][1][2],image[15][1][3],image[15][1][4],image[15][1][5],image[15][2][1],image[15][2][2],image[15][2][3],image[15][2][4],image[15][2][5],image[15][3][1],image[15][3][2],image[15][3][3],image[15][3][4],image[15][3][5],image[15][4][1],image[15][4][2],image[15][4][3],image[15][4][4],image[15][4][5],image[16][0][1],image[16][0][2],image[16][0][3],image[16][0][4],image[16][0][5],image[16][1][1],image[16][1][2],image[16][1][3],image[16][1][4],image[16][1][5],image[16][2][1],image[16][2][2],image[16][2][3],image[16][2][4],image[16][2][5],image[16][3][1],image[16][3][2],image[16][3][3],image[16][3][4],image[16][3][5],image[16][4][1],image[16][4][2],image[16][4][3],image[16][4][4],image[16][4][5],image[17][0][1],image[17][0][2],image[17][0][3],image[17][0][4],image[17][0][5],image[17][1][1],image[17][1][2],image[17][1][3],image[17][1][4],image[17][1][5],image[17][2][1],image[17][2][2],image[17][2][3],image[17][2][4],image[17][2][5],image[17][3][1],image[17][3][2],image[17][3][3],image[17][3][4],image[17][3][5],image[17][4][1],image[17][4][2],image[17][4][3],image[17][4][4],image[17][4][5]};
logic [chan*5*5-1:0] image_slice4;
assign image_slice4 = {image[0][1][1],image[0][1][2],image[0][1][3],image[0][1][4],image[0][1][5],image[0][2][1],image[0][2][2],image[0][2][3],image[0][2][4],image[0][2][5],image[0][3][1],image[0][3][2],image[0][3][3],image[0][3][4],image[0][3][5],image[0][4][1],image[0][4][2],image[0][4][3],image[0][4][4],image[0][4][5],image[0][5][1],image[0][5][2],image[0][5][3],image[0][5][4],image[0][5][5],image[1][1][1],image[1][1][2],image[1][1][3],image[1][1][4],image[1][1][5],image[1][2][1],image[1][2][2],image[1][2][3],image[1][2][4],image[1][2][5],image[1][3][1],image[1][3][2],image[1][3][3],image[1][3][4],image[1][3][5],image[1][4][1],image[1][4][2],image[1][4][3],image[1][4][4],image[1][4][5],image[1][5][1],image[1][5][2],image[1][5][3],image[1][5][4],image[1][5][5],image[2][1][1],image[2][1][2],image[2][1][3],image[2][1][4],image[2][1][5],image[2][2][1],image[2][2][2],image[2][2][3],image[2][2][4],image[2][2][5],image[2][3][1],image[2][3][2],image[2][3][3],image[2][3][4],image[2][3][5],image[2][4][1],image[2][4][2],image[2][4][3],image[2][4][4],image[2][4][5],image[2][5][1],image[2][5][2],image[2][5][3],image[2][5][4],image[2][5][5],image[3][1][1],image[3][1][2],image[3][1][3],image[3][1][4],image[3][1][5],image[3][2][1],image[3][2][2],image[3][2][3],image[3][2][4],image[3][2][5],image[3][3][1],image[3][3][2],image[3][3][3],image[3][3][4],image[3][3][5],image[3][4][1],image[3][4][2],image[3][4][3],image[3][4][4],image[3][4][5],image[3][5][1],image[3][5][2],image[3][5][3],image[3][5][4],image[3][5][5],image[4][1][1],image[4][1][2],image[4][1][3],image[4][1][4],image[4][1][5],image[4][2][1],image[4][2][2],image[4][2][3],image[4][2][4],image[4][2][5],image[4][3][1],image[4][3][2],image[4][3][3],image[4][3][4],image[4][3][5],image[4][4][1],image[4][4][2],image[4][4][3],image[4][4][4],image[4][4][5],image[4][5][1],image[4][5][2],image[4][5][3],image[4][5][4],image[4][5][5],image[5][1][1],image[5][1][2],image[5][1][3],image[5][1][4],image[5][1][5],image[5][2][1],image[5][2][2],image[5][2][3],image[5][2][4],image[5][2][5],image[5][3][1],image[5][3][2],image[5][3][3],image[5][3][4],image[5][3][5],image[5][4][1],image[5][4][2],image[5][4][3],image[5][4][4],image[5][4][5],image[5][5][1],image[5][5][2],image[5][5][3],image[5][5][4],image[5][5][5],image[6][1][1],image[6][1][2],image[6][1][3],image[6][1][4],image[6][1][5],image[6][2][1],image[6][2][2],image[6][2][3],image[6][2][4],image[6][2][5],image[6][3][1],image[6][3][2],image[6][3][3],image[6][3][4],image[6][3][5],image[6][4][1],image[6][4][2],image[6][4][3],image[6][4][4],image[6][4][5],image[6][5][1],image[6][5][2],image[6][5][3],image[6][5][4],image[6][5][5],image[7][1][1],image[7][1][2],image[7][1][3],image[7][1][4],image[7][1][5],image[7][2][1],image[7][2][2],image[7][2][3],image[7][2][4],image[7][2][5],image[7][3][1],image[7][3][2],image[7][3][3],image[7][3][4],image[7][3][5],image[7][4][1],image[7][4][2],image[7][4][3],image[7][4][4],image[7][4][5],image[7][5][1],image[7][5][2],image[7][5][3],image[7][5][4],image[7][5][5],image[8][1][1],image[8][1][2],image[8][1][3],image[8][1][4],image[8][1][5],image[8][2][1],image[8][2][2],image[8][2][3],image[8][2][4],image[8][2][5],image[8][3][1],image[8][3][2],image[8][3][3],image[8][3][4],image[8][3][5],image[8][4][1],image[8][4][2],image[8][4][3],image[8][4][4],image[8][4][5],image[8][5][1],image[8][5][2],image[8][5][3],image[8][5][4],image[8][5][5],image[9][1][1],image[9][1][2],image[9][1][3],image[9][1][4],image[9][1][5],image[9][2][1],image[9][2][2],image[9][2][3],image[9][2][4],image[9][2][5],image[9][3][1],image[9][3][2],image[9][3][3],image[9][3][4],image[9][3][5],image[9][4][1],image[9][4][2],image[9][4][3],image[9][4][4],image[9][4][5],image[9][5][1],image[9][5][2],image[9][5][3],image[9][5][4],image[9][5][5],image[10][1][1],image[10][1][2],image[10][1][3],image[10][1][4],image[10][1][5],image[10][2][1],image[10][2][2],image[10][2][3],image[10][2][4],image[10][2][5],image[10][3][1],image[10][3][2],image[10][3][3],image[10][3][4],image[10][3][5],image[10][4][1],image[10][4][2],image[10][4][3],image[10][4][4],image[10][4][5],image[10][5][1],image[10][5][2],image[10][5][3],image[10][5][4],image[10][5][5],image[11][1][1],image[11][1][2],image[11][1][3],image[11][1][4],image[11][1][5],image[11][2][1],image[11][2][2],image[11][2][3],image[11][2][4],image[11][2][5],image[11][3][1],image[11][3][2],image[11][3][3],image[11][3][4],image[11][3][5],image[11][4][1],image[11][4][2],image[11][4][3],image[11][4][4],image[11][4][5],image[11][5][1],image[11][5][2],image[11][5][3],image[11][5][4],image[11][5][5],image[12][1][1],image[12][1][2],image[12][1][3],image[12][1][4],image[12][1][5],image[12][2][1],image[12][2][2],image[12][2][3],image[12][2][4],image[12][2][5],image[12][3][1],image[12][3][2],image[12][3][3],image[12][3][4],image[12][3][5],image[12][4][1],image[12][4][2],image[12][4][3],image[12][4][4],image[12][4][5],image[12][5][1],image[12][5][2],image[12][5][3],image[12][5][4],image[12][5][5],image[13][1][1],image[13][1][2],image[13][1][3],image[13][1][4],image[13][1][5],image[13][2][1],image[13][2][2],image[13][2][3],image[13][2][4],image[13][2][5],image[13][3][1],image[13][3][2],image[13][3][3],image[13][3][4],image[13][3][5],image[13][4][1],image[13][4][2],image[13][4][3],image[13][4][4],image[13][4][5],image[13][5][1],image[13][5][2],image[13][5][3],image[13][5][4],image[13][5][5],image[14][1][1],image[14][1][2],image[14][1][3],image[14][1][4],image[14][1][5],image[14][2][1],image[14][2][2],image[14][2][3],image[14][2][4],image[14][2][5],image[14][3][1],image[14][3][2],image[14][3][3],image[14][3][4],image[14][3][5],image[14][4][1],image[14][4][2],image[14][4][3],image[14][4][4],image[14][4][5],image[14][5][1],image[14][5][2],image[14][5][3],image[14][5][4],image[14][5][5],image[15][1][1],image[15][1][2],image[15][1][3],image[15][1][4],image[15][1][5],image[15][2][1],image[15][2][2],image[15][2][3],image[15][2][4],image[15][2][5],image[15][3][1],image[15][3][2],image[15][3][3],image[15][3][4],image[15][3][5],image[15][4][1],image[15][4][2],image[15][4][3],image[15][4][4],image[15][4][5],image[15][5][1],image[15][5][2],image[15][5][3],image[15][5][4],image[15][5][5],image[16][1][1],image[16][1][2],image[16][1][3],image[16][1][4],image[16][1][5],image[16][2][1],image[16][2][2],image[16][2][3],image[16][2][4],image[16][2][5],image[16][3][1],image[16][3][2],image[16][3][3],image[16][3][4],image[16][3][5],image[16][4][1],image[16][4][2],image[16][4][3],image[16][4][4],image[16][4][5],image[16][5][1],image[16][5][2],image[16][5][3],image[16][5][4],image[16][5][5],image[17][1][1],image[17][1][2],image[17][1][3],image[17][1][4],image[17][1][5],image[17][2][1],image[17][2][2],image[17][2][3],image[17][2][4],image[17][2][5],image[17][3][1],image[17][3][2],image[17][3][3],image[17][3][4],image[17][3][5],image[17][4][1],image[17][4][2],image[17][4][3],image[17][4][4],image[17][4][5],image[17][5][1],image[17][5][2],image[17][5][3],image[17][5][4],image[17][5][5]};


logic [0:chan*5*5-1] kernel_slice;
assign kernel_slice = {kernels[0][0][0],kernels[0][0][1],kernels[0][0][2],kernels[0][0][3],kernels[0][0][4],kernels[0][1][0],kernels[0][1][1],kernels[0][1][2],kernels[0][1][3],kernels[0][1][4],kernels[0][2][0],kernels[0][2][1],kernels[0][2][2],kernels[0][2][3],kernels[0][2][4],kernels[0][3][0],kernels[0][3][1],kernels[0][3][2],kernels[0][3][3],kernels[0][3][4],kernels[0][4][0],kernels[0][4][1],kernels[0][4][2],kernels[0][4][3],kernels[0][4][4],kernels[1][0][0],kernels[1][0][1],kernels[1][0][2],kernels[1][0][3],kernels[1][0][4],kernels[1][1][0],kernels[1][1][1],kernels[1][1][2],kernels[1][1][3],kernels[1][1][4],kernels[1][2][0],kernels[1][2][1],kernels[1][2][2],kernels[1][2][3],kernels[1][2][4],kernels[1][3][0],kernels[1][3][1],kernels[1][3][2],kernels[1][3][3],kernels[1][3][4],kernels[1][4][0],kernels[1][4][1],kernels[1][4][2],kernels[1][4][3],kernels[1][4][4],kernels[2][0][0],kernels[2][0][1],kernels[2][0][2],kernels[2][0][3],kernels[2][0][4],kernels[2][1][0],kernels[2][1][1],kernels[2][1][2],kernels[2][1][3],kernels[2][1][4],kernels[2][2][0],kernels[2][2][1],kernels[2][2][2],kernels[2][2][3],kernels[2][2][4],kernels[2][3][0],kernels[2][3][1],kernels[2][3][2],kernels[2][3][3],kernels[2][3][4],kernels[2][4][0],kernels[2][4][1],kernels[2][4][2],kernels[2][4][3],kernels[2][4][4],kernels[3][0][0],kernels[3][0][1],kernels[3][0][2],kernels[3][0][3],kernels[3][0][4],kernels[3][1][0],kernels[3][1][1],kernels[3][1][2],kernels[3][1][3],kernels[3][1][4],kernels[3][2][0],kernels[3][2][1],kernels[3][2][2],kernels[3][2][3],kernels[3][2][4],kernels[3][3][0],kernels[3][3][1],kernels[3][3][2],kernels[3][3][3],kernels[3][3][4],kernels[3][4][0],kernels[3][4][1],kernels[3][4][2],kernels[3][4][3],kernels[3][4][4],kernels[4][0][0],kernels[4][0][1],kernels[4][0][2],kernels[4][0][3],kernels[4][0][4],kernels[4][1][0],kernels[4][1][1],kernels[4][1][2],kernels[4][1][3],kernels[4][1][4],kernels[4][2][0],kernels[4][2][1],kernels[4][2][2],kernels[4][2][3],kernels[4][2][4],kernels[4][3][0],kernels[4][3][1],kernels[4][3][2],kernels[4][3][3],kernels[4][3][4],kernels[4][4][0],kernels[4][4][1],kernels[4][4][2],kernels[4][4][3],kernels[4][4][4],kernels[5][0][0],kernels[5][0][1],kernels[5][0][2],kernels[5][0][3],kernels[5][0][4],kernels[5][1][0],kernels[5][1][1],kernels[5][1][2],kernels[5][1][3],kernels[5][1][4],kernels[5][2][0],kernels[5][2][1],kernels[5][2][2],kernels[5][2][3],kernels[5][2][4],kernels[5][3][0],kernels[5][3][1],kernels[5][3][2],kernels[5][3][3],kernels[5][3][4],kernels[5][4][0],kernels[5][4][1],kernels[5][4][2],kernels[5][4][3],kernels[5][4][4],kernels[6][0][0],kernels[6][0][1],kernels[6][0][2],kernels[6][0][3],kernels[6][0][4],kernels[6][1][0],kernels[6][1][1],kernels[6][1][2],kernels[6][1][3],kernels[6][1][4],kernels[6][2][0],kernels[6][2][1],kernels[6][2][2],kernels[6][2][3],kernels[6][2][4],kernels[6][3][0],kernels[6][3][1],kernels[6][3][2],kernels[6][3][3],kernels[6][3][4],kernels[6][4][0],kernels[6][4][1],kernels[6][4][2],kernels[6][4][3],kernels[6][4][4],kernels[7][0][0],kernels[7][0][1],kernels[7][0][2],kernels[7][0][3],kernels[7][0][4],kernels[7][1][0],kernels[7][1][1],kernels[7][1][2],kernels[7][1][3],kernels[7][1][4],kernels[7][2][0],kernels[7][2][1],kernels[7][2][2],kernels[7][2][3],kernels[7][2][4],kernels[7][3][0],kernels[7][3][1],kernels[7][3][2],kernels[7][3][3],kernels[7][3][4],kernels[7][4][0],kernels[7][4][1],kernels[7][4][2],kernels[7][4][3],kernels[7][4][4],kernels[8][0][0],kernels[8][0][1],kernels[8][0][2],kernels[8][0][3],kernels[8][0][4],kernels[8][1][0],kernels[8][1][1],kernels[8][1][2],kernels[8][1][3],kernels[8][1][4],kernels[8][2][0],kernels[8][2][1],kernels[8][2][2],kernels[8][2][3],kernels[8][2][4],kernels[8][3][0],kernels[8][3][1],kernels[8][3][2],kernels[8][3][3],kernels[8][3][4],kernels[8][4][0],kernels[8][4][1],kernels[8][4][2],kernels[8][4][3],kernels[8][4][4],kernels[9][0][0],kernels[9][0][1],kernels[9][0][2],kernels[9][0][3],kernels[9][0][4],kernels[9][1][0],kernels[9][1][1],kernels[9][1][2],kernels[9][1][3],kernels[9][1][4],kernels[9][2][0],kernels[9][2][1],kernels[9][2][2],kernels[9][2][3],kernels[9][2][4],kernels[9][3][0],kernels[9][3][1],kernels[9][3][2],kernels[9][3][3],kernels[9][3][4],kernels[9][4][0],kernels[9][4][1],kernels[9][4][2],kernels[9][4][3],kernels[9][4][4],kernels[10][0][0],kernels[10][0][1],kernels[10][0][2],kernels[10][0][3],kernels[10][0][4],kernels[10][1][0],kernels[10][1][1],kernels[10][1][2],kernels[10][1][3],kernels[10][1][4],kernels[10][2][0],kernels[10][2][1],kernels[10][2][2],kernels[10][2][3],kernels[10][2][4],kernels[10][3][0],kernels[10][3][1],kernels[10][3][2],kernels[10][3][3],kernels[10][3][4],kernels[10][4][0],kernels[10][4][1],kernels[10][4][2],kernels[10][4][3],kernels[10][4][4],kernels[11][0][0],kernels[11][0][1],kernels[11][0][2],kernels[11][0][3],kernels[11][0][4],kernels[11][1][0],kernels[11][1][1],kernels[11][1][2],kernels[11][1][3],kernels[11][1][4],kernels[11][2][0],kernels[11][2][1],kernels[11][2][2],kernels[11][2][3],kernels[11][2][4],kernels[11][3][0],kernels[11][3][1],kernels[11][3][2],kernels[11][3][3],kernels[11][3][4],kernels[11][4][0],kernels[11][4][1],kernels[11][4][2],kernels[11][4][3],kernels[11][4][4],kernels[12][0][0],kernels[12][0][1],kernels[12][0][2],kernels[12][0][3],kernels[12][0][4],kernels[12][1][0],kernels[12][1][1],kernels[12][1][2],kernels[12][1][3],kernels[12][1][4],kernels[12][2][0],kernels[12][2][1],kernels[12][2][2],kernels[12][2][3],kernels[12][2][4],kernels[12][3][0],kernels[12][3][1],kernels[12][3][2],kernels[12][3][3],kernels[12][3][4],kernels[12][4][0],kernels[12][4][1],kernels[12][4][2],kernels[12][4][3],kernels[12][4][4],kernels[13][0][0],kernels[13][0][1],kernels[13][0][2],kernels[13][0][3],kernels[13][0][4],kernels[13][1][0],kernels[13][1][1],kernels[13][1][2],kernels[13][1][3],kernels[13][1][4],kernels[13][2][0],kernels[13][2][1],kernels[13][2][2],kernels[13][2][3],kernels[13][2][4],kernels[13][3][0],kernels[13][3][1],kernels[13][3][2],kernels[13][3][3],kernels[13][3][4],kernels[13][4][0],kernels[13][4][1],kernels[13][4][2],kernels[13][4][3],kernels[13][4][4],kernels[14][0][0],kernels[14][0][1],kernels[14][0][2],kernels[14][0][3],kernels[14][0][4],kernels[14][1][0],kernels[14][1][1],kernels[14][1][2],kernels[14][1][3],kernels[14][1][4],kernels[14][2][0],kernels[14][2][1],kernels[14][2][2],kernels[14][2][3],kernels[14][2][4],kernels[14][3][0],kernels[14][3][1],kernels[14][3][2],kernels[14][3][3],kernels[14][3][4],kernels[14][4][0],kernels[14][4][1],kernels[14][4][2],kernels[14][4][3],kernels[14][4][4],kernels[15][0][0],kernels[15][0][1],kernels[15][0][2],kernels[15][0][3],kernels[15][0][4],kernels[15][1][0],kernels[15][1][1],kernels[15][1][2],kernels[15][1][3],kernels[15][1][4],kernels[15][2][0],kernels[15][2][1],kernels[15][2][2],kernels[15][2][3],kernels[15][2][4],kernels[15][3][0],kernels[15][3][1],kernels[15][3][2],kernels[15][3][3],kernels[15][3][4],kernels[15][4][0],kernels[15][4][1],kernels[15][4][2],kernels[15][4][3],kernels[15][4][4],kernels[16][0][0],kernels[16][0][1],kernels[16][0][2],kernels[16][0][3],kernels[16][0][4],kernels[16][1][0],kernels[16][1][1],kernels[16][1][2],kernels[16][1][3],kernels[16][1][4],kernels[16][2][0],kernels[16][2][1],kernels[16][2][2],kernels[16][2][3],kernels[16][2][4],kernels[16][3][0],kernels[16][3][1],kernels[16][3][2],kernels[16][3][3],kernels[16][3][4],kernels[16][4][0],kernels[16][4][1],kernels[16][4][2],kernels[16][4][3],kernels[16][4][4],kernels[17][0][0],kernels[17][0][1],kernels[17][0][2],kernels[17][0][3],kernels[17][0][4],kernels[17][1][0],kernels[17][1][1],kernels[17][1][2],kernels[17][1][3],kernels[17][1][4],kernels[17][2][0],kernels[17][2][1],kernels[17][2][2],kernels[17][2][3],kernels[17][2][4],kernels[17][3][0],kernels[17][3][1],kernels[17][3][2],kernels[17][3][3],kernels[17][3][4],kernels[17][4][0],kernels[17][4][1],kernels[17][4][2],kernels[17][4][3],kernels[17][4][4]};

logic [0:chan*5*5-1] xnor1, xnor2, xnor3, xnor4;
assign xnor1 = image_slice1 ~^ kernel_slice;
assign xnor2 = image_slice2 ~^ kernel_slice;
assign xnor3 = image_slice3 ~^ kernel_slice;
assign xnor4 = image_slice4 ~^ kernel_slice;

logic [bW-1:0] sum1;
logic [bW-1:0] sum2;
logic [bW-1:0] sum3;
logic [bW-1:0] sum4;

popadd450 p1 (.bits(xnor1), .cnt(sum1));
popadd450 p2 (.bits(xnor2), .cnt(sum2));
popadd450 p3 (.bits(xnor3), .cnt(sum3));
popadd450 p4 (.bits(xnor4), .cnt(sum4));

logic bin1, bin2, bin3, bin4;

assign bin1 = sum1 > offset;
assign bin2 = sum2 > offset;
assign bin3 = sum3 > offset;
assign bin4 = sum4 > offset;

assign pixel = bin1 | bin2 | bin3 | bin4;


endmodule
