module convchan1 
    #( parameter bW = 8 )
    ( 
    input  logic [0:28*28-1]    i_image    ,
    input  logic [0:5*5-1]      i_kernel   ,
    output logic [0:24*24*bW-1] o_out_fmap
    );

logic          image    [0:27][0:27];
logic          kernel   [0: 4][0: 4];
logic [bW-1:0] out_fmap [0:23][0:23];

genvar i,j,k;
for (i=0; i<28; i=i+1) begin
    for (j=0; j<28; j=j+1) begin
        assign image[i][j] = i_image[ 28*i + j ];
    end
end

for (i=0; i<5; i=i+1) begin
    for (j=0; j<5; j=j+1) begin
        assign kernel[i][j] = i_kernel[ 5*i + j ];
    end
end

for (i=0; i<24; i=i+1) begin
    for (j=0; j<24; j=j+1) begin
        for (k=0; k<bW; k=k+1) begin
            assign o_out_fmap[ 24*bW*i + bW*j + k ] = out_fmap[i][j][k];
        end
    end
end

assign out_fmap[0][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][0])} + {7'd0,(kernel[0][1] ~^ image[0][1])} + {7'd0,(kernel[0][2] ~^ image[0][2])} + {7'd0,(kernel[0][3] ~^ image[0][3])} + {7'd0,(kernel[0][4] ~^ image[0][4])} + {7'd0,(kernel[1][0] ~^ image[1][0])} + {7'd0,(kernel[1][1] ~^ image[1][1])} + {7'd0,(kernel[1][2] ~^ image[1][2])} + {7'd0,(kernel[1][3] ~^ image[1][3])} + {7'd0,(kernel[1][4] ~^ image[1][4])} + {7'd0,(kernel[2][0] ~^ image[2][0])} + {7'd0,(kernel[2][1] ~^ image[2][1])} + {7'd0,(kernel[2][2] ~^ image[2][2])} + {7'd0,(kernel[2][3] ~^ image[2][3])} + {7'd0,(kernel[2][4] ~^ image[2][4])} + {7'd0,(kernel[3][0] ~^ image[3][0])} + {7'd0,(kernel[3][1] ~^ image[3][1])} + {7'd0,(kernel[3][2] ~^ image[3][2])} + {7'd0,(kernel[3][3] ~^ image[3][3])} + {7'd0,(kernel[3][4] ~^ image[3][4])} + {7'd0,(kernel[4][0] ~^ image[4][0])} + {7'd0,(kernel[4][1] ~^ image[4][1])} + {7'd0,(kernel[4][2] ~^ image[4][2])} + {7'd0,(kernel[4][3] ~^ image[4][3])} + {7'd0,(kernel[4][4] ~^ image[4][4])};
assign out_fmap[0][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][1])} + {7'd0,(kernel[0][1] ~^ image[0][2])} + {7'd0,(kernel[0][2] ~^ image[0][3])} + {7'd0,(kernel[0][3] ~^ image[0][4])} + {7'd0,(kernel[0][4] ~^ image[0][5])} + {7'd0,(kernel[1][0] ~^ image[1][1])} + {7'd0,(kernel[1][1] ~^ image[1][2])} + {7'd0,(kernel[1][2] ~^ image[1][3])} + {7'd0,(kernel[1][3] ~^ image[1][4])} + {7'd0,(kernel[1][4] ~^ image[1][5])} + {7'd0,(kernel[2][0] ~^ image[2][1])} + {7'd0,(kernel[2][1] ~^ image[2][2])} + {7'd0,(kernel[2][2] ~^ image[2][3])} + {7'd0,(kernel[2][3] ~^ image[2][4])} + {7'd0,(kernel[2][4] ~^ image[2][5])} + {7'd0,(kernel[3][0] ~^ image[3][1])} + {7'd0,(kernel[3][1] ~^ image[3][2])} + {7'd0,(kernel[3][2] ~^ image[3][3])} + {7'd0,(kernel[3][3] ~^ image[3][4])} + {7'd0,(kernel[3][4] ~^ image[3][5])} + {7'd0,(kernel[4][0] ~^ image[4][1])} + {7'd0,(kernel[4][1] ~^ image[4][2])} + {7'd0,(kernel[4][2] ~^ image[4][3])} + {7'd0,(kernel[4][3] ~^ image[4][4])} + {7'd0,(kernel[4][4] ~^ image[4][5])};
assign out_fmap[0][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][2])} + {7'd0,(kernel[0][1] ~^ image[0][3])} + {7'd0,(kernel[0][2] ~^ image[0][4])} + {7'd0,(kernel[0][3] ~^ image[0][5])} + {7'd0,(kernel[0][4] ~^ image[0][6])} + {7'd0,(kernel[1][0] ~^ image[1][2])} + {7'd0,(kernel[1][1] ~^ image[1][3])} + {7'd0,(kernel[1][2] ~^ image[1][4])} + {7'd0,(kernel[1][3] ~^ image[1][5])} + {7'd0,(kernel[1][4] ~^ image[1][6])} + {7'd0,(kernel[2][0] ~^ image[2][2])} + {7'd0,(kernel[2][1] ~^ image[2][3])} + {7'd0,(kernel[2][2] ~^ image[2][4])} + {7'd0,(kernel[2][3] ~^ image[2][5])} + {7'd0,(kernel[2][4] ~^ image[2][6])} + {7'd0,(kernel[3][0] ~^ image[3][2])} + {7'd0,(kernel[3][1] ~^ image[3][3])} + {7'd0,(kernel[3][2] ~^ image[3][4])} + {7'd0,(kernel[3][3] ~^ image[3][5])} + {7'd0,(kernel[3][4] ~^ image[3][6])} + {7'd0,(kernel[4][0] ~^ image[4][2])} + {7'd0,(kernel[4][1] ~^ image[4][3])} + {7'd0,(kernel[4][2] ~^ image[4][4])} + {7'd0,(kernel[4][3] ~^ image[4][5])} + {7'd0,(kernel[4][4] ~^ image[4][6])};
assign out_fmap[0][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][3])} + {7'd0,(kernel[0][1] ~^ image[0][4])} + {7'd0,(kernel[0][2] ~^ image[0][5])} + {7'd0,(kernel[0][3] ~^ image[0][6])} + {7'd0,(kernel[0][4] ~^ image[0][7])} + {7'd0,(kernel[1][0] ~^ image[1][3])} + {7'd0,(kernel[1][1] ~^ image[1][4])} + {7'd0,(kernel[1][2] ~^ image[1][5])} + {7'd0,(kernel[1][3] ~^ image[1][6])} + {7'd0,(kernel[1][4] ~^ image[1][7])} + {7'd0,(kernel[2][0] ~^ image[2][3])} + {7'd0,(kernel[2][1] ~^ image[2][4])} + {7'd0,(kernel[2][2] ~^ image[2][5])} + {7'd0,(kernel[2][3] ~^ image[2][6])} + {7'd0,(kernel[2][4] ~^ image[2][7])} + {7'd0,(kernel[3][0] ~^ image[3][3])} + {7'd0,(kernel[3][1] ~^ image[3][4])} + {7'd0,(kernel[3][2] ~^ image[3][5])} + {7'd0,(kernel[3][3] ~^ image[3][6])} + {7'd0,(kernel[3][4] ~^ image[3][7])} + {7'd0,(kernel[4][0] ~^ image[4][3])} + {7'd0,(kernel[4][1] ~^ image[4][4])} + {7'd0,(kernel[4][2] ~^ image[4][5])} + {7'd0,(kernel[4][3] ~^ image[4][6])} + {7'd0,(kernel[4][4] ~^ image[4][7])};
assign out_fmap[0][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][4])} + {7'd0,(kernel[0][1] ~^ image[0][5])} + {7'd0,(kernel[0][2] ~^ image[0][6])} + {7'd0,(kernel[0][3] ~^ image[0][7])} + {7'd0,(kernel[0][4] ~^ image[0][8])} + {7'd0,(kernel[1][0] ~^ image[1][4])} + {7'd0,(kernel[1][1] ~^ image[1][5])} + {7'd0,(kernel[1][2] ~^ image[1][6])} + {7'd0,(kernel[1][3] ~^ image[1][7])} + {7'd0,(kernel[1][4] ~^ image[1][8])} + {7'd0,(kernel[2][0] ~^ image[2][4])} + {7'd0,(kernel[2][1] ~^ image[2][5])} + {7'd0,(kernel[2][2] ~^ image[2][6])} + {7'd0,(kernel[2][3] ~^ image[2][7])} + {7'd0,(kernel[2][4] ~^ image[2][8])} + {7'd0,(kernel[3][0] ~^ image[3][4])} + {7'd0,(kernel[3][1] ~^ image[3][5])} + {7'd0,(kernel[3][2] ~^ image[3][6])} + {7'd0,(kernel[3][3] ~^ image[3][7])} + {7'd0,(kernel[3][4] ~^ image[3][8])} + {7'd0,(kernel[4][0] ~^ image[4][4])} + {7'd0,(kernel[4][1] ~^ image[4][5])} + {7'd0,(kernel[4][2] ~^ image[4][6])} + {7'd0,(kernel[4][3] ~^ image[4][7])} + {7'd0,(kernel[4][4] ~^ image[4][8])};
assign out_fmap[0][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][5])} + {7'd0,(kernel[0][1] ~^ image[0][6])} + {7'd0,(kernel[0][2] ~^ image[0][7])} + {7'd0,(kernel[0][3] ~^ image[0][8])} + {7'd0,(kernel[0][4] ~^ image[0][9])} + {7'd0,(kernel[1][0] ~^ image[1][5])} + {7'd0,(kernel[1][1] ~^ image[1][6])} + {7'd0,(kernel[1][2] ~^ image[1][7])} + {7'd0,(kernel[1][3] ~^ image[1][8])} + {7'd0,(kernel[1][4] ~^ image[1][9])} + {7'd0,(kernel[2][0] ~^ image[2][5])} + {7'd0,(kernel[2][1] ~^ image[2][6])} + {7'd0,(kernel[2][2] ~^ image[2][7])} + {7'd0,(kernel[2][3] ~^ image[2][8])} + {7'd0,(kernel[2][4] ~^ image[2][9])} + {7'd0,(kernel[3][0] ~^ image[3][5])} + {7'd0,(kernel[3][1] ~^ image[3][6])} + {7'd0,(kernel[3][2] ~^ image[3][7])} + {7'd0,(kernel[3][3] ~^ image[3][8])} + {7'd0,(kernel[3][4] ~^ image[3][9])} + {7'd0,(kernel[4][0] ~^ image[4][5])} + {7'd0,(kernel[4][1] ~^ image[4][6])} + {7'd0,(kernel[4][2] ~^ image[4][7])} + {7'd0,(kernel[4][3] ~^ image[4][8])} + {7'd0,(kernel[4][4] ~^ image[4][9])};
assign out_fmap[0][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][6])} + {7'd0,(kernel[0][1] ~^ image[0][7])} + {7'd0,(kernel[0][2] ~^ image[0][8])} + {7'd0,(kernel[0][3] ~^ image[0][9])} + {7'd0,(kernel[0][4] ~^ image[0][10])} + {7'd0,(kernel[1][0] ~^ image[1][6])} + {7'd0,(kernel[1][1] ~^ image[1][7])} + {7'd0,(kernel[1][2] ~^ image[1][8])} + {7'd0,(kernel[1][3] ~^ image[1][9])} + {7'd0,(kernel[1][4] ~^ image[1][10])} + {7'd0,(kernel[2][0] ~^ image[2][6])} + {7'd0,(kernel[2][1] ~^ image[2][7])} + {7'd0,(kernel[2][2] ~^ image[2][8])} + {7'd0,(kernel[2][3] ~^ image[2][9])} + {7'd0,(kernel[2][4] ~^ image[2][10])} + {7'd0,(kernel[3][0] ~^ image[3][6])} + {7'd0,(kernel[3][1] ~^ image[3][7])} + {7'd0,(kernel[3][2] ~^ image[3][8])} + {7'd0,(kernel[3][3] ~^ image[3][9])} + {7'd0,(kernel[3][4] ~^ image[3][10])} + {7'd0,(kernel[4][0] ~^ image[4][6])} + {7'd0,(kernel[4][1] ~^ image[4][7])} + {7'd0,(kernel[4][2] ~^ image[4][8])} + {7'd0,(kernel[4][3] ~^ image[4][9])} + {7'd0,(kernel[4][4] ~^ image[4][10])};
assign out_fmap[0][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][7])} + {7'd0,(kernel[0][1] ~^ image[0][8])} + {7'd0,(kernel[0][2] ~^ image[0][9])} + {7'd0,(kernel[0][3] ~^ image[0][10])} + {7'd0,(kernel[0][4] ~^ image[0][11])} + {7'd0,(kernel[1][0] ~^ image[1][7])} + {7'd0,(kernel[1][1] ~^ image[1][8])} + {7'd0,(kernel[1][2] ~^ image[1][9])} + {7'd0,(kernel[1][3] ~^ image[1][10])} + {7'd0,(kernel[1][4] ~^ image[1][11])} + {7'd0,(kernel[2][0] ~^ image[2][7])} + {7'd0,(kernel[2][1] ~^ image[2][8])} + {7'd0,(kernel[2][2] ~^ image[2][9])} + {7'd0,(kernel[2][3] ~^ image[2][10])} + {7'd0,(kernel[2][4] ~^ image[2][11])} + {7'd0,(kernel[3][0] ~^ image[3][7])} + {7'd0,(kernel[3][1] ~^ image[3][8])} + {7'd0,(kernel[3][2] ~^ image[3][9])} + {7'd0,(kernel[3][3] ~^ image[3][10])} + {7'd0,(kernel[3][4] ~^ image[3][11])} + {7'd0,(kernel[4][0] ~^ image[4][7])} + {7'd0,(kernel[4][1] ~^ image[4][8])} + {7'd0,(kernel[4][2] ~^ image[4][9])} + {7'd0,(kernel[4][3] ~^ image[4][10])} + {7'd0,(kernel[4][4] ~^ image[4][11])};
assign out_fmap[0][8][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][8])} + {7'd0,(kernel[0][1] ~^ image[0][9])} + {7'd0,(kernel[0][2] ~^ image[0][10])} + {7'd0,(kernel[0][3] ~^ image[0][11])} + {7'd0,(kernel[0][4] ~^ image[0][12])} + {7'd0,(kernel[1][0] ~^ image[1][8])} + {7'd0,(kernel[1][1] ~^ image[1][9])} + {7'd0,(kernel[1][2] ~^ image[1][10])} + {7'd0,(kernel[1][3] ~^ image[1][11])} + {7'd0,(kernel[1][4] ~^ image[1][12])} + {7'd0,(kernel[2][0] ~^ image[2][8])} + {7'd0,(kernel[2][1] ~^ image[2][9])} + {7'd0,(kernel[2][2] ~^ image[2][10])} + {7'd0,(kernel[2][3] ~^ image[2][11])} + {7'd0,(kernel[2][4] ~^ image[2][12])} + {7'd0,(kernel[3][0] ~^ image[3][8])} + {7'd0,(kernel[3][1] ~^ image[3][9])} + {7'd0,(kernel[3][2] ~^ image[3][10])} + {7'd0,(kernel[3][3] ~^ image[3][11])} + {7'd0,(kernel[3][4] ~^ image[3][12])} + {7'd0,(kernel[4][0] ~^ image[4][8])} + {7'd0,(kernel[4][1] ~^ image[4][9])} + {7'd0,(kernel[4][2] ~^ image[4][10])} + {7'd0,(kernel[4][3] ~^ image[4][11])} + {7'd0,(kernel[4][4] ~^ image[4][12])};
assign out_fmap[0][9][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][9])} + {7'd0,(kernel[0][1] ~^ image[0][10])} + {7'd0,(kernel[0][2] ~^ image[0][11])} + {7'd0,(kernel[0][3] ~^ image[0][12])} + {7'd0,(kernel[0][4] ~^ image[0][13])} + {7'd0,(kernel[1][0] ~^ image[1][9])} + {7'd0,(kernel[1][1] ~^ image[1][10])} + {7'd0,(kernel[1][2] ~^ image[1][11])} + {7'd0,(kernel[1][3] ~^ image[1][12])} + {7'd0,(kernel[1][4] ~^ image[1][13])} + {7'd0,(kernel[2][0] ~^ image[2][9])} + {7'd0,(kernel[2][1] ~^ image[2][10])} + {7'd0,(kernel[2][2] ~^ image[2][11])} + {7'd0,(kernel[2][3] ~^ image[2][12])} + {7'd0,(kernel[2][4] ~^ image[2][13])} + {7'd0,(kernel[3][0] ~^ image[3][9])} + {7'd0,(kernel[3][1] ~^ image[3][10])} + {7'd0,(kernel[3][2] ~^ image[3][11])} + {7'd0,(kernel[3][3] ~^ image[3][12])} + {7'd0,(kernel[3][4] ~^ image[3][13])} + {7'd0,(kernel[4][0] ~^ image[4][9])} + {7'd0,(kernel[4][1] ~^ image[4][10])} + {7'd0,(kernel[4][2] ~^ image[4][11])} + {7'd0,(kernel[4][3] ~^ image[4][12])} + {7'd0,(kernel[4][4] ~^ image[4][13])};
assign out_fmap[0][10][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][10])} + {7'd0,(kernel[0][1] ~^ image[0][11])} + {7'd0,(kernel[0][2] ~^ image[0][12])} + {7'd0,(kernel[0][3] ~^ image[0][13])} + {7'd0,(kernel[0][4] ~^ image[0][14])} + {7'd0,(kernel[1][0] ~^ image[1][10])} + {7'd0,(kernel[1][1] ~^ image[1][11])} + {7'd0,(kernel[1][2] ~^ image[1][12])} + {7'd0,(kernel[1][3] ~^ image[1][13])} + {7'd0,(kernel[1][4] ~^ image[1][14])} + {7'd0,(kernel[2][0] ~^ image[2][10])} + {7'd0,(kernel[2][1] ~^ image[2][11])} + {7'd0,(kernel[2][2] ~^ image[2][12])} + {7'd0,(kernel[2][3] ~^ image[2][13])} + {7'd0,(kernel[2][4] ~^ image[2][14])} + {7'd0,(kernel[3][0] ~^ image[3][10])} + {7'd0,(kernel[3][1] ~^ image[3][11])} + {7'd0,(kernel[3][2] ~^ image[3][12])} + {7'd0,(kernel[3][3] ~^ image[3][13])} + {7'd0,(kernel[3][4] ~^ image[3][14])} + {7'd0,(kernel[4][0] ~^ image[4][10])} + {7'd0,(kernel[4][1] ~^ image[4][11])} + {7'd0,(kernel[4][2] ~^ image[4][12])} + {7'd0,(kernel[4][3] ~^ image[4][13])} + {7'd0,(kernel[4][4] ~^ image[4][14])};
assign out_fmap[0][11][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][11])} + {7'd0,(kernel[0][1] ~^ image[0][12])} + {7'd0,(kernel[0][2] ~^ image[0][13])} + {7'd0,(kernel[0][3] ~^ image[0][14])} + {7'd0,(kernel[0][4] ~^ image[0][15])} + {7'd0,(kernel[1][0] ~^ image[1][11])} + {7'd0,(kernel[1][1] ~^ image[1][12])} + {7'd0,(kernel[1][2] ~^ image[1][13])} + {7'd0,(kernel[1][3] ~^ image[1][14])} + {7'd0,(kernel[1][4] ~^ image[1][15])} + {7'd0,(kernel[2][0] ~^ image[2][11])} + {7'd0,(kernel[2][1] ~^ image[2][12])} + {7'd0,(kernel[2][2] ~^ image[2][13])} + {7'd0,(kernel[2][3] ~^ image[2][14])} + {7'd0,(kernel[2][4] ~^ image[2][15])} + {7'd0,(kernel[3][0] ~^ image[3][11])} + {7'd0,(kernel[3][1] ~^ image[3][12])} + {7'd0,(kernel[3][2] ~^ image[3][13])} + {7'd0,(kernel[3][3] ~^ image[3][14])} + {7'd0,(kernel[3][4] ~^ image[3][15])} + {7'd0,(kernel[4][0] ~^ image[4][11])} + {7'd0,(kernel[4][1] ~^ image[4][12])} + {7'd0,(kernel[4][2] ~^ image[4][13])} + {7'd0,(kernel[4][3] ~^ image[4][14])} + {7'd0,(kernel[4][4] ~^ image[4][15])};
assign out_fmap[0][12][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][12])} + {7'd0,(kernel[0][1] ~^ image[0][13])} + {7'd0,(kernel[0][2] ~^ image[0][14])} + {7'd0,(kernel[0][3] ~^ image[0][15])} + {7'd0,(kernel[0][4] ~^ image[0][16])} + {7'd0,(kernel[1][0] ~^ image[1][12])} + {7'd0,(kernel[1][1] ~^ image[1][13])} + {7'd0,(kernel[1][2] ~^ image[1][14])} + {7'd0,(kernel[1][3] ~^ image[1][15])} + {7'd0,(kernel[1][4] ~^ image[1][16])} + {7'd0,(kernel[2][0] ~^ image[2][12])} + {7'd0,(kernel[2][1] ~^ image[2][13])} + {7'd0,(kernel[2][2] ~^ image[2][14])} + {7'd0,(kernel[2][3] ~^ image[2][15])} + {7'd0,(kernel[2][4] ~^ image[2][16])} + {7'd0,(kernel[3][0] ~^ image[3][12])} + {7'd0,(kernel[3][1] ~^ image[3][13])} + {7'd0,(kernel[3][2] ~^ image[3][14])} + {7'd0,(kernel[3][3] ~^ image[3][15])} + {7'd0,(kernel[3][4] ~^ image[3][16])} + {7'd0,(kernel[4][0] ~^ image[4][12])} + {7'd0,(kernel[4][1] ~^ image[4][13])} + {7'd0,(kernel[4][2] ~^ image[4][14])} + {7'd0,(kernel[4][3] ~^ image[4][15])} + {7'd0,(kernel[4][4] ~^ image[4][16])};
assign out_fmap[0][13][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][13])} + {7'd0,(kernel[0][1] ~^ image[0][14])} + {7'd0,(kernel[0][2] ~^ image[0][15])} + {7'd0,(kernel[0][3] ~^ image[0][16])} + {7'd0,(kernel[0][4] ~^ image[0][17])} + {7'd0,(kernel[1][0] ~^ image[1][13])} + {7'd0,(kernel[1][1] ~^ image[1][14])} + {7'd0,(kernel[1][2] ~^ image[1][15])} + {7'd0,(kernel[1][3] ~^ image[1][16])} + {7'd0,(kernel[1][4] ~^ image[1][17])} + {7'd0,(kernel[2][0] ~^ image[2][13])} + {7'd0,(kernel[2][1] ~^ image[2][14])} + {7'd0,(kernel[2][2] ~^ image[2][15])} + {7'd0,(kernel[2][3] ~^ image[2][16])} + {7'd0,(kernel[2][4] ~^ image[2][17])} + {7'd0,(kernel[3][0] ~^ image[3][13])} + {7'd0,(kernel[3][1] ~^ image[3][14])} + {7'd0,(kernel[3][2] ~^ image[3][15])} + {7'd0,(kernel[3][3] ~^ image[3][16])} + {7'd0,(kernel[3][4] ~^ image[3][17])} + {7'd0,(kernel[4][0] ~^ image[4][13])} + {7'd0,(kernel[4][1] ~^ image[4][14])} + {7'd0,(kernel[4][2] ~^ image[4][15])} + {7'd0,(kernel[4][3] ~^ image[4][16])} + {7'd0,(kernel[4][4] ~^ image[4][17])};
assign out_fmap[0][14][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][14])} + {7'd0,(kernel[0][1] ~^ image[0][15])} + {7'd0,(kernel[0][2] ~^ image[0][16])} + {7'd0,(kernel[0][3] ~^ image[0][17])} + {7'd0,(kernel[0][4] ~^ image[0][18])} + {7'd0,(kernel[1][0] ~^ image[1][14])} + {7'd0,(kernel[1][1] ~^ image[1][15])} + {7'd0,(kernel[1][2] ~^ image[1][16])} + {7'd0,(kernel[1][3] ~^ image[1][17])} + {7'd0,(kernel[1][4] ~^ image[1][18])} + {7'd0,(kernel[2][0] ~^ image[2][14])} + {7'd0,(kernel[2][1] ~^ image[2][15])} + {7'd0,(kernel[2][2] ~^ image[2][16])} + {7'd0,(kernel[2][3] ~^ image[2][17])} + {7'd0,(kernel[2][4] ~^ image[2][18])} + {7'd0,(kernel[3][0] ~^ image[3][14])} + {7'd0,(kernel[3][1] ~^ image[3][15])} + {7'd0,(kernel[3][2] ~^ image[3][16])} + {7'd0,(kernel[3][3] ~^ image[3][17])} + {7'd0,(kernel[3][4] ~^ image[3][18])} + {7'd0,(kernel[4][0] ~^ image[4][14])} + {7'd0,(kernel[4][1] ~^ image[4][15])} + {7'd0,(kernel[4][2] ~^ image[4][16])} + {7'd0,(kernel[4][3] ~^ image[4][17])} + {7'd0,(kernel[4][4] ~^ image[4][18])};
assign out_fmap[0][15][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][15])} + {7'd0,(kernel[0][1] ~^ image[0][16])} + {7'd0,(kernel[0][2] ~^ image[0][17])} + {7'd0,(kernel[0][3] ~^ image[0][18])} + {7'd0,(kernel[0][4] ~^ image[0][19])} + {7'd0,(kernel[1][0] ~^ image[1][15])} + {7'd0,(kernel[1][1] ~^ image[1][16])} + {7'd0,(kernel[1][2] ~^ image[1][17])} + {7'd0,(kernel[1][3] ~^ image[1][18])} + {7'd0,(kernel[1][4] ~^ image[1][19])} + {7'd0,(kernel[2][0] ~^ image[2][15])} + {7'd0,(kernel[2][1] ~^ image[2][16])} + {7'd0,(kernel[2][2] ~^ image[2][17])} + {7'd0,(kernel[2][3] ~^ image[2][18])} + {7'd0,(kernel[2][4] ~^ image[2][19])} + {7'd0,(kernel[3][0] ~^ image[3][15])} + {7'd0,(kernel[3][1] ~^ image[3][16])} + {7'd0,(kernel[3][2] ~^ image[3][17])} + {7'd0,(kernel[3][3] ~^ image[3][18])} + {7'd0,(kernel[3][4] ~^ image[3][19])} + {7'd0,(kernel[4][0] ~^ image[4][15])} + {7'd0,(kernel[4][1] ~^ image[4][16])} + {7'd0,(kernel[4][2] ~^ image[4][17])} + {7'd0,(kernel[4][3] ~^ image[4][18])} + {7'd0,(kernel[4][4] ~^ image[4][19])};
assign out_fmap[0][16][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][16])} + {7'd0,(kernel[0][1] ~^ image[0][17])} + {7'd0,(kernel[0][2] ~^ image[0][18])} + {7'd0,(kernel[0][3] ~^ image[0][19])} + {7'd0,(kernel[0][4] ~^ image[0][20])} + {7'd0,(kernel[1][0] ~^ image[1][16])} + {7'd0,(kernel[1][1] ~^ image[1][17])} + {7'd0,(kernel[1][2] ~^ image[1][18])} + {7'd0,(kernel[1][3] ~^ image[1][19])} + {7'd0,(kernel[1][4] ~^ image[1][20])} + {7'd0,(kernel[2][0] ~^ image[2][16])} + {7'd0,(kernel[2][1] ~^ image[2][17])} + {7'd0,(kernel[2][2] ~^ image[2][18])} + {7'd0,(kernel[2][3] ~^ image[2][19])} + {7'd0,(kernel[2][4] ~^ image[2][20])} + {7'd0,(kernel[3][0] ~^ image[3][16])} + {7'd0,(kernel[3][1] ~^ image[3][17])} + {7'd0,(kernel[3][2] ~^ image[3][18])} + {7'd0,(kernel[3][3] ~^ image[3][19])} + {7'd0,(kernel[3][4] ~^ image[3][20])} + {7'd0,(kernel[4][0] ~^ image[4][16])} + {7'd0,(kernel[4][1] ~^ image[4][17])} + {7'd0,(kernel[4][2] ~^ image[4][18])} + {7'd0,(kernel[4][3] ~^ image[4][19])} + {7'd0,(kernel[4][4] ~^ image[4][20])};
assign out_fmap[0][17][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][17])} + {7'd0,(kernel[0][1] ~^ image[0][18])} + {7'd0,(kernel[0][2] ~^ image[0][19])} + {7'd0,(kernel[0][3] ~^ image[0][20])} + {7'd0,(kernel[0][4] ~^ image[0][21])} + {7'd0,(kernel[1][0] ~^ image[1][17])} + {7'd0,(kernel[1][1] ~^ image[1][18])} + {7'd0,(kernel[1][2] ~^ image[1][19])} + {7'd0,(kernel[1][3] ~^ image[1][20])} + {7'd0,(kernel[1][4] ~^ image[1][21])} + {7'd0,(kernel[2][0] ~^ image[2][17])} + {7'd0,(kernel[2][1] ~^ image[2][18])} + {7'd0,(kernel[2][2] ~^ image[2][19])} + {7'd0,(kernel[2][3] ~^ image[2][20])} + {7'd0,(kernel[2][4] ~^ image[2][21])} + {7'd0,(kernel[3][0] ~^ image[3][17])} + {7'd0,(kernel[3][1] ~^ image[3][18])} + {7'd0,(kernel[3][2] ~^ image[3][19])} + {7'd0,(kernel[3][3] ~^ image[3][20])} + {7'd0,(kernel[3][4] ~^ image[3][21])} + {7'd0,(kernel[4][0] ~^ image[4][17])} + {7'd0,(kernel[4][1] ~^ image[4][18])} + {7'd0,(kernel[4][2] ~^ image[4][19])} + {7'd0,(kernel[4][3] ~^ image[4][20])} + {7'd0,(kernel[4][4] ~^ image[4][21])};
assign out_fmap[0][18][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][18])} + {7'd0,(kernel[0][1] ~^ image[0][19])} + {7'd0,(kernel[0][2] ~^ image[0][20])} + {7'd0,(kernel[0][3] ~^ image[0][21])} + {7'd0,(kernel[0][4] ~^ image[0][22])} + {7'd0,(kernel[1][0] ~^ image[1][18])} + {7'd0,(kernel[1][1] ~^ image[1][19])} + {7'd0,(kernel[1][2] ~^ image[1][20])} + {7'd0,(kernel[1][3] ~^ image[1][21])} + {7'd0,(kernel[1][4] ~^ image[1][22])} + {7'd0,(kernel[2][0] ~^ image[2][18])} + {7'd0,(kernel[2][1] ~^ image[2][19])} + {7'd0,(kernel[2][2] ~^ image[2][20])} + {7'd0,(kernel[2][3] ~^ image[2][21])} + {7'd0,(kernel[2][4] ~^ image[2][22])} + {7'd0,(kernel[3][0] ~^ image[3][18])} + {7'd0,(kernel[3][1] ~^ image[3][19])} + {7'd0,(kernel[3][2] ~^ image[3][20])} + {7'd0,(kernel[3][3] ~^ image[3][21])} + {7'd0,(kernel[3][4] ~^ image[3][22])} + {7'd0,(kernel[4][0] ~^ image[4][18])} + {7'd0,(kernel[4][1] ~^ image[4][19])} + {7'd0,(kernel[4][2] ~^ image[4][20])} + {7'd0,(kernel[4][3] ~^ image[4][21])} + {7'd0,(kernel[4][4] ~^ image[4][22])};
assign out_fmap[0][19][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][19])} + {7'd0,(kernel[0][1] ~^ image[0][20])} + {7'd0,(kernel[0][2] ~^ image[0][21])} + {7'd0,(kernel[0][3] ~^ image[0][22])} + {7'd0,(kernel[0][4] ~^ image[0][23])} + {7'd0,(kernel[1][0] ~^ image[1][19])} + {7'd0,(kernel[1][1] ~^ image[1][20])} + {7'd0,(kernel[1][2] ~^ image[1][21])} + {7'd0,(kernel[1][3] ~^ image[1][22])} + {7'd0,(kernel[1][4] ~^ image[1][23])} + {7'd0,(kernel[2][0] ~^ image[2][19])} + {7'd0,(kernel[2][1] ~^ image[2][20])} + {7'd0,(kernel[2][2] ~^ image[2][21])} + {7'd0,(kernel[2][3] ~^ image[2][22])} + {7'd0,(kernel[2][4] ~^ image[2][23])} + {7'd0,(kernel[3][0] ~^ image[3][19])} + {7'd0,(kernel[3][1] ~^ image[3][20])} + {7'd0,(kernel[3][2] ~^ image[3][21])} + {7'd0,(kernel[3][3] ~^ image[3][22])} + {7'd0,(kernel[3][4] ~^ image[3][23])} + {7'd0,(kernel[4][0] ~^ image[4][19])} + {7'd0,(kernel[4][1] ~^ image[4][20])} + {7'd0,(kernel[4][2] ~^ image[4][21])} + {7'd0,(kernel[4][3] ~^ image[4][22])} + {7'd0,(kernel[4][4] ~^ image[4][23])};
assign out_fmap[0][20][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][20])} + {7'd0,(kernel[0][1] ~^ image[0][21])} + {7'd0,(kernel[0][2] ~^ image[0][22])} + {7'd0,(kernel[0][3] ~^ image[0][23])} + {7'd0,(kernel[0][4] ~^ image[0][24])} + {7'd0,(kernel[1][0] ~^ image[1][20])} + {7'd0,(kernel[1][1] ~^ image[1][21])} + {7'd0,(kernel[1][2] ~^ image[1][22])} + {7'd0,(kernel[1][3] ~^ image[1][23])} + {7'd0,(kernel[1][4] ~^ image[1][24])} + {7'd0,(kernel[2][0] ~^ image[2][20])} + {7'd0,(kernel[2][1] ~^ image[2][21])} + {7'd0,(kernel[2][2] ~^ image[2][22])} + {7'd0,(kernel[2][3] ~^ image[2][23])} + {7'd0,(kernel[2][4] ~^ image[2][24])} + {7'd0,(kernel[3][0] ~^ image[3][20])} + {7'd0,(kernel[3][1] ~^ image[3][21])} + {7'd0,(kernel[3][2] ~^ image[3][22])} + {7'd0,(kernel[3][3] ~^ image[3][23])} + {7'd0,(kernel[3][4] ~^ image[3][24])} + {7'd0,(kernel[4][0] ~^ image[4][20])} + {7'd0,(kernel[4][1] ~^ image[4][21])} + {7'd0,(kernel[4][2] ~^ image[4][22])} + {7'd0,(kernel[4][3] ~^ image[4][23])} + {7'd0,(kernel[4][4] ~^ image[4][24])};
assign out_fmap[0][21][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][21])} + {7'd0,(kernel[0][1] ~^ image[0][22])} + {7'd0,(kernel[0][2] ~^ image[0][23])} + {7'd0,(kernel[0][3] ~^ image[0][24])} + {7'd0,(kernel[0][4] ~^ image[0][25])} + {7'd0,(kernel[1][0] ~^ image[1][21])} + {7'd0,(kernel[1][1] ~^ image[1][22])} + {7'd0,(kernel[1][2] ~^ image[1][23])} + {7'd0,(kernel[1][3] ~^ image[1][24])} + {7'd0,(kernel[1][4] ~^ image[1][25])} + {7'd0,(kernel[2][0] ~^ image[2][21])} + {7'd0,(kernel[2][1] ~^ image[2][22])} + {7'd0,(kernel[2][2] ~^ image[2][23])} + {7'd0,(kernel[2][3] ~^ image[2][24])} + {7'd0,(kernel[2][4] ~^ image[2][25])} + {7'd0,(kernel[3][0] ~^ image[3][21])} + {7'd0,(kernel[3][1] ~^ image[3][22])} + {7'd0,(kernel[3][2] ~^ image[3][23])} + {7'd0,(kernel[3][3] ~^ image[3][24])} + {7'd0,(kernel[3][4] ~^ image[3][25])} + {7'd0,(kernel[4][0] ~^ image[4][21])} + {7'd0,(kernel[4][1] ~^ image[4][22])} + {7'd0,(kernel[4][2] ~^ image[4][23])} + {7'd0,(kernel[4][3] ~^ image[4][24])} + {7'd0,(kernel[4][4] ~^ image[4][25])};
assign out_fmap[0][22][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][22])} + {7'd0,(kernel[0][1] ~^ image[0][23])} + {7'd0,(kernel[0][2] ~^ image[0][24])} + {7'd0,(kernel[0][3] ~^ image[0][25])} + {7'd0,(kernel[0][4] ~^ image[0][26])} + {7'd0,(kernel[1][0] ~^ image[1][22])} + {7'd0,(kernel[1][1] ~^ image[1][23])} + {7'd0,(kernel[1][2] ~^ image[1][24])} + {7'd0,(kernel[1][3] ~^ image[1][25])} + {7'd0,(kernel[1][4] ~^ image[1][26])} + {7'd0,(kernel[2][0] ~^ image[2][22])} + {7'd0,(kernel[2][1] ~^ image[2][23])} + {7'd0,(kernel[2][2] ~^ image[2][24])} + {7'd0,(kernel[2][3] ~^ image[2][25])} + {7'd0,(kernel[2][4] ~^ image[2][26])} + {7'd0,(kernel[3][0] ~^ image[3][22])} + {7'd0,(kernel[3][1] ~^ image[3][23])} + {7'd0,(kernel[3][2] ~^ image[3][24])} + {7'd0,(kernel[3][3] ~^ image[3][25])} + {7'd0,(kernel[3][4] ~^ image[3][26])} + {7'd0,(kernel[4][0] ~^ image[4][22])} + {7'd0,(kernel[4][1] ~^ image[4][23])} + {7'd0,(kernel[4][2] ~^ image[4][24])} + {7'd0,(kernel[4][3] ~^ image[4][25])} + {7'd0,(kernel[4][4] ~^ image[4][26])};
assign out_fmap[0][23][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[0][23])} + {7'd0,(kernel[0][1] ~^ image[0][24])} + {7'd0,(kernel[0][2] ~^ image[0][25])} + {7'd0,(kernel[0][3] ~^ image[0][26])} + {7'd0,(kernel[0][4] ~^ image[0][27])} + {7'd0,(kernel[1][0] ~^ image[1][23])} + {7'd0,(kernel[1][1] ~^ image[1][24])} + {7'd0,(kernel[1][2] ~^ image[1][25])} + {7'd0,(kernel[1][3] ~^ image[1][26])} + {7'd0,(kernel[1][4] ~^ image[1][27])} + {7'd0,(kernel[2][0] ~^ image[2][23])} + {7'd0,(kernel[2][1] ~^ image[2][24])} + {7'd0,(kernel[2][2] ~^ image[2][25])} + {7'd0,(kernel[2][3] ~^ image[2][26])} + {7'd0,(kernel[2][4] ~^ image[2][27])} + {7'd0,(kernel[3][0] ~^ image[3][23])} + {7'd0,(kernel[3][1] ~^ image[3][24])} + {7'd0,(kernel[3][2] ~^ image[3][25])} + {7'd0,(kernel[3][3] ~^ image[3][26])} + {7'd0,(kernel[3][4] ~^ image[3][27])} + {7'd0,(kernel[4][0] ~^ image[4][23])} + {7'd0,(kernel[4][1] ~^ image[4][24])} + {7'd0,(kernel[4][2] ~^ image[4][25])} + {7'd0,(kernel[4][3] ~^ image[4][26])} + {7'd0,(kernel[4][4] ~^ image[4][27])};
assign out_fmap[1][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][0])} + {7'd0,(kernel[0][1] ~^ image[1][1])} + {7'd0,(kernel[0][2] ~^ image[1][2])} + {7'd0,(kernel[0][3] ~^ image[1][3])} + {7'd0,(kernel[0][4] ~^ image[1][4])} + {7'd0,(kernel[1][0] ~^ image[2][0])} + {7'd0,(kernel[1][1] ~^ image[2][1])} + {7'd0,(kernel[1][2] ~^ image[2][2])} + {7'd0,(kernel[1][3] ~^ image[2][3])} + {7'd0,(kernel[1][4] ~^ image[2][4])} + {7'd0,(kernel[2][0] ~^ image[3][0])} + {7'd0,(kernel[2][1] ~^ image[3][1])} + {7'd0,(kernel[2][2] ~^ image[3][2])} + {7'd0,(kernel[2][3] ~^ image[3][3])} + {7'd0,(kernel[2][4] ~^ image[3][4])} + {7'd0,(kernel[3][0] ~^ image[4][0])} + {7'd0,(kernel[3][1] ~^ image[4][1])} + {7'd0,(kernel[3][2] ~^ image[4][2])} + {7'd0,(kernel[3][3] ~^ image[4][3])} + {7'd0,(kernel[3][4] ~^ image[4][4])} + {7'd0,(kernel[4][0] ~^ image[5][0])} + {7'd0,(kernel[4][1] ~^ image[5][1])} + {7'd0,(kernel[4][2] ~^ image[5][2])} + {7'd0,(kernel[4][3] ~^ image[5][3])} + {7'd0,(kernel[4][4] ~^ image[5][4])};
assign out_fmap[1][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][1])} + {7'd0,(kernel[0][1] ~^ image[1][2])} + {7'd0,(kernel[0][2] ~^ image[1][3])} + {7'd0,(kernel[0][3] ~^ image[1][4])} + {7'd0,(kernel[0][4] ~^ image[1][5])} + {7'd0,(kernel[1][0] ~^ image[2][1])} + {7'd0,(kernel[1][1] ~^ image[2][2])} + {7'd0,(kernel[1][2] ~^ image[2][3])} + {7'd0,(kernel[1][3] ~^ image[2][4])} + {7'd0,(kernel[1][4] ~^ image[2][5])} + {7'd0,(kernel[2][0] ~^ image[3][1])} + {7'd0,(kernel[2][1] ~^ image[3][2])} + {7'd0,(kernel[2][2] ~^ image[3][3])} + {7'd0,(kernel[2][3] ~^ image[3][4])} + {7'd0,(kernel[2][4] ~^ image[3][5])} + {7'd0,(kernel[3][0] ~^ image[4][1])} + {7'd0,(kernel[3][1] ~^ image[4][2])} + {7'd0,(kernel[3][2] ~^ image[4][3])} + {7'd0,(kernel[3][3] ~^ image[4][4])} + {7'd0,(kernel[3][4] ~^ image[4][5])} + {7'd0,(kernel[4][0] ~^ image[5][1])} + {7'd0,(kernel[4][1] ~^ image[5][2])} + {7'd0,(kernel[4][2] ~^ image[5][3])} + {7'd0,(kernel[4][3] ~^ image[5][4])} + {7'd0,(kernel[4][4] ~^ image[5][5])};
assign out_fmap[1][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][2])} + {7'd0,(kernel[0][1] ~^ image[1][3])} + {7'd0,(kernel[0][2] ~^ image[1][4])} + {7'd0,(kernel[0][3] ~^ image[1][5])} + {7'd0,(kernel[0][4] ~^ image[1][6])} + {7'd0,(kernel[1][0] ~^ image[2][2])} + {7'd0,(kernel[1][1] ~^ image[2][3])} + {7'd0,(kernel[1][2] ~^ image[2][4])} + {7'd0,(kernel[1][3] ~^ image[2][5])} + {7'd0,(kernel[1][4] ~^ image[2][6])} + {7'd0,(kernel[2][0] ~^ image[3][2])} + {7'd0,(kernel[2][1] ~^ image[3][3])} + {7'd0,(kernel[2][2] ~^ image[3][4])} + {7'd0,(kernel[2][3] ~^ image[3][5])} + {7'd0,(kernel[2][4] ~^ image[3][6])} + {7'd0,(kernel[3][0] ~^ image[4][2])} + {7'd0,(kernel[3][1] ~^ image[4][3])} + {7'd0,(kernel[3][2] ~^ image[4][4])} + {7'd0,(kernel[3][3] ~^ image[4][5])} + {7'd0,(kernel[3][4] ~^ image[4][6])} + {7'd0,(kernel[4][0] ~^ image[5][2])} + {7'd0,(kernel[4][1] ~^ image[5][3])} + {7'd0,(kernel[4][2] ~^ image[5][4])} + {7'd0,(kernel[4][3] ~^ image[5][5])} + {7'd0,(kernel[4][4] ~^ image[5][6])};
assign out_fmap[1][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][3])} + {7'd0,(kernel[0][1] ~^ image[1][4])} + {7'd0,(kernel[0][2] ~^ image[1][5])} + {7'd0,(kernel[0][3] ~^ image[1][6])} + {7'd0,(kernel[0][4] ~^ image[1][7])} + {7'd0,(kernel[1][0] ~^ image[2][3])} + {7'd0,(kernel[1][1] ~^ image[2][4])} + {7'd0,(kernel[1][2] ~^ image[2][5])} + {7'd0,(kernel[1][3] ~^ image[2][6])} + {7'd0,(kernel[1][4] ~^ image[2][7])} + {7'd0,(kernel[2][0] ~^ image[3][3])} + {7'd0,(kernel[2][1] ~^ image[3][4])} + {7'd0,(kernel[2][2] ~^ image[3][5])} + {7'd0,(kernel[2][3] ~^ image[3][6])} + {7'd0,(kernel[2][4] ~^ image[3][7])} + {7'd0,(kernel[3][0] ~^ image[4][3])} + {7'd0,(kernel[3][1] ~^ image[4][4])} + {7'd0,(kernel[3][2] ~^ image[4][5])} + {7'd0,(kernel[3][3] ~^ image[4][6])} + {7'd0,(kernel[3][4] ~^ image[4][7])} + {7'd0,(kernel[4][0] ~^ image[5][3])} + {7'd0,(kernel[4][1] ~^ image[5][4])} + {7'd0,(kernel[4][2] ~^ image[5][5])} + {7'd0,(kernel[4][3] ~^ image[5][6])} + {7'd0,(kernel[4][4] ~^ image[5][7])};
assign out_fmap[1][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][4])} + {7'd0,(kernel[0][1] ~^ image[1][5])} + {7'd0,(kernel[0][2] ~^ image[1][6])} + {7'd0,(kernel[0][3] ~^ image[1][7])} + {7'd0,(kernel[0][4] ~^ image[1][8])} + {7'd0,(kernel[1][0] ~^ image[2][4])} + {7'd0,(kernel[1][1] ~^ image[2][5])} + {7'd0,(kernel[1][2] ~^ image[2][6])} + {7'd0,(kernel[1][3] ~^ image[2][7])} + {7'd0,(kernel[1][4] ~^ image[2][8])} + {7'd0,(kernel[2][0] ~^ image[3][4])} + {7'd0,(kernel[2][1] ~^ image[3][5])} + {7'd0,(kernel[2][2] ~^ image[3][6])} + {7'd0,(kernel[2][3] ~^ image[3][7])} + {7'd0,(kernel[2][4] ~^ image[3][8])} + {7'd0,(kernel[3][0] ~^ image[4][4])} + {7'd0,(kernel[3][1] ~^ image[4][5])} + {7'd0,(kernel[3][2] ~^ image[4][6])} + {7'd0,(kernel[3][3] ~^ image[4][7])} + {7'd0,(kernel[3][4] ~^ image[4][8])} + {7'd0,(kernel[4][0] ~^ image[5][4])} + {7'd0,(kernel[4][1] ~^ image[5][5])} + {7'd0,(kernel[4][2] ~^ image[5][6])} + {7'd0,(kernel[4][3] ~^ image[5][7])} + {7'd0,(kernel[4][4] ~^ image[5][8])};
assign out_fmap[1][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][5])} + {7'd0,(kernel[0][1] ~^ image[1][6])} + {7'd0,(kernel[0][2] ~^ image[1][7])} + {7'd0,(kernel[0][3] ~^ image[1][8])} + {7'd0,(kernel[0][4] ~^ image[1][9])} + {7'd0,(kernel[1][0] ~^ image[2][5])} + {7'd0,(kernel[1][1] ~^ image[2][6])} + {7'd0,(kernel[1][2] ~^ image[2][7])} + {7'd0,(kernel[1][3] ~^ image[2][8])} + {7'd0,(kernel[1][4] ~^ image[2][9])} + {7'd0,(kernel[2][0] ~^ image[3][5])} + {7'd0,(kernel[2][1] ~^ image[3][6])} + {7'd0,(kernel[2][2] ~^ image[3][7])} + {7'd0,(kernel[2][3] ~^ image[3][8])} + {7'd0,(kernel[2][4] ~^ image[3][9])} + {7'd0,(kernel[3][0] ~^ image[4][5])} + {7'd0,(kernel[3][1] ~^ image[4][6])} + {7'd0,(kernel[3][2] ~^ image[4][7])} + {7'd0,(kernel[3][3] ~^ image[4][8])} + {7'd0,(kernel[3][4] ~^ image[4][9])} + {7'd0,(kernel[4][0] ~^ image[5][5])} + {7'd0,(kernel[4][1] ~^ image[5][6])} + {7'd0,(kernel[4][2] ~^ image[5][7])} + {7'd0,(kernel[4][3] ~^ image[5][8])} + {7'd0,(kernel[4][4] ~^ image[5][9])};
assign out_fmap[1][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][6])} + {7'd0,(kernel[0][1] ~^ image[1][7])} + {7'd0,(kernel[0][2] ~^ image[1][8])} + {7'd0,(kernel[0][3] ~^ image[1][9])} + {7'd0,(kernel[0][4] ~^ image[1][10])} + {7'd0,(kernel[1][0] ~^ image[2][6])} + {7'd0,(kernel[1][1] ~^ image[2][7])} + {7'd0,(kernel[1][2] ~^ image[2][8])} + {7'd0,(kernel[1][3] ~^ image[2][9])} + {7'd0,(kernel[1][4] ~^ image[2][10])} + {7'd0,(kernel[2][0] ~^ image[3][6])} + {7'd0,(kernel[2][1] ~^ image[3][7])} + {7'd0,(kernel[2][2] ~^ image[3][8])} + {7'd0,(kernel[2][3] ~^ image[3][9])} + {7'd0,(kernel[2][4] ~^ image[3][10])} + {7'd0,(kernel[3][0] ~^ image[4][6])} + {7'd0,(kernel[3][1] ~^ image[4][7])} + {7'd0,(kernel[3][2] ~^ image[4][8])} + {7'd0,(kernel[3][3] ~^ image[4][9])} + {7'd0,(kernel[3][4] ~^ image[4][10])} + {7'd0,(kernel[4][0] ~^ image[5][6])} + {7'd0,(kernel[4][1] ~^ image[5][7])} + {7'd0,(kernel[4][2] ~^ image[5][8])} + {7'd0,(kernel[4][3] ~^ image[5][9])} + {7'd0,(kernel[4][4] ~^ image[5][10])};
assign out_fmap[1][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][7])} + {7'd0,(kernel[0][1] ~^ image[1][8])} + {7'd0,(kernel[0][2] ~^ image[1][9])} + {7'd0,(kernel[0][3] ~^ image[1][10])} + {7'd0,(kernel[0][4] ~^ image[1][11])} + {7'd0,(kernel[1][0] ~^ image[2][7])} + {7'd0,(kernel[1][1] ~^ image[2][8])} + {7'd0,(kernel[1][2] ~^ image[2][9])} + {7'd0,(kernel[1][3] ~^ image[2][10])} + {7'd0,(kernel[1][4] ~^ image[2][11])} + {7'd0,(kernel[2][0] ~^ image[3][7])} + {7'd0,(kernel[2][1] ~^ image[3][8])} + {7'd0,(kernel[2][2] ~^ image[3][9])} + {7'd0,(kernel[2][3] ~^ image[3][10])} + {7'd0,(kernel[2][4] ~^ image[3][11])} + {7'd0,(kernel[3][0] ~^ image[4][7])} + {7'd0,(kernel[3][1] ~^ image[4][8])} + {7'd0,(kernel[3][2] ~^ image[4][9])} + {7'd0,(kernel[3][3] ~^ image[4][10])} + {7'd0,(kernel[3][4] ~^ image[4][11])} + {7'd0,(kernel[4][0] ~^ image[5][7])} + {7'd0,(kernel[4][1] ~^ image[5][8])} + {7'd0,(kernel[4][2] ~^ image[5][9])} + {7'd0,(kernel[4][3] ~^ image[5][10])} + {7'd0,(kernel[4][4] ~^ image[5][11])};
assign out_fmap[1][8][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][8])} + {7'd0,(kernel[0][1] ~^ image[1][9])} + {7'd0,(kernel[0][2] ~^ image[1][10])} + {7'd0,(kernel[0][3] ~^ image[1][11])} + {7'd0,(kernel[0][4] ~^ image[1][12])} + {7'd0,(kernel[1][0] ~^ image[2][8])} + {7'd0,(kernel[1][1] ~^ image[2][9])} + {7'd0,(kernel[1][2] ~^ image[2][10])} + {7'd0,(kernel[1][3] ~^ image[2][11])} + {7'd0,(kernel[1][4] ~^ image[2][12])} + {7'd0,(kernel[2][0] ~^ image[3][8])} + {7'd0,(kernel[2][1] ~^ image[3][9])} + {7'd0,(kernel[2][2] ~^ image[3][10])} + {7'd0,(kernel[2][3] ~^ image[3][11])} + {7'd0,(kernel[2][4] ~^ image[3][12])} + {7'd0,(kernel[3][0] ~^ image[4][8])} + {7'd0,(kernel[3][1] ~^ image[4][9])} + {7'd0,(kernel[3][2] ~^ image[4][10])} + {7'd0,(kernel[3][3] ~^ image[4][11])} + {7'd0,(kernel[3][4] ~^ image[4][12])} + {7'd0,(kernel[4][0] ~^ image[5][8])} + {7'd0,(kernel[4][1] ~^ image[5][9])} + {7'd0,(kernel[4][2] ~^ image[5][10])} + {7'd0,(kernel[4][3] ~^ image[5][11])} + {7'd0,(kernel[4][4] ~^ image[5][12])};
assign out_fmap[1][9][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][9])} + {7'd0,(kernel[0][1] ~^ image[1][10])} + {7'd0,(kernel[0][2] ~^ image[1][11])} + {7'd0,(kernel[0][3] ~^ image[1][12])} + {7'd0,(kernel[0][4] ~^ image[1][13])} + {7'd0,(kernel[1][0] ~^ image[2][9])} + {7'd0,(kernel[1][1] ~^ image[2][10])} + {7'd0,(kernel[1][2] ~^ image[2][11])} + {7'd0,(kernel[1][3] ~^ image[2][12])} + {7'd0,(kernel[1][4] ~^ image[2][13])} + {7'd0,(kernel[2][0] ~^ image[3][9])} + {7'd0,(kernel[2][1] ~^ image[3][10])} + {7'd0,(kernel[2][2] ~^ image[3][11])} + {7'd0,(kernel[2][3] ~^ image[3][12])} + {7'd0,(kernel[2][4] ~^ image[3][13])} + {7'd0,(kernel[3][0] ~^ image[4][9])} + {7'd0,(kernel[3][1] ~^ image[4][10])} + {7'd0,(kernel[3][2] ~^ image[4][11])} + {7'd0,(kernel[3][3] ~^ image[4][12])} + {7'd0,(kernel[3][4] ~^ image[4][13])} + {7'd0,(kernel[4][0] ~^ image[5][9])} + {7'd0,(kernel[4][1] ~^ image[5][10])} + {7'd0,(kernel[4][2] ~^ image[5][11])} + {7'd0,(kernel[4][3] ~^ image[5][12])} + {7'd0,(kernel[4][4] ~^ image[5][13])};
assign out_fmap[1][10][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][10])} + {7'd0,(kernel[0][1] ~^ image[1][11])} + {7'd0,(kernel[0][2] ~^ image[1][12])} + {7'd0,(kernel[0][3] ~^ image[1][13])} + {7'd0,(kernel[0][4] ~^ image[1][14])} + {7'd0,(kernel[1][0] ~^ image[2][10])} + {7'd0,(kernel[1][1] ~^ image[2][11])} + {7'd0,(kernel[1][2] ~^ image[2][12])} + {7'd0,(kernel[1][3] ~^ image[2][13])} + {7'd0,(kernel[1][4] ~^ image[2][14])} + {7'd0,(kernel[2][0] ~^ image[3][10])} + {7'd0,(kernel[2][1] ~^ image[3][11])} + {7'd0,(kernel[2][2] ~^ image[3][12])} + {7'd0,(kernel[2][3] ~^ image[3][13])} + {7'd0,(kernel[2][4] ~^ image[3][14])} + {7'd0,(kernel[3][0] ~^ image[4][10])} + {7'd0,(kernel[3][1] ~^ image[4][11])} + {7'd0,(kernel[3][2] ~^ image[4][12])} + {7'd0,(kernel[3][3] ~^ image[4][13])} + {7'd0,(kernel[3][4] ~^ image[4][14])} + {7'd0,(kernel[4][0] ~^ image[5][10])} + {7'd0,(kernel[4][1] ~^ image[5][11])} + {7'd0,(kernel[4][2] ~^ image[5][12])} + {7'd0,(kernel[4][3] ~^ image[5][13])} + {7'd0,(kernel[4][4] ~^ image[5][14])};
assign out_fmap[1][11][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][11])} + {7'd0,(kernel[0][1] ~^ image[1][12])} + {7'd0,(kernel[0][2] ~^ image[1][13])} + {7'd0,(kernel[0][3] ~^ image[1][14])} + {7'd0,(kernel[0][4] ~^ image[1][15])} + {7'd0,(kernel[1][0] ~^ image[2][11])} + {7'd0,(kernel[1][1] ~^ image[2][12])} + {7'd0,(kernel[1][2] ~^ image[2][13])} + {7'd0,(kernel[1][3] ~^ image[2][14])} + {7'd0,(kernel[1][4] ~^ image[2][15])} + {7'd0,(kernel[2][0] ~^ image[3][11])} + {7'd0,(kernel[2][1] ~^ image[3][12])} + {7'd0,(kernel[2][2] ~^ image[3][13])} + {7'd0,(kernel[2][3] ~^ image[3][14])} + {7'd0,(kernel[2][4] ~^ image[3][15])} + {7'd0,(kernel[3][0] ~^ image[4][11])} + {7'd0,(kernel[3][1] ~^ image[4][12])} + {7'd0,(kernel[3][2] ~^ image[4][13])} + {7'd0,(kernel[3][3] ~^ image[4][14])} + {7'd0,(kernel[3][4] ~^ image[4][15])} + {7'd0,(kernel[4][0] ~^ image[5][11])} + {7'd0,(kernel[4][1] ~^ image[5][12])} + {7'd0,(kernel[4][2] ~^ image[5][13])} + {7'd0,(kernel[4][3] ~^ image[5][14])} + {7'd0,(kernel[4][4] ~^ image[5][15])};
assign out_fmap[1][12][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][12])} + {7'd0,(kernel[0][1] ~^ image[1][13])} + {7'd0,(kernel[0][2] ~^ image[1][14])} + {7'd0,(kernel[0][3] ~^ image[1][15])} + {7'd0,(kernel[0][4] ~^ image[1][16])} + {7'd0,(kernel[1][0] ~^ image[2][12])} + {7'd0,(kernel[1][1] ~^ image[2][13])} + {7'd0,(kernel[1][2] ~^ image[2][14])} + {7'd0,(kernel[1][3] ~^ image[2][15])} + {7'd0,(kernel[1][4] ~^ image[2][16])} + {7'd0,(kernel[2][0] ~^ image[3][12])} + {7'd0,(kernel[2][1] ~^ image[3][13])} + {7'd0,(kernel[2][2] ~^ image[3][14])} + {7'd0,(kernel[2][3] ~^ image[3][15])} + {7'd0,(kernel[2][4] ~^ image[3][16])} + {7'd0,(kernel[3][0] ~^ image[4][12])} + {7'd0,(kernel[3][1] ~^ image[4][13])} + {7'd0,(kernel[3][2] ~^ image[4][14])} + {7'd0,(kernel[3][3] ~^ image[4][15])} + {7'd0,(kernel[3][4] ~^ image[4][16])} + {7'd0,(kernel[4][0] ~^ image[5][12])} + {7'd0,(kernel[4][1] ~^ image[5][13])} + {7'd0,(kernel[4][2] ~^ image[5][14])} + {7'd0,(kernel[4][3] ~^ image[5][15])} + {7'd0,(kernel[4][4] ~^ image[5][16])};
assign out_fmap[1][13][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][13])} + {7'd0,(kernel[0][1] ~^ image[1][14])} + {7'd0,(kernel[0][2] ~^ image[1][15])} + {7'd0,(kernel[0][3] ~^ image[1][16])} + {7'd0,(kernel[0][4] ~^ image[1][17])} + {7'd0,(kernel[1][0] ~^ image[2][13])} + {7'd0,(kernel[1][1] ~^ image[2][14])} + {7'd0,(kernel[1][2] ~^ image[2][15])} + {7'd0,(kernel[1][3] ~^ image[2][16])} + {7'd0,(kernel[1][4] ~^ image[2][17])} + {7'd0,(kernel[2][0] ~^ image[3][13])} + {7'd0,(kernel[2][1] ~^ image[3][14])} + {7'd0,(kernel[2][2] ~^ image[3][15])} + {7'd0,(kernel[2][3] ~^ image[3][16])} + {7'd0,(kernel[2][4] ~^ image[3][17])} + {7'd0,(kernel[3][0] ~^ image[4][13])} + {7'd0,(kernel[3][1] ~^ image[4][14])} + {7'd0,(kernel[3][2] ~^ image[4][15])} + {7'd0,(kernel[3][3] ~^ image[4][16])} + {7'd0,(kernel[3][4] ~^ image[4][17])} + {7'd0,(kernel[4][0] ~^ image[5][13])} + {7'd0,(kernel[4][1] ~^ image[5][14])} + {7'd0,(kernel[4][2] ~^ image[5][15])} + {7'd0,(kernel[4][3] ~^ image[5][16])} + {7'd0,(kernel[4][4] ~^ image[5][17])};
assign out_fmap[1][14][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][14])} + {7'd0,(kernel[0][1] ~^ image[1][15])} + {7'd0,(kernel[0][2] ~^ image[1][16])} + {7'd0,(kernel[0][3] ~^ image[1][17])} + {7'd0,(kernel[0][4] ~^ image[1][18])} + {7'd0,(kernel[1][0] ~^ image[2][14])} + {7'd0,(kernel[1][1] ~^ image[2][15])} + {7'd0,(kernel[1][2] ~^ image[2][16])} + {7'd0,(kernel[1][3] ~^ image[2][17])} + {7'd0,(kernel[1][4] ~^ image[2][18])} + {7'd0,(kernel[2][0] ~^ image[3][14])} + {7'd0,(kernel[2][1] ~^ image[3][15])} + {7'd0,(kernel[2][2] ~^ image[3][16])} + {7'd0,(kernel[2][3] ~^ image[3][17])} + {7'd0,(kernel[2][4] ~^ image[3][18])} + {7'd0,(kernel[3][0] ~^ image[4][14])} + {7'd0,(kernel[3][1] ~^ image[4][15])} + {7'd0,(kernel[3][2] ~^ image[4][16])} + {7'd0,(kernel[3][3] ~^ image[4][17])} + {7'd0,(kernel[3][4] ~^ image[4][18])} + {7'd0,(kernel[4][0] ~^ image[5][14])} + {7'd0,(kernel[4][1] ~^ image[5][15])} + {7'd0,(kernel[4][2] ~^ image[5][16])} + {7'd0,(kernel[4][3] ~^ image[5][17])} + {7'd0,(kernel[4][4] ~^ image[5][18])};
assign out_fmap[1][15][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][15])} + {7'd0,(kernel[0][1] ~^ image[1][16])} + {7'd0,(kernel[0][2] ~^ image[1][17])} + {7'd0,(kernel[0][3] ~^ image[1][18])} + {7'd0,(kernel[0][4] ~^ image[1][19])} + {7'd0,(kernel[1][0] ~^ image[2][15])} + {7'd0,(kernel[1][1] ~^ image[2][16])} + {7'd0,(kernel[1][2] ~^ image[2][17])} + {7'd0,(kernel[1][3] ~^ image[2][18])} + {7'd0,(kernel[1][4] ~^ image[2][19])} + {7'd0,(kernel[2][0] ~^ image[3][15])} + {7'd0,(kernel[2][1] ~^ image[3][16])} + {7'd0,(kernel[2][2] ~^ image[3][17])} + {7'd0,(kernel[2][3] ~^ image[3][18])} + {7'd0,(kernel[2][4] ~^ image[3][19])} + {7'd0,(kernel[3][0] ~^ image[4][15])} + {7'd0,(kernel[3][1] ~^ image[4][16])} + {7'd0,(kernel[3][2] ~^ image[4][17])} + {7'd0,(kernel[3][3] ~^ image[4][18])} + {7'd0,(kernel[3][4] ~^ image[4][19])} + {7'd0,(kernel[4][0] ~^ image[5][15])} + {7'd0,(kernel[4][1] ~^ image[5][16])} + {7'd0,(kernel[4][2] ~^ image[5][17])} + {7'd0,(kernel[4][3] ~^ image[5][18])} + {7'd0,(kernel[4][4] ~^ image[5][19])};
assign out_fmap[1][16][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][16])} + {7'd0,(kernel[0][1] ~^ image[1][17])} + {7'd0,(kernel[0][2] ~^ image[1][18])} + {7'd0,(kernel[0][3] ~^ image[1][19])} + {7'd0,(kernel[0][4] ~^ image[1][20])} + {7'd0,(kernel[1][0] ~^ image[2][16])} + {7'd0,(kernel[1][1] ~^ image[2][17])} + {7'd0,(kernel[1][2] ~^ image[2][18])} + {7'd0,(kernel[1][3] ~^ image[2][19])} + {7'd0,(kernel[1][4] ~^ image[2][20])} + {7'd0,(kernel[2][0] ~^ image[3][16])} + {7'd0,(kernel[2][1] ~^ image[3][17])} + {7'd0,(kernel[2][2] ~^ image[3][18])} + {7'd0,(kernel[2][3] ~^ image[3][19])} + {7'd0,(kernel[2][4] ~^ image[3][20])} + {7'd0,(kernel[3][0] ~^ image[4][16])} + {7'd0,(kernel[3][1] ~^ image[4][17])} + {7'd0,(kernel[3][2] ~^ image[4][18])} + {7'd0,(kernel[3][3] ~^ image[4][19])} + {7'd0,(kernel[3][4] ~^ image[4][20])} + {7'd0,(kernel[4][0] ~^ image[5][16])} + {7'd0,(kernel[4][1] ~^ image[5][17])} + {7'd0,(kernel[4][2] ~^ image[5][18])} + {7'd0,(kernel[4][3] ~^ image[5][19])} + {7'd0,(kernel[4][4] ~^ image[5][20])};
assign out_fmap[1][17][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][17])} + {7'd0,(kernel[0][1] ~^ image[1][18])} + {7'd0,(kernel[0][2] ~^ image[1][19])} + {7'd0,(kernel[0][3] ~^ image[1][20])} + {7'd0,(kernel[0][4] ~^ image[1][21])} + {7'd0,(kernel[1][0] ~^ image[2][17])} + {7'd0,(kernel[1][1] ~^ image[2][18])} + {7'd0,(kernel[1][2] ~^ image[2][19])} + {7'd0,(kernel[1][3] ~^ image[2][20])} + {7'd0,(kernel[1][4] ~^ image[2][21])} + {7'd0,(kernel[2][0] ~^ image[3][17])} + {7'd0,(kernel[2][1] ~^ image[3][18])} + {7'd0,(kernel[2][2] ~^ image[3][19])} + {7'd0,(kernel[2][3] ~^ image[3][20])} + {7'd0,(kernel[2][4] ~^ image[3][21])} + {7'd0,(kernel[3][0] ~^ image[4][17])} + {7'd0,(kernel[3][1] ~^ image[4][18])} + {7'd0,(kernel[3][2] ~^ image[4][19])} + {7'd0,(kernel[3][3] ~^ image[4][20])} + {7'd0,(kernel[3][4] ~^ image[4][21])} + {7'd0,(kernel[4][0] ~^ image[5][17])} + {7'd0,(kernel[4][1] ~^ image[5][18])} + {7'd0,(kernel[4][2] ~^ image[5][19])} + {7'd0,(kernel[4][3] ~^ image[5][20])} + {7'd0,(kernel[4][4] ~^ image[5][21])};
assign out_fmap[1][18][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][18])} + {7'd0,(kernel[0][1] ~^ image[1][19])} + {7'd0,(kernel[0][2] ~^ image[1][20])} + {7'd0,(kernel[0][3] ~^ image[1][21])} + {7'd0,(kernel[0][4] ~^ image[1][22])} + {7'd0,(kernel[1][0] ~^ image[2][18])} + {7'd0,(kernel[1][1] ~^ image[2][19])} + {7'd0,(kernel[1][2] ~^ image[2][20])} + {7'd0,(kernel[1][3] ~^ image[2][21])} + {7'd0,(kernel[1][4] ~^ image[2][22])} + {7'd0,(kernel[2][0] ~^ image[3][18])} + {7'd0,(kernel[2][1] ~^ image[3][19])} + {7'd0,(kernel[2][2] ~^ image[3][20])} + {7'd0,(kernel[2][3] ~^ image[3][21])} + {7'd0,(kernel[2][4] ~^ image[3][22])} + {7'd0,(kernel[3][0] ~^ image[4][18])} + {7'd0,(kernel[3][1] ~^ image[4][19])} + {7'd0,(kernel[3][2] ~^ image[4][20])} + {7'd0,(kernel[3][3] ~^ image[4][21])} + {7'd0,(kernel[3][4] ~^ image[4][22])} + {7'd0,(kernel[4][0] ~^ image[5][18])} + {7'd0,(kernel[4][1] ~^ image[5][19])} + {7'd0,(kernel[4][2] ~^ image[5][20])} + {7'd0,(kernel[4][3] ~^ image[5][21])} + {7'd0,(kernel[4][4] ~^ image[5][22])};
assign out_fmap[1][19][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][19])} + {7'd0,(kernel[0][1] ~^ image[1][20])} + {7'd0,(kernel[0][2] ~^ image[1][21])} + {7'd0,(kernel[0][3] ~^ image[1][22])} + {7'd0,(kernel[0][4] ~^ image[1][23])} + {7'd0,(kernel[1][0] ~^ image[2][19])} + {7'd0,(kernel[1][1] ~^ image[2][20])} + {7'd0,(kernel[1][2] ~^ image[2][21])} + {7'd0,(kernel[1][3] ~^ image[2][22])} + {7'd0,(kernel[1][4] ~^ image[2][23])} + {7'd0,(kernel[2][0] ~^ image[3][19])} + {7'd0,(kernel[2][1] ~^ image[3][20])} + {7'd0,(kernel[2][2] ~^ image[3][21])} + {7'd0,(kernel[2][3] ~^ image[3][22])} + {7'd0,(kernel[2][4] ~^ image[3][23])} + {7'd0,(kernel[3][0] ~^ image[4][19])} + {7'd0,(kernel[3][1] ~^ image[4][20])} + {7'd0,(kernel[3][2] ~^ image[4][21])} + {7'd0,(kernel[3][3] ~^ image[4][22])} + {7'd0,(kernel[3][4] ~^ image[4][23])} + {7'd0,(kernel[4][0] ~^ image[5][19])} + {7'd0,(kernel[4][1] ~^ image[5][20])} + {7'd0,(kernel[4][2] ~^ image[5][21])} + {7'd0,(kernel[4][3] ~^ image[5][22])} + {7'd0,(kernel[4][4] ~^ image[5][23])};
assign out_fmap[1][20][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][20])} + {7'd0,(kernel[0][1] ~^ image[1][21])} + {7'd0,(kernel[0][2] ~^ image[1][22])} + {7'd0,(kernel[0][3] ~^ image[1][23])} + {7'd0,(kernel[0][4] ~^ image[1][24])} + {7'd0,(kernel[1][0] ~^ image[2][20])} + {7'd0,(kernel[1][1] ~^ image[2][21])} + {7'd0,(kernel[1][2] ~^ image[2][22])} + {7'd0,(kernel[1][3] ~^ image[2][23])} + {7'd0,(kernel[1][4] ~^ image[2][24])} + {7'd0,(kernel[2][0] ~^ image[3][20])} + {7'd0,(kernel[2][1] ~^ image[3][21])} + {7'd0,(kernel[2][2] ~^ image[3][22])} + {7'd0,(kernel[2][3] ~^ image[3][23])} + {7'd0,(kernel[2][4] ~^ image[3][24])} + {7'd0,(kernel[3][0] ~^ image[4][20])} + {7'd0,(kernel[3][1] ~^ image[4][21])} + {7'd0,(kernel[3][2] ~^ image[4][22])} + {7'd0,(kernel[3][3] ~^ image[4][23])} + {7'd0,(kernel[3][4] ~^ image[4][24])} + {7'd0,(kernel[4][0] ~^ image[5][20])} + {7'd0,(kernel[4][1] ~^ image[5][21])} + {7'd0,(kernel[4][2] ~^ image[5][22])} + {7'd0,(kernel[4][3] ~^ image[5][23])} + {7'd0,(kernel[4][4] ~^ image[5][24])};
assign out_fmap[1][21][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][21])} + {7'd0,(kernel[0][1] ~^ image[1][22])} + {7'd0,(kernel[0][2] ~^ image[1][23])} + {7'd0,(kernel[0][3] ~^ image[1][24])} + {7'd0,(kernel[0][4] ~^ image[1][25])} + {7'd0,(kernel[1][0] ~^ image[2][21])} + {7'd0,(kernel[1][1] ~^ image[2][22])} + {7'd0,(kernel[1][2] ~^ image[2][23])} + {7'd0,(kernel[1][3] ~^ image[2][24])} + {7'd0,(kernel[1][4] ~^ image[2][25])} + {7'd0,(kernel[2][0] ~^ image[3][21])} + {7'd0,(kernel[2][1] ~^ image[3][22])} + {7'd0,(kernel[2][2] ~^ image[3][23])} + {7'd0,(kernel[2][3] ~^ image[3][24])} + {7'd0,(kernel[2][4] ~^ image[3][25])} + {7'd0,(kernel[3][0] ~^ image[4][21])} + {7'd0,(kernel[3][1] ~^ image[4][22])} + {7'd0,(kernel[3][2] ~^ image[4][23])} + {7'd0,(kernel[3][3] ~^ image[4][24])} + {7'd0,(kernel[3][4] ~^ image[4][25])} + {7'd0,(kernel[4][0] ~^ image[5][21])} + {7'd0,(kernel[4][1] ~^ image[5][22])} + {7'd0,(kernel[4][2] ~^ image[5][23])} + {7'd0,(kernel[4][3] ~^ image[5][24])} + {7'd0,(kernel[4][4] ~^ image[5][25])};
assign out_fmap[1][22][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][22])} + {7'd0,(kernel[0][1] ~^ image[1][23])} + {7'd0,(kernel[0][2] ~^ image[1][24])} + {7'd0,(kernel[0][3] ~^ image[1][25])} + {7'd0,(kernel[0][4] ~^ image[1][26])} + {7'd0,(kernel[1][0] ~^ image[2][22])} + {7'd0,(kernel[1][1] ~^ image[2][23])} + {7'd0,(kernel[1][2] ~^ image[2][24])} + {7'd0,(kernel[1][3] ~^ image[2][25])} + {7'd0,(kernel[1][4] ~^ image[2][26])} + {7'd0,(kernel[2][0] ~^ image[3][22])} + {7'd0,(kernel[2][1] ~^ image[3][23])} + {7'd0,(kernel[2][2] ~^ image[3][24])} + {7'd0,(kernel[2][3] ~^ image[3][25])} + {7'd0,(kernel[2][4] ~^ image[3][26])} + {7'd0,(kernel[3][0] ~^ image[4][22])} + {7'd0,(kernel[3][1] ~^ image[4][23])} + {7'd0,(kernel[3][2] ~^ image[4][24])} + {7'd0,(kernel[3][3] ~^ image[4][25])} + {7'd0,(kernel[3][4] ~^ image[4][26])} + {7'd0,(kernel[4][0] ~^ image[5][22])} + {7'd0,(kernel[4][1] ~^ image[5][23])} + {7'd0,(kernel[4][2] ~^ image[5][24])} + {7'd0,(kernel[4][3] ~^ image[5][25])} + {7'd0,(kernel[4][4] ~^ image[5][26])};
assign out_fmap[1][23][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[1][23])} + {7'd0,(kernel[0][1] ~^ image[1][24])} + {7'd0,(kernel[0][2] ~^ image[1][25])} + {7'd0,(kernel[0][3] ~^ image[1][26])} + {7'd0,(kernel[0][4] ~^ image[1][27])} + {7'd0,(kernel[1][0] ~^ image[2][23])} + {7'd0,(kernel[1][1] ~^ image[2][24])} + {7'd0,(kernel[1][2] ~^ image[2][25])} + {7'd0,(kernel[1][3] ~^ image[2][26])} + {7'd0,(kernel[1][4] ~^ image[2][27])} + {7'd0,(kernel[2][0] ~^ image[3][23])} + {7'd0,(kernel[2][1] ~^ image[3][24])} + {7'd0,(kernel[2][2] ~^ image[3][25])} + {7'd0,(kernel[2][3] ~^ image[3][26])} + {7'd0,(kernel[2][4] ~^ image[3][27])} + {7'd0,(kernel[3][0] ~^ image[4][23])} + {7'd0,(kernel[3][1] ~^ image[4][24])} + {7'd0,(kernel[3][2] ~^ image[4][25])} + {7'd0,(kernel[3][3] ~^ image[4][26])} + {7'd0,(kernel[3][4] ~^ image[4][27])} + {7'd0,(kernel[4][0] ~^ image[5][23])} + {7'd0,(kernel[4][1] ~^ image[5][24])} + {7'd0,(kernel[4][2] ~^ image[5][25])} + {7'd0,(kernel[4][3] ~^ image[5][26])} + {7'd0,(kernel[4][4] ~^ image[5][27])};
assign out_fmap[2][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][0])} + {7'd0,(kernel[0][1] ~^ image[2][1])} + {7'd0,(kernel[0][2] ~^ image[2][2])} + {7'd0,(kernel[0][3] ~^ image[2][3])} + {7'd0,(kernel[0][4] ~^ image[2][4])} + {7'd0,(kernel[1][0] ~^ image[3][0])} + {7'd0,(kernel[1][1] ~^ image[3][1])} + {7'd0,(kernel[1][2] ~^ image[3][2])} + {7'd0,(kernel[1][3] ~^ image[3][3])} + {7'd0,(kernel[1][4] ~^ image[3][4])} + {7'd0,(kernel[2][0] ~^ image[4][0])} + {7'd0,(kernel[2][1] ~^ image[4][1])} + {7'd0,(kernel[2][2] ~^ image[4][2])} + {7'd0,(kernel[2][3] ~^ image[4][3])} + {7'd0,(kernel[2][4] ~^ image[4][4])} + {7'd0,(kernel[3][0] ~^ image[5][0])} + {7'd0,(kernel[3][1] ~^ image[5][1])} + {7'd0,(kernel[3][2] ~^ image[5][2])} + {7'd0,(kernel[3][3] ~^ image[5][3])} + {7'd0,(kernel[3][4] ~^ image[5][4])} + {7'd0,(kernel[4][0] ~^ image[6][0])} + {7'd0,(kernel[4][1] ~^ image[6][1])} + {7'd0,(kernel[4][2] ~^ image[6][2])} + {7'd0,(kernel[4][3] ~^ image[6][3])} + {7'd0,(kernel[4][4] ~^ image[6][4])};
assign out_fmap[2][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][1])} + {7'd0,(kernel[0][1] ~^ image[2][2])} + {7'd0,(kernel[0][2] ~^ image[2][3])} + {7'd0,(kernel[0][3] ~^ image[2][4])} + {7'd0,(kernel[0][4] ~^ image[2][5])} + {7'd0,(kernel[1][0] ~^ image[3][1])} + {7'd0,(kernel[1][1] ~^ image[3][2])} + {7'd0,(kernel[1][2] ~^ image[3][3])} + {7'd0,(kernel[1][3] ~^ image[3][4])} + {7'd0,(kernel[1][4] ~^ image[3][5])} + {7'd0,(kernel[2][0] ~^ image[4][1])} + {7'd0,(kernel[2][1] ~^ image[4][2])} + {7'd0,(kernel[2][2] ~^ image[4][3])} + {7'd0,(kernel[2][3] ~^ image[4][4])} + {7'd0,(kernel[2][4] ~^ image[4][5])} + {7'd0,(kernel[3][0] ~^ image[5][1])} + {7'd0,(kernel[3][1] ~^ image[5][2])} + {7'd0,(kernel[3][2] ~^ image[5][3])} + {7'd0,(kernel[3][3] ~^ image[5][4])} + {7'd0,(kernel[3][4] ~^ image[5][5])} + {7'd0,(kernel[4][0] ~^ image[6][1])} + {7'd0,(kernel[4][1] ~^ image[6][2])} + {7'd0,(kernel[4][2] ~^ image[6][3])} + {7'd0,(kernel[4][3] ~^ image[6][4])} + {7'd0,(kernel[4][4] ~^ image[6][5])};
assign out_fmap[2][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][2])} + {7'd0,(kernel[0][1] ~^ image[2][3])} + {7'd0,(kernel[0][2] ~^ image[2][4])} + {7'd0,(kernel[0][3] ~^ image[2][5])} + {7'd0,(kernel[0][4] ~^ image[2][6])} + {7'd0,(kernel[1][0] ~^ image[3][2])} + {7'd0,(kernel[1][1] ~^ image[3][3])} + {7'd0,(kernel[1][2] ~^ image[3][4])} + {7'd0,(kernel[1][3] ~^ image[3][5])} + {7'd0,(kernel[1][4] ~^ image[3][6])} + {7'd0,(kernel[2][0] ~^ image[4][2])} + {7'd0,(kernel[2][1] ~^ image[4][3])} + {7'd0,(kernel[2][2] ~^ image[4][4])} + {7'd0,(kernel[2][3] ~^ image[4][5])} + {7'd0,(kernel[2][4] ~^ image[4][6])} + {7'd0,(kernel[3][0] ~^ image[5][2])} + {7'd0,(kernel[3][1] ~^ image[5][3])} + {7'd0,(kernel[3][2] ~^ image[5][4])} + {7'd0,(kernel[3][3] ~^ image[5][5])} + {7'd0,(kernel[3][4] ~^ image[5][6])} + {7'd0,(kernel[4][0] ~^ image[6][2])} + {7'd0,(kernel[4][1] ~^ image[6][3])} + {7'd0,(kernel[4][2] ~^ image[6][4])} + {7'd0,(kernel[4][3] ~^ image[6][5])} + {7'd0,(kernel[4][4] ~^ image[6][6])};
assign out_fmap[2][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][3])} + {7'd0,(kernel[0][1] ~^ image[2][4])} + {7'd0,(kernel[0][2] ~^ image[2][5])} + {7'd0,(kernel[0][3] ~^ image[2][6])} + {7'd0,(kernel[0][4] ~^ image[2][7])} + {7'd0,(kernel[1][0] ~^ image[3][3])} + {7'd0,(kernel[1][1] ~^ image[3][4])} + {7'd0,(kernel[1][2] ~^ image[3][5])} + {7'd0,(kernel[1][3] ~^ image[3][6])} + {7'd0,(kernel[1][4] ~^ image[3][7])} + {7'd0,(kernel[2][0] ~^ image[4][3])} + {7'd0,(kernel[2][1] ~^ image[4][4])} + {7'd0,(kernel[2][2] ~^ image[4][5])} + {7'd0,(kernel[2][3] ~^ image[4][6])} + {7'd0,(kernel[2][4] ~^ image[4][7])} + {7'd0,(kernel[3][0] ~^ image[5][3])} + {7'd0,(kernel[3][1] ~^ image[5][4])} + {7'd0,(kernel[3][2] ~^ image[5][5])} + {7'd0,(kernel[3][3] ~^ image[5][6])} + {7'd0,(kernel[3][4] ~^ image[5][7])} + {7'd0,(kernel[4][0] ~^ image[6][3])} + {7'd0,(kernel[4][1] ~^ image[6][4])} + {7'd0,(kernel[4][2] ~^ image[6][5])} + {7'd0,(kernel[4][3] ~^ image[6][6])} + {7'd0,(kernel[4][4] ~^ image[6][7])};
assign out_fmap[2][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][4])} + {7'd0,(kernel[0][1] ~^ image[2][5])} + {7'd0,(kernel[0][2] ~^ image[2][6])} + {7'd0,(kernel[0][3] ~^ image[2][7])} + {7'd0,(kernel[0][4] ~^ image[2][8])} + {7'd0,(kernel[1][0] ~^ image[3][4])} + {7'd0,(kernel[1][1] ~^ image[3][5])} + {7'd0,(kernel[1][2] ~^ image[3][6])} + {7'd0,(kernel[1][3] ~^ image[3][7])} + {7'd0,(kernel[1][4] ~^ image[3][8])} + {7'd0,(kernel[2][0] ~^ image[4][4])} + {7'd0,(kernel[2][1] ~^ image[4][5])} + {7'd0,(kernel[2][2] ~^ image[4][6])} + {7'd0,(kernel[2][3] ~^ image[4][7])} + {7'd0,(kernel[2][4] ~^ image[4][8])} + {7'd0,(kernel[3][0] ~^ image[5][4])} + {7'd0,(kernel[3][1] ~^ image[5][5])} + {7'd0,(kernel[3][2] ~^ image[5][6])} + {7'd0,(kernel[3][3] ~^ image[5][7])} + {7'd0,(kernel[3][4] ~^ image[5][8])} + {7'd0,(kernel[4][0] ~^ image[6][4])} + {7'd0,(kernel[4][1] ~^ image[6][5])} + {7'd0,(kernel[4][2] ~^ image[6][6])} + {7'd0,(kernel[4][3] ~^ image[6][7])} + {7'd0,(kernel[4][4] ~^ image[6][8])};
assign out_fmap[2][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][5])} + {7'd0,(kernel[0][1] ~^ image[2][6])} + {7'd0,(kernel[0][2] ~^ image[2][7])} + {7'd0,(kernel[0][3] ~^ image[2][8])} + {7'd0,(kernel[0][4] ~^ image[2][9])} + {7'd0,(kernel[1][0] ~^ image[3][5])} + {7'd0,(kernel[1][1] ~^ image[3][6])} + {7'd0,(kernel[1][2] ~^ image[3][7])} + {7'd0,(kernel[1][3] ~^ image[3][8])} + {7'd0,(kernel[1][4] ~^ image[3][9])} + {7'd0,(kernel[2][0] ~^ image[4][5])} + {7'd0,(kernel[2][1] ~^ image[4][6])} + {7'd0,(kernel[2][2] ~^ image[4][7])} + {7'd0,(kernel[2][3] ~^ image[4][8])} + {7'd0,(kernel[2][4] ~^ image[4][9])} + {7'd0,(kernel[3][0] ~^ image[5][5])} + {7'd0,(kernel[3][1] ~^ image[5][6])} + {7'd0,(kernel[3][2] ~^ image[5][7])} + {7'd0,(kernel[3][3] ~^ image[5][8])} + {7'd0,(kernel[3][4] ~^ image[5][9])} + {7'd0,(kernel[4][0] ~^ image[6][5])} + {7'd0,(kernel[4][1] ~^ image[6][6])} + {7'd0,(kernel[4][2] ~^ image[6][7])} + {7'd0,(kernel[4][3] ~^ image[6][8])} + {7'd0,(kernel[4][4] ~^ image[6][9])};
assign out_fmap[2][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][6])} + {7'd0,(kernel[0][1] ~^ image[2][7])} + {7'd0,(kernel[0][2] ~^ image[2][8])} + {7'd0,(kernel[0][3] ~^ image[2][9])} + {7'd0,(kernel[0][4] ~^ image[2][10])} + {7'd0,(kernel[1][0] ~^ image[3][6])} + {7'd0,(kernel[1][1] ~^ image[3][7])} + {7'd0,(kernel[1][2] ~^ image[3][8])} + {7'd0,(kernel[1][3] ~^ image[3][9])} + {7'd0,(kernel[1][4] ~^ image[3][10])} + {7'd0,(kernel[2][0] ~^ image[4][6])} + {7'd0,(kernel[2][1] ~^ image[4][7])} + {7'd0,(kernel[2][2] ~^ image[4][8])} + {7'd0,(kernel[2][3] ~^ image[4][9])} + {7'd0,(kernel[2][4] ~^ image[4][10])} + {7'd0,(kernel[3][0] ~^ image[5][6])} + {7'd0,(kernel[3][1] ~^ image[5][7])} + {7'd0,(kernel[3][2] ~^ image[5][8])} + {7'd0,(kernel[3][3] ~^ image[5][9])} + {7'd0,(kernel[3][4] ~^ image[5][10])} + {7'd0,(kernel[4][0] ~^ image[6][6])} + {7'd0,(kernel[4][1] ~^ image[6][7])} + {7'd0,(kernel[4][2] ~^ image[6][8])} + {7'd0,(kernel[4][3] ~^ image[6][9])} + {7'd0,(kernel[4][4] ~^ image[6][10])};
assign out_fmap[2][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][7])} + {7'd0,(kernel[0][1] ~^ image[2][8])} + {7'd0,(kernel[0][2] ~^ image[2][9])} + {7'd0,(kernel[0][3] ~^ image[2][10])} + {7'd0,(kernel[0][4] ~^ image[2][11])} + {7'd0,(kernel[1][0] ~^ image[3][7])} + {7'd0,(kernel[1][1] ~^ image[3][8])} + {7'd0,(kernel[1][2] ~^ image[3][9])} + {7'd0,(kernel[1][3] ~^ image[3][10])} + {7'd0,(kernel[1][4] ~^ image[3][11])} + {7'd0,(kernel[2][0] ~^ image[4][7])} + {7'd0,(kernel[2][1] ~^ image[4][8])} + {7'd0,(kernel[2][2] ~^ image[4][9])} + {7'd0,(kernel[2][3] ~^ image[4][10])} + {7'd0,(kernel[2][4] ~^ image[4][11])} + {7'd0,(kernel[3][0] ~^ image[5][7])} + {7'd0,(kernel[3][1] ~^ image[5][8])} + {7'd0,(kernel[3][2] ~^ image[5][9])} + {7'd0,(kernel[3][3] ~^ image[5][10])} + {7'd0,(kernel[3][4] ~^ image[5][11])} + {7'd0,(kernel[4][0] ~^ image[6][7])} + {7'd0,(kernel[4][1] ~^ image[6][8])} + {7'd0,(kernel[4][2] ~^ image[6][9])} + {7'd0,(kernel[4][3] ~^ image[6][10])} + {7'd0,(kernel[4][4] ~^ image[6][11])};
assign out_fmap[2][8][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][8])} + {7'd0,(kernel[0][1] ~^ image[2][9])} + {7'd0,(kernel[0][2] ~^ image[2][10])} + {7'd0,(kernel[0][3] ~^ image[2][11])} + {7'd0,(kernel[0][4] ~^ image[2][12])} + {7'd0,(kernel[1][0] ~^ image[3][8])} + {7'd0,(kernel[1][1] ~^ image[3][9])} + {7'd0,(kernel[1][2] ~^ image[3][10])} + {7'd0,(kernel[1][3] ~^ image[3][11])} + {7'd0,(kernel[1][4] ~^ image[3][12])} + {7'd0,(kernel[2][0] ~^ image[4][8])} + {7'd0,(kernel[2][1] ~^ image[4][9])} + {7'd0,(kernel[2][2] ~^ image[4][10])} + {7'd0,(kernel[2][3] ~^ image[4][11])} + {7'd0,(kernel[2][4] ~^ image[4][12])} + {7'd0,(kernel[3][0] ~^ image[5][8])} + {7'd0,(kernel[3][1] ~^ image[5][9])} + {7'd0,(kernel[3][2] ~^ image[5][10])} + {7'd0,(kernel[3][3] ~^ image[5][11])} + {7'd0,(kernel[3][4] ~^ image[5][12])} + {7'd0,(kernel[4][0] ~^ image[6][8])} + {7'd0,(kernel[4][1] ~^ image[6][9])} + {7'd0,(kernel[4][2] ~^ image[6][10])} + {7'd0,(kernel[4][3] ~^ image[6][11])} + {7'd0,(kernel[4][4] ~^ image[6][12])};
assign out_fmap[2][9][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][9])} + {7'd0,(kernel[0][1] ~^ image[2][10])} + {7'd0,(kernel[0][2] ~^ image[2][11])} + {7'd0,(kernel[0][3] ~^ image[2][12])} + {7'd0,(kernel[0][4] ~^ image[2][13])} + {7'd0,(kernel[1][0] ~^ image[3][9])} + {7'd0,(kernel[1][1] ~^ image[3][10])} + {7'd0,(kernel[1][2] ~^ image[3][11])} + {7'd0,(kernel[1][3] ~^ image[3][12])} + {7'd0,(kernel[1][4] ~^ image[3][13])} + {7'd0,(kernel[2][0] ~^ image[4][9])} + {7'd0,(kernel[2][1] ~^ image[4][10])} + {7'd0,(kernel[2][2] ~^ image[4][11])} + {7'd0,(kernel[2][3] ~^ image[4][12])} + {7'd0,(kernel[2][4] ~^ image[4][13])} + {7'd0,(kernel[3][0] ~^ image[5][9])} + {7'd0,(kernel[3][1] ~^ image[5][10])} + {7'd0,(kernel[3][2] ~^ image[5][11])} + {7'd0,(kernel[3][3] ~^ image[5][12])} + {7'd0,(kernel[3][4] ~^ image[5][13])} + {7'd0,(kernel[4][0] ~^ image[6][9])} + {7'd0,(kernel[4][1] ~^ image[6][10])} + {7'd0,(kernel[4][2] ~^ image[6][11])} + {7'd0,(kernel[4][3] ~^ image[6][12])} + {7'd0,(kernel[4][4] ~^ image[6][13])};
assign out_fmap[2][10][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][10])} + {7'd0,(kernel[0][1] ~^ image[2][11])} + {7'd0,(kernel[0][2] ~^ image[2][12])} + {7'd0,(kernel[0][3] ~^ image[2][13])} + {7'd0,(kernel[0][4] ~^ image[2][14])} + {7'd0,(kernel[1][0] ~^ image[3][10])} + {7'd0,(kernel[1][1] ~^ image[3][11])} + {7'd0,(kernel[1][2] ~^ image[3][12])} + {7'd0,(kernel[1][3] ~^ image[3][13])} + {7'd0,(kernel[1][4] ~^ image[3][14])} + {7'd0,(kernel[2][0] ~^ image[4][10])} + {7'd0,(kernel[2][1] ~^ image[4][11])} + {7'd0,(kernel[2][2] ~^ image[4][12])} + {7'd0,(kernel[2][3] ~^ image[4][13])} + {7'd0,(kernel[2][4] ~^ image[4][14])} + {7'd0,(kernel[3][0] ~^ image[5][10])} + {7'd0,(kernel[3][1] ~^ image[5][11])} + {7'd0,(kernel[3][2] ~^ image[5][12])} + {7'd0,(kernel[3][3] ~^ image[5][13])} + {7'd0,(kernel[3][4] ~^ image[5][14])} + {7'd0,(kernel[4][0] ~^ image[6][10])} + {7'd0,(kernel[4][1] ~^ image[6][11])} + {7'd0,(kernel[4][2] ~^ image[6][12])} + {7'd0,(kernel[4][3] ~^ image[6][13])} + {7'd0,(kernel[4][4] ~^ image[6][14])};
assign out_fmap[2][11][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][11])} + {7'd0,(kernel[0][1] ~^ image[2][12])} + {7'd0,(kernel[0][2] ~^ image[2][13])} + {7'd0,(kernel[0][3] ~^ image[2][14])} + {7'd0,(kernel[0][4] ~^ image[2][15])} + {7'd0,(kernel[1][0] ~^ image[3][11])} + {7'd0,(kernel[1][1] ~^ image[3][12])} + {7'd0,(kernel[1][2] ~^ image[3][13])} + {7'd0,(kernel[1][3] ~^ image[3][14])} + {7'd0,(kernel[1][4] ~^ image[3][15])} + {7'd0,(kernel[2][0] ~^ image[4][11])} + {7'd0,(kernel[2][1] ~^ image[4][12])} + {7'd0,(kernel[2][2] ~^ image[4][13])} + {7'd0,(kernel[2][3] ~^ image[4][14])} + {7'd0,(kernel[2][4] ~^ image[4][15])} + {7'd0,(kernel[3][0] ~^ image[5][11])} + {7'd0,(kernel[3][1] ~^ image[5][12])} + {7'd0,(kernel[3][2] ~^ image[5][13])} + {7'd0,(kernel[3][3] ~^ image[5][14])} + {7'd0,(kernel[3][4] ~^ image[5][15])} + {7'd0,(kernel[4][0] ~^ image[6][11])} + {7'd0,(kernel[4][1] ~^ image[6][12])} + {7'd0,(kernel[4][2] ~^ image[6][13])} + {7'd0,(kernel[4][3] ~^ image[6][14])} + {7'd0,(kernel[4][4] ~^ image[6][15])};
assign out_fmap[2][12][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][12])} + {7'd0,(kernel[0][1] ~^ image[2][13])} + {7'd0,(kernel[0][2] ~^ image[2][14])} + {7'd0,(kernel[0][3] ~^ image[2][15])} + {7'd0,(kernel[0][4] ~^ image[2][16])} + {7'd0,(kernel[1][0] ~^ image[3][12])} + {7'd0,(kernel[1][1] ~^ image[3][13])} + {7'd0,(kernel[1][2] ~^ image[3][14])} + {7'd0,(kernel[1][3] ~^ image[3][15])} + {7'd0,(kernel[1][4] ~^ image[3][16])} + {7'd0,(kernel[2][0] ~^ image[4][12])} + {7'd0,(kernel[2][1] ~^ image[4][13])} + {7'd0,(kernel[2][2] ~^ image[4][14])} + {7'd0,(kernel[2][3] ~^ image[4][15])} + {7'd0,(kernel[2][4] ~^ image[4][16])} + {7'd0,(kernel[3][0] ~^ image[5][12])} + {7'd0,(kernel[3][1] ~^ image[5][13])} + {7'd0,(kernel[3][2] ~^ image[5][14])} + {7'd0,(kernel[3][3] ~^ image[5][15])} + {7'd0,(kernel[3][4] ~^ image[5][16])} + {7'd0,(kernel[4][0] ~^ image[6][12])} + {7'd0,(kernel[4][1] ~^ image[6][13])} + {7'd0,(kernel[4][2] ~^ image[6][14])} + {7'd0,(kernel[4][3] ~^ image[6][15])} + {7'd0,(kernel[4][4] ~^ image[6][16])};
assign out_fmap[2][13][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][13])} + {7'd0,(kernel[0][1] ~^ image[2][14])} + {7'd0,(kernel[0][2] ~^ image[2][15])} + {7'd0,(kernel[0][3] ~^ image[2][16])} + {7'd0,(kernel[0][4] ~^ image[2][17])} + {7'd0,(kernel[1][0] ~^ image[3][13])} + {7'd0,(kernel[1][1] ~^ image[3][14])} + {7'd0,(kernel[1][2] ~^ image[3][15])} + {7'd0,(kernel[1][3] ~^ image[3][16])} + {7'd0,(kernel[1][4] ~^ image[3][17])} + {7'd0,(kernel[2][0] ~^ image[4][13])} + {7'd0,(kernel[2][1] ~^ image[4][14])} + {7'd0,(kernel[2][2] ~^ image[4][15])} + {7'd0,(kernel[2][3] ~^ image[4][16])} + {7'd0,(kernel[2][4] ~^ image[4][17])} + {7'd0,(kernel[3][0] ~^ image[5][13])} + {7'd0,(kernel[3][1] ~^ image[5][14])} + {7'd0,(kernel[3][2] ~^ image[5][15])} + {7'd0,(kernel[3][3] ~^ image[5][16])} + {7'd0,(kernel[3][4] ~^ image[5][17])} + {7'd0,(kernel[4][0] ~^ image[6][13])} + {7'd0,(kernel[4][1] ~^ image[6][14])} + {7'd0,(kernel[4][2] ~^ image[6][15])} + {7'd0,(kernel[4][3] ~^ image[6][16])} + {7'd0,(kernel[4][4] ~^ image[6][17])};
assign out_fmap[2][14][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][14])} + {7'd0,(kernel[0][1] ~^ image[2][15])} + {7'd0,(kernel[0][2] ~^ image[2][16])} + {7'd0,(kernel[0][3] ~^ image[2][17])} + {7'd0,(kernel[0][4] ~^ image[2][18])} + {7'd0,(kernel[1][0] ~^ image[3][14])} + {7'd0,(kernel[1][1] ~^ image[3][15])} + {7'd0,(kernel[1][2] ~^ image[3][16])} + {7'd0,(kernel[1][3] ~^ image[3][17])} + {7'd0,(kernel[1][4] ~^ image[3][18])} + {7'd0,(kernel[2][0] ~^ image[4][14])} + {7'd0,(kernel[2][1] ~^ image[4][15])} + {7'd0,(kernel[2][2] ~^ image[4][16])} + {7'd0,(kernel[2][3] ~^ image[4][17])} + {7'd0,(kernel[2][4] ~^ image[4][18])} + {7'd0,(kernel[3][0] ~^ image[5][14])} + {7'd0,(kernel[3][1] ~^ image[5][15])} + {7'd0,(kernel[3][2] ~^ image[5][16])} + {7'd0,(kernel[3][3] ~^ image[5][17])} + {7'd0,(kernel[3][4] ~^ image[5][18])} + {7'd0,(kernel[4][0] ~^ image[6][14])} + {7'd0,(kernel[4][1] ~^ image[6][15])} + {7'd0,(kernel[4][2] ~^ image[6][16])} + {7'd0,(kernel[4][3] ~^ image[6][17])} + {7'd0,(kernel[4][4] ~^ image[6][18])};
assign out_fmap[2][15][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][15])} + {7'd0,(kernel[0][1] ~^ image[2][16])} + {7'd0,(kernel[0][2] ~^ image[2][17])} + {7'd0,(kernel[0][3] ~^ image[2][18])} + {7'd0,(kernel[0][4] ~^ image[2][19])} + {7'd0,(kernel[1][0] ~^ image[3][15])} + {7'd0,(kernel[1][1] ~^ image[3][16])} + {7'd0,(kernel[1][2] ~^ image[3][17])} + {7'd0,(kernel[1][3] ~^ image[3][18])} + {7'd0,(kernel[1][4] ~^ image[3][19])} + {7'd0,(kernel[2][0] ~^ image[4][15])} + {7'd0,(kernel[2][1] ~^ image[4][16])} + {7'd0,(kernel[2][2] ~^ image[4][17])} + {7'd0,(kernel[2][3] ~^ image[4][18])} + {7'd0,(kernel[2][4] ~^ image[4][19])} + {7'd0,(kernel[3][0] ~^ image[5][15])} + {7'd0,(kernel[3][1] ~^ image[5][16])} + {7'd0,(kernel[3][2] ~^ image[5][17])} + {7'd0,(kernel[3][3] ~^ image[5][18])} + {7'd0,(kernel[3][4] ~^ image[5][19])} + {7'd0,(kernel[4][0] ~^ image[6][15])} + {7'd0,(kernel[4][1] ~^ image[6][16])} + {7'd0,(kernel[4][2] ~^ image[6][17])} + {7'd0,(kernel[4][3] ~^ image[6][18])} + {7'd0,(kernel[4][4] ~^ image[6][19])};
assign out_fmap[2][16][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][16])} + {7'd0,(kernel[0][1] ~^ image[2][17])} + {7'd0,(kernel[0][2] ~^ image[2][18])} + {7'd0,(kernel[0][3] ~^ image[2][19])} + {7'd0,(kernel[0][4] ~^ image[2][20])} + {7'd0,(kernel[1][0] ~^ image[3][16])} + {7'd0,(kernel[1][1] ~^ image[3][17])} + {7'd0,(kernel[1][2] ~^ image[3][18])} + {7'd0,(kernel[1][3] ~^ image[3][19])} + {7'd0,(kernel[1][4] ~^ image[3][20])} + {7'd0,(kernel[2][0] ~^ image[4][16])} + {7'd0,(kernel[2][1] ~^ image[4][17])} + {7'd0,(kernel[2][2] ~^ image[4][18])} + {7'd0,(kernel[2][3] ~^ image[4][19])} + {7'd0,(kernel[2][4] ~^ image[4][20])} + {7'd0,(kernel[3][0] ~^ image[5][16])} + {7'd0,(kernel[3][1] ~^ image[5][17])} + {7'd0,(kernel[3][2] ~^ image[5][18])} + {7'd0,(kernel[3][3] ~^ image[5][19])} + {7'd0,(kernel[3][4] ~^ image[5][20])} + {7'd0,(kernel[4][0] ~^ image[6][16])} + {7'd0,(kernel[4][1] ~^ image[6][17])} + {7'd0,(kernel[4][2] ~^ image[6][18])} + {7'd0,(kernel[4][3] ~^ image[6][19])} + {7'd0,(kernel[4][4] ~^ image[6][20])};
assign out_fmap[2][17][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][17])} + {7'd0,(kernel[0][1] ~^ image[2][18])} + {7'd0,(kernel[0][2] ~^ image[2][19])} + {7'd0,(kernel[0][3] ~^ image[2][20])} + {7'd0,(kernel[0][4] ~^ image[2][21])} + {7'd0,(kernel[1][0] ~^ image[3][17])} + {7'd0,(kernel[1][1] ~^ image[3][18])} + {7'd0,(kernel[1][2] ~^ image[3][19])} + {7'd0,(kernel[1][3] ~^ image[3][20])} + {7'd0,(kernel[1][4] ~^ image[3][21])} + {7'd0,(kernel[2][0] ~^ image[4][17])} + {7'd0,(kernel[2][1] ~^ image[4][18])} + {7'd0,(kernel[2][2] ~^ image[4][19])} + {7'd0,(kernel[2][3] ~^ image[4][20])} + {7'd0,(kernel[2][4] ~^ image[4][21])} + {7'd0,(kernel[3][0] ~^ image[5][17])} + {7'd0,(kernel[3][1] ~^ image[5][18])} + {7'd0,(kernel[3][2] ~^ image[5][19])} + {7'd0,(kernel[3][3] ~^ image[5][20])} + {7'd0,(kernel[3][4] ~^ image[5][21])} + {7'd0,(kernel[4][0] ~^ image[6][17])} + {7'd0,(kernel[4][1] ~^ image[6][18])} + {7'd0,(kernel[4][2] ~^ image[6][19])} + {7'd0,(kernel[4][3] ~^ image[6][20])} + {7'd0,(kernel[4][4] ~^ image[6][21])};
assign out_fmap[2][18][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][18])} + {7'd0,(kernel[0][1] ~^ image[2][19])} + {7'd0,(kernel[0][2] ~^ image[2][20])} + {7'd0,(kernel[0][3] ~^ image[2][21])} + {7'd0,(kernel[0][4] ~^ image[2][22])} + {7'd0,(kernel[1][0] ~^ image[3][18])} + {7'd0,(kernel[1][1] ~^ image[3][19])} + {7'd0,(kernel[1][2] ~^ image[3][20])} + {7'd0,(kernel[1][3] ~^ image[3][21])} + {7'd0,(kernel[1][4] ~^ image[3][22])} + {7'd0,(kernel[2][0] ~^ image[4][18])} + {7'd0,(kernel[2][1] ~^ image[4][19])} + {7'd0,(kernel[2][2] ~^ image[4][20])} + {7'd0,(kernel[2][3] ~^ image[4][21])} + {7'd0,(kernel[2][4] ~^ image[4][22])} + {7'd0,(kernel[3][0] ~^ image[5][18])} + {7'd0,(kernel[3][1] ~^ image[5][19])} + {7'd0,(kernel[3][2] ~^ image[5][20])} + {7'd0,(kernel[3][3] ~^ image[5][21])} + {7'd0,(kernel[3][4] ~^ image[5][22])} + {7'd0,(kernel[4][0] ~^ image[6][18])} + {7'd0,(kernel[4][1] ~^ image[6][19])} + {7'd0,(kernel[4][2] ~^ image[6][20])} + {7'd0,(kernel[4][3] ~^ image[6][21])} + {7'd0,(kernel[4][4] ~^ image[6][22])};
assign out_fmap[2][19][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][19])} + {7'd0,(kernel[0][1] ~^ image[2][20])} + {7'd0,(kernel[0][2] ~^ image[2][21])} + {7'd0,(kernel[0][3] ~^ image[2][22])} + {7'd0,(kernel[0][4] ~^ image[2][23])} + {7'd0,(kernel[1][0] ~^ image[3][19])} + {7'd0,(kernel[1][1] ~^ image[3][20])} + {7'd0,(kernel[1][2] ~^ image[3][21])} + {7'd0,(kernel[1][3] ~^ image[3][22])} + {7'd0,(kernel[1][4] ~^ image[3][23])} + {7'd0,(kernel[2][0] ~^ image[4][19])} + {7'd0,(kernel[2][1] ~^ image[4][20])} + {7'd0,(kernel[2][2] ~^ image[4][21])} + {7'd0,(kernel[2][3] ~^ image[4][22])} + {7'd0,(kernel[2][4] ~^ image[4][23])} + {7'd0,(kernel[3][0] ~^ image[5][19])} + {7'd0,(kernel[3][1] ~^ image[5][20])} + {7'd0,(kernel[3][2] ~^ image[5][21])} + {7'd0,(kernel[3][3] ~^ image[5][22])} + {7'd0,(kernel[3][4] ~^ image[5][23])} + {7'd0,(kernel[4][0] ~^ image[6][19])} + {7'd0,(kernel[4][1] ~^ image[6][20])} + {7'd0,(kernel[4][2] ~^ image[6][21])} + {7'd0,(kernel[4][3] ~^ image[6][22])} + {7'd0,(kernel[4][4] ~^ image[6][23])};
assign out_fmap[2][20][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][20])} + {7'd0,(kernel[0][1] ~^ image[2][21])} + {7'd0,(kernel[0][2] ~^ image[2][22])} + {7'd0,(kernel[0][3] ~^ image[2][23])} + {7'd0,(kernel[0][4] ~^ image[2][24])} + {7'd0,(kernel[1][0] ~^ image[3][20])} + {7'd0,(kernel[1][1] ~^ image[3][21])} + {7'd0,(kernel[1][2] ~^ image[3][22])} + {7'd0,(kernel[1][3] ~^ image[3][23])} + {7'd0,(kernel[1][4] ~^ image[3][24])} + {7'd0,(kernel[2][0] ~^ image[4][20])} + {7'd0,(kernel[2][1] ~^ image[4][21])} + {7'd0,(kernel[2][2] ~^ image[4][22])} + {7'd0,(kernel[2][3] ~^ image[4][23])} + {7'd0,(kernel[2][4] ~^ image[4][24])} + {7'd0,(kernel[3][0] ~^ image[5][20])} + {7'd0,(kernel[3][1] ~^ image[5][21])} + {7'd0,(kernel[3][2] ~^ image[5][22])} + {7'd0,(kernel[3][3] ~^ image[5][23])} + {7'd0,(kernel[3][4] ~^ image[5][24])} + {7'd0,(kernel[4][0] ~^ image[6][20])} + {7'd0,(kernel[4][1] ~^ image[6][21])} + {7'd0,(kernel[4][2] ~^ image[6][22])} + {7'd0,(kernel[4][3] ~^ image[6][23])} + {7'd0,(kernel[4][4] ~^ image[6][24])};
assign out_fmap[2][21][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][21])} + {7'd0,(kernel[0][1] ~^ image[2][22])} + {7'd0,(kernel[0][2] ~^ image[2][23])} + {7'd0,(kernel[0][3] ~^ image[2][24])} + {7'd0,(kernel[0][4] ~^ image[2][25])} + {7'd0,(kernel[1][0] ~^ image[3][21])} + {7'd0,(kernel[1][1] ~^ image[3][22])} + {7'd0,(kernel[1][2] ~^ image[3][23])} + {7'd0,(kernel[1][3] ~^ image[3][24])} + {7'd0,(kernel[1][4] ~^ image[3][25])} + {7'd0,(kernel[2][0] ~^ image[4][21])} + {7'd0,(kernel[2][1] ~^ image[4][22])} + {7'd0,(kernel[2][2] ~^ image[4][23])} + {7'd0,(kernel[2][3] ~^ image[4][24])} + {7'd0,(kernel[2][4] ~^ image[4][25])} + {7'd0,(kernel[3][0] ~^ image[5][21])} + {7'd0,(kernel[3][1] ~^ image[5][22])} + {7'd0,(kernel[3][2] ~^ image[5][23])} + {7'd0,(kernel[3][3] ~^ image[5][24])} + {7'd0,(kernel[3][4] ~^ image[5][25])} + {7'd0,(kernel[4][0] ~^ image[6][21])} + {7'd0,(kernel[4][1] ~^ image[6][22])} + {7'd0,(kernel[4][2] ~^ image[6][23])} + {7'd0,(kernel[4][3] ~^ image[6][24])} + {7'd0,(kernel[4][4] ~^ image[6][25])};
assign out_fmap[2][22][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][22])} + {7'd0,(kernel[0][1] ~^ image[2][23])} + {7'd0,(kernel[0][2] ~^ image[2][24])} + {7'd0,(kernel[0][3] ~^ image[2][25])} + {7'd0,(kernel[0][4] ~^ image[2][26])} + {7'd0,(kernel[1][0] ~^ image[3][22])} + {7'd0,(kernel[1][1] ~^ image[3][23])} + {7'd0,(kernel[1][2] ~^ image[3][24])} + {7'd0,(kernel[1][3] ~^ image[3][25])} + {7'd0,(kernel[1][4] ~^ image[3][26])} + {7'd0,(kernel[2][0] ~^ image[4][22])} + {7'd0,(kernel[2][1] ~^ image[4][23])} + {7'd0,(kernel[2][2] ~^ image[4][24])} + {7'd0,(kernel[2][3] ~^ image[4][25])} + {7'd0,(kernel[2][4] ~^ image[4][26])} + {7'd0,(kernel[3][0] ~^ image[5][22])} + {7'd0,(kernel[3][1] ~^ image[5][23])} + {7'd0,(kernel[3][2] ~^ image[5][24])} + {7'd0,(kernel[3][3] ~^ image[5][25])} + {7'd0,(kernel[3][4] ~^ image[5][26])} + {7'd0,(kernel[4][0] ~^ image[6][22])} + {7'd0,(kernel[4][1] ~^ image[6][23])} + {7'd0,(kernel[4][2] ~^ image[6][24])} + {7'd0,(kernel[4][3] ~^ image[6][25])} + {7'd0,(kernel[4][4] ~^ image[6][26])};
assign out_fmap[2][23][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[2][23])} + {7'd0,(kernel[0][1] ~^ image[2][24])} + {7'd0,(kernel[0][2] ~^ image[2][25])} + {7'd0,(kernel[0][3] ~^ image[2][26])} + {7'd0,(kernel[0][4] ~^ image[2][27])} + {7'd0,(kernel[1][0] ~^ image[3][23])} + {7'd0,(kernel[1][1] ~^ image[3][24])} + {7'd0,(kernel[1][2] ~^ image[3][25])} + {7'd0,(kernel[1][3] ~^ image[3][26])} + {7'd0,(kernel[1][4] ~^ image[3][27])} + {7'd0,(kernel[2][0] ~^ image[4][23])} + {7'd0,(kernel[2][1] ~^ image[4][24])} + {7'd0,(kernel[2][2] ~^ image[4][25])} + {7'd0,(kernel[2][3] ~^ image[4][26])} + {7'd0,(kernel[2][4] ~^ image[4][27])} + {7'd0,(kernel[3][0] ~^ image[5][23])} + {7'd0,(kernel[3][1] ~^ image[5][24])} + {7'd0,(kernel[3][2] ~^ image[5][25])} + {7'd0,(kernel[3][3] ~^ image[5][26])} + {7'd0,(kernel[3][4] ~^ image[5][27])} + {7'd0,(kernel[4][0] ~^ image[6][23])} + {7'd0,(kernel[4][1] ~^ image[6][24])} + {7'd0,(kernel[4][2] ~^ image[6][25])} + {7'd0,(kernel[4][3] ~^ image[6][26])} + {7'd0,(kernel[4][4] ~^ image[6][27])};
assign out_fmap[3][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][0])} + {7'd0,(kernel[0][1] ~^ image[3][1])} + {7'd0,(kernel[0][2] ~^ image[3][2])} + {7'd0,(kernel[0][3] ~^ image[3][3])} + {7'd0,(kernel[0][4] ~^ image[3][4])} + {7'd0,(kernel[1][0] ~^ image[4][0])} + {7'd0,(kernel[1][1] ~^ image[4][1])} + {7'd0,(kernel[1][2] ~^ image[4][2])} + {7'd0,(kernel[1][3] ~^ image[4][3])} + {7'd0,(kernel[1][4] ~^ image[4][4])} + {7'd0,(kernel[2][0] ~^ image[5][0])} + {7'd0,(kernel[2][1] ~^ image[5][1])} + {7'd0,(kernel[2][2] ~^ image[5][2])} + {7'd0,(kernel[2][3] ~^ image[5][3])} + {7'd0,(kernel[2][4] ~^ image[5][4])} + {7'd0,(kernel[3][0] ~^ image[6][0])} + {7'd0,(kernel[3][1] ~^ image[6][1])} + {7'd0,(kernel[3][2] ~^ image[6][2])} + {7'd0,(kernel[3][3] ~^ image[6][3])} + {7'd0,(kernel[3][4] ~^ image[6][4])} + {7'd0,(kernel[4][0] ~^ image[7][0])} + {7'd0,(kernel[4][1] ~^ image[7][1])} + {7'd0,(kernel[4][2] ~^ image[7][2])} + {7'd0,(kernel[4][3] ~^ image[7][3])} + {7'd0,(kernel[4][4] ~^ image[7][4])};
assign out_fmap[3][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][1])} + {7'd0,(kernel[0][1] ~^ image[3][2])} + {7'd0,(kernel[0][2] ~^ image[3][3])} + {7'd0,(kernel[0][3] ~^ image[3][4])} + {7'd0,(kernel[0][4] ~^ image[3][5])} + {7'd0,(kernel[1][0] ~^ image[4][1])} + {7'd0,(kernel[1][1] ~^ image[4][2])} + {7'd0,(kernel[1][2] ~^ image[4][3])} + {7'd0,(kernel[1][3] ~^ image[4][4])} + {7'd0,(kernel[1][4] ~^ image[4][5])} + {7'd0,(kernel[2][0] ~^ image[5][1])} + {7'd0,(kernel[2][1] ~^ image[5][2])} + {7'd0,(kernel[2][2] ~^ image[5][3])} + {7'd0,(kernel[2][3] ~^ image[5][4])} + {7'd0,(kernel[2][4] ~^ image[5][5])} + {7'd0,(kernel[3][0] ~^ image[6][1])} + {7'd0,(kernel[3][1] ~^ image[6][2])} + {7'd0,(kernel[3][2] ~^ image[6][3])} + {7'd0,(kernel[3][3] ~^ image[6][4])} + {7'd0,(kernel[3][4] ~^ image[6][5])} + {7'd0,(kernel[4][0] ~^ image[7][1])} + {7'd0,(kernel[4][1] ~^ image[7][2])} + {7'd0,(kernel[4][2] ~^ image[7][3])} + {7'd0,(kernel[4][3] ~^ image[7][4])} + {7'd0,(kernel[4][4] ~^ image[7][5])};
assign out_fmap[3][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][2])} + {7'd0,(kernel[0][1] ~^ image[3][3])} + {7'd0,(kernel[0][2] ~^ image[3][4])} + {7'd0,(kernel[0][3] ~^ image[3][5])} + {7'd0,(kernel[0][4] ~^ image[3][6])} + {7'd0,(kernel[1][0] ~^ image[4][2])} + {7'd0,(kernel[1][1] ~^ image[4][3])} + {7'd0,(kernel[1][2] ~^ image[4][4])} + {7'd0,(kernel[1][3] ~^ image[4][5])} + {7'd0,(kernel[1][4] ~^ image[4][6])} + {7'd0,(kernel[2][0] ~^ image[5][2])} + {7'd0,(kernel[2][1] ~^ image[5][3])} + {7'd0,(kernel[2][2] ~^ image[5][4])} + {7'd0,(kernel[2][3] ~^ image[5][5])} + {7'd0,(kernel[2][4] ~^ image[5][6])} + {7'd0,(kernel[3][0] ~^ image[6][2])} + {7'd0,(kernel[3][1] ~^ image[6][3])} + {7'd0,(kernel[3][2] ~^ image[6][4])} + {7'd0,(kernel[3][3] ~^ image[6][5])} + {7'd0,(kernel[3][4] ~^ image[6][6])} + {7'd0,(kernel[4][0] ~^ image[7][2])} + {7'd0,(kernel[4][1] ~^ image[7][3])} + {7'd0,(kernel[4][2] ~^ image[7][4])} + {7'd0,(kernel[4][3] ~^ image[7][5])} + {7'd0,(kernel[4][4] ~^ image[7][6])};
assign out_fmap[3][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][3])} + {7'd0,(kernel[0][1] ~^ image[3][4])} + {7'd0,(kernel[0][2] ~^ image[3][5])} + {7'd0,(kernel[0][3] ~^ image[3][6])} + {7'd0,(kernel[0][4] ~^ image[3][7])} + {7'd0,(kernel[1][0] ~^ image[4][3])} + {7'd0,(kernel[1][1] ~^ image[4][4])} + {7'd0,(kernel[1][2] ~^ image[4][5])} + {7'd0,(kernel[1][3] ~^ image[4][6])} + {7'd0,(kernel[1][4] ~^ image[4][7])} + {7'd0,(kernel[2][0] ~^ image[5][3])} + {7'd0,(kernel[2][1] ~^ image[5][4])} + {7'd0,(kernel[2][2] ~^ image[5][5])} + {7'd0,(kernel[2][3] ~^ image[5][6])} + {7'd0,(kernel[2][4] ~^ image[5][7])} + {7'd0,(kernel[3][0] ~^ image[6][3])} + {7'd0,(kernel[3][1] ~^ image[6][4])} + {7'd0,(kernel[3][2] ~^ image[6][5])} + {7'd0,(kernel[3][3] ~^ image[6][6])} + {7'd0,(kernel[3][4] ~^ image[6][7])} + {7'd0,(kernel[4][0] ~^ image[7][3])} + {7'd0,(kernel[4][1] ~^ image[7][4])} + {7'd0,(kernel[4][2] ~^ image[7][5])} + {7'd0,(kernel[4][3] ~^ image[7][6])} + {7'd0,(kernel[4][4] ~^ image[7][7])};
assign out_fmap[3][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][4])} + {7'd0,(kernel[0][1] ~^ image[3][5])} + {7'd0,(kernel[0][2] ~^ image[3][6])} + {7'd0,(kernel[0][3] ~^ image[3][7])} + {7'd0,(kernel[0][4] ~^ image[3][8])} + {7'd0,(kernel[1][0] ~^ image[4][4])} + {7'd0,(kernel[1][1] ~^ image[4][5])} + {7'd0,(kernel[1][2] ~^ image[4][6])} + {7'd0,(kernel[1][3] ~^ image[4][7])} + {7'd0,(kernel[1][4] ~^ image[4][8])} + {7'd0,(kernel[2][0] ~^ image[5][4])} + {7'd0,(kernel[2][1] ~^ image[5][5])} + {7'd0,(kernel[2][2] ~^ image[5][6])} + {7'd0,(kernel[2][3] ~^ image[5][7])} + {7'd0,(kernel[2][4] ~^ image[5][8])} + {7'd0,(kernel[3][0] ~^ image[6][4])} + {7'd0,(kernel[3][1] ~^ image[6][5])} + {7'd0,(kernel[3][2] ~^ image[6][6])} + {7'd0,(kernel[3][3] ~^ image[6][7])} + {7'd0,(kernel[3][4] ~^ image[6][8])} + {7'd0,(kernel[4][0] ~^ image[7][4])} + {7'd0,(kernel[4][1] ~^ image[7][5])} + {7'd0,(kernel[4][2] ~^ image[7][6])} + {7'd0,(kernel[4][3] ~^ image[7][7])} + {7'd0,(kernel[4][4] ~^ image[7][8])};
assign out_fmap[3][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][5])} + {7'd0,(kernel[0][1] ~^ image[3][6])} + {7'd0,(kernel[0][2] ~^ image[3][7])} + {7'd0,(kernel[0][3] ~^ image[3][8])} + {7'd0,(kernel[0][4] ~^ image[3][9])} + {7'd0,(kernel[1][0] ~^ image[4][5])} + {7'd0,(kernel[1][1] ~^ image[4][6])} + {7'd0,(kernel[1][2] ~^ image[4][7])} + {7'd0,(kernel[1][3] ~^ image[4][8])} + {7'd0,(kernel[1][4] ~^ image[4][9])} + {7'd0,(kernel[2][0] ~^ image[5][5])} + {7'd0,(kernel[2][1] ~^ image[5][6])} + {7'd0,(kernel[2][2] ~^ image[5][7])} + {7'd0,(kernel[2][3] ~^ image[5][8])} + {7'd0,(kernel[2][4] ~^ image[5][9])} + {7'd0,(kernel[3][0] ~^ image[6][5])} + {7'd0,(kernel[3][1] ~^ image[6][6])} + {7'd0,(kernel[3][2] ~^ image[6][7])} + {7'd0,(kernel[3][3] ~^ image[6][8])} + {7'd0,(kernel[3][4] ~^ image[6][9])} + {7'd0,(kernel[4][0] ~^ image[7][5])} + {7'd0,(kernel[4][1] ~^ image[7][6])} + {7'd0,(kernel[4][2] ~^ image[7][7])} + {7'd0,(kernel[4][3] ~^ image[7][8])} + {7'd0,(kernel[4][4] ~^ image[7][9])};
assign out_fmap[3][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][6])} + {7'd0,(kernel[0][1] ~^ image[3][7])} + {7'd0,(kernel[0][2] ~^ image[3][8])} + {7'd0,(kernel[0][3] ~^ image[3][9])} + {7'd0,(kernel[0][4] ~^ image[3][10])} + {7'd0,(kernel[1][0] ~^ image[4][6])} + {7'd0,(kernel[1][1] ~^ image[4][7])} + {7'd0,(kernel[1][2] ~^ image[4][8])} + {7'd0,(kernel[1][3] ~^ image[4][9])} + {7'd0,(kernel[1][4] ~^ image[4][10])} + {7'd0,(kernel[2][0] ~^ image[5][6])} + {7'd0,(kernel[2][1] ~^ image[5][7])} + {7'd0,(kernel[2][2] ~^ image[5][8])} + {7'd0,(kernel[2][3] ~^ image[5][9])} + {7'd0,(kernel[2][4] ~^ image[5][10])} + {7'd0,(kernel[3][0] ~^ image[6][6])} + {7'd0,(kernel[3][1] ~^ image[6][7])} + {7'd0,(kernel[3][2] ~^ image[6][8])} + {7'd0,(kernel[3][3] ~^ image[6][9])} + {7'd0,(kernel[3][4] ~^ image[6][10])} + {7'd0,(kernel[4][0] ~^ image[7][6])} + {7'd0,(kernel[4][1] ~^ image[7][7])} + {7'd0,(kernel[4][2] ~^ image[7][8])} + {7'd0,(kernel[4][3] ~^ image[7][9])} + {7'd0,(kernel[4][4] ~^ image[7][10])};
assign out_fmap[3][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][7])} + {7'd0,(kernel[0][1] ~^ image[3][8])} + {7'd0,(kernel[0][2] ~^ image[3][9])} + {7'd0,(kernel[0][3] ~^ image[3][10])} + {7'd0,(kernel[0][4] ~^ image[3][11])} + {7'd0,(kernel[1][0] ~^ image[4][7])} + {7'd0,(kernel[1][1] ~^ image[4][8])} + {7'd0,(kernel[1][2] ~^ image[4][9])} + {7'd0,(kernel[1][3] ~^ image[4][10])} + {7'd0,(kernel[1][4] ~^ image[4][11])} + {7'd0,(kernel[2][0] ~^ image[5][7])} + {7'd0,(kernel[2][1] ~^ image[5][8])} + {7'd0,(kernel[2][2] ~^ image[5][9])} + {7'd0,(kernel[2][3] ~^ image[5][10])} + {7'd0,(kernel[2][4] ~^ image[5][11])} + {7'd0,(kernel[3][0] ~^ image[6][7])} + {7'd0,(kernel[3][1] ~^ image[6][8])} + {7'd0,(kernel[3][2] ~^ image[6][9])} + {7'd0,(kernel[3][3] ~^ image[6][10])} + {7'd0,(kernel[3][4] ~^ image[6][11])} + {7'd0,(kernel[4][0] ~^ image[7][7])} + {7'd0,(kernel[4][1] ~^ image[7][8])} + {7'd0,(kernel[4][2] ~^ image[7][9])} + {7'd0,(kernel[4][3] ~^ image[7][10])} + {7'd0,(kernel[4][4] ~^ image[7][11])};
assign out_fmap[3][8][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][8])} + {7'd0,(kernel[0][1] ~^ image[3][9])} + {7'd0,(kernel[0][2] ~^ image[3][10])} + {7'd0,(kernel[0][3] ~^ image[3][11])} + {7'd0,(kernel[0][4] ~^ image[3][12])} + {7'd0,(kernel[1][0] ~^ image[4][8])} + {7'd0,(kernel[1][1] ~^ image[4][9])} + {7'd0,(kernel[1][2] ~^ image[4][10])} + {7'd0,(kernel[1][3] ~^ image[4][11])} + {7'd0,(kernel[1][4] ~^ image[4][12])} + {7'd0,(kernel[2][0] ~^ image[5][8])} + {7'd0,(kernel[2][1] ~^ image[5][9])} + {7'd0,(kernel[2][2] ~^ image[5][10])} + {7'd0,(kernel[2][3] ~^ image[5][11])} + {7'd0,(kernel[2][4] ~^ image[5][12])} + {7'd0,(kernel[3][0] ~^ image[6][8])} + {7'd0,(kernel[3][1] ~^ image[6][9])} + {7'd0,(kernel[3][2] ~^ image[6][10])} + {7'd0,(kernel[3][3] ~^ image[6][11])} + {7'd0,(kernel[3][4] ~^ image[6][12])} + {7'd0,(kernel[4][0] ~^ image[7][8])} + {7'd0,(kernel[4][1] ~^ image[7][9])} + {7'd0,(kernel[4][2] ~^ image[7][10])} + {7'd0,(kernel[4][3] ~^ image[7][11])} + {7'd0,(kernel[4][4] ~^ image[7][12])};
assign out_fmap[3][9][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][9])} + {7'd0,(kernel[0][1] ~^ image[3][10])} + {7'd0,(kernel[0][2] ~^ image[3][11])} + {7'd0,(kernel[0][3] ~^ image[3][12])} + {7'd0,(kernel[0][4] ~^ image[3][13])} + {7'd0,(kernel[1][0] ~^ image[4][9])} + {7'd0,(kernel[1][1] ~^ image[4][10])} + {7'd0,(kernel[1][2] ~^ image[4][11])} + {7'd0,(kernel[1][3] ~^ image[4][12])} + {7'd0,(kernel[1][4] ~^ image[4][13])} + {7'd0,(kernel[2][0] ~^ image[5][9])} + {7'd0,(kernel[2][1] ~^ image[5][10])} + {7'd0,(kernel[2][2] ~^ image[5][11])} + {7'd0,(kernel[2][3] ~^ image[5][12])} + {7'd0,(kernel[2][4] ~^ image[5][13])} + {7'd0,(kernel[3][0] ~^ image[6][9])} + {7'd0,(kernel[3][1] ~^ image[6][10])} + {7'd0,(kernel[3][2] ~^ image[6][11])} + {7'd0,(kernel[3][3] ~^ image[6][12])} + {7'd0,(kernel[3][4] ~^ image[6][13])} + {7'd0,(kernel[4][0] ~^ image[7][9])} + {7'd0,(kernel[4][1] ~^ image[7][10])} + {7'd0,(kernel[4][2] ~^ image[7][11])} + {7'd0,(kernel[4][3] ~^ image[7][12])} + {7'd0,(kernel[4][4] ~^ image[7][13])};
assign out_fmap[3][10][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][10])} + {7'd0,(kernel[0][1] ~^ image[3][11])} + {7'd0,(kernel[0][2] ~^ image[3][12])} + {7'd0,(kernel[0][3] ~^ image[3][13])} + {7'd0,(kernel[0][4] ~^ image[3][14])} + {7'd0,(kernel[1][0] ~^ image[4][10])} + {7'd0,(kernel[1][1] ~^ image[4][11])} + {7'd0,(kernel[1][2] ~^ image[4][12])} + {7'd0,(kernel[1][3] ~^ image[4][13])} + {7'd0,(kernel[1][4] ~^ image[4][14])} + {7'd0,(kernel[2][0] ~^ image[5][10])} + {7'd0,(kernel[2][1] ~^ image[5][11])} + {7'd0,(kernel[2][2] ~^ image[5][12])} + {7'd0,(kernel[2][3] ~^ image[5][13])} + {7'd0,(kernel[2][4] ~^ image[5][14])} + {7'd0,(kernel[3][0] ~^ image[6][10])} + {7'd0,(kernel[3][1] ~^ image[6][11])} + {7'd0,(kernel[3][2] ~^ image[6][12])} + {7'd0,(kernel[3][3] ~^ image[6][13])} + {7'd0,(kernel[3][4] ~^ image[6][14])} + {7'd0,(kernel[4][0] ~^ image[7][10])} + {7'd0,(kernel[4][1] ~^ image[7][11])} + {7'd0,(kernel[4][2] ~^ image[7][12])} + {7'd0,(kernel[4][3] ~^ image[7][13])} + {7'd0,(kernel[4][4] ~^ image[7][14])};
assign out_fmap[3][11][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][11])} + {7'd0,(kernel[0][1] ~^ image[3][12])} + {7'd0,(kernel[0][2] ~^ image[3][13])} + {7'd0,(kernel[0][3] ~^ image[3][14])} + {7'd0,(kernel[0][4] ~^ image[3][15])} + {7'd0,(kernel[1][0] ~^ image[4][11])} + {7'd0,(kernel[1][1] ~^ image[4][12])} + {7'd0,(kernel[1][2] ~^ image[4][13])} + {7'd0,(kernel[1][3] ~^ image[4][14])} + {7'd0,(kernel[1][4] ~^ image[4][15])} + {7'd0,(kernel[2][0] ~^ image[5][11])} + {7'd0,(kernel[2][1] ~^ image[5][12])} + {7'd0,(kernel[2][2] ~^ image[5][13])} + {7'd0,(kernel[2][3] ~^ image[5][14])} + {7'd0,(kernel[2][4] ~^ image[5][15])} + {7'd0,(kernel[3][0] ~^ image[6][11])} + {7'd0,(kernel[3][1] ~^ image[6][12])} + {7'd0,(kernel[3][2] ~^ image[6][13])} + {7'd0,(kernel[3][3] ~^ image[6][14])} + {7'd0,(kernel[3][4] ~^ image[6][15])} + {7'd0,(kernel[4][0] ~^ image[7][11])} + {7'd0,(kernel[4][1] ~^ image[7][12])} + {7'd0,(kernel[4][2] ~^ image[7][13])} + {7'd0,(kernel[4][3] ~^ image[7][14])} + {7'd0,(kernel[4][4] ~^ image[7][15])};
assign out_fmap[3][12][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][12])} + {7'd0,(kernel[0][1] ~^ image[3][13])} + {7'd0,(kernel[0][2] ~^ image[3][14])} + {7'd0,(kernel[0][3] ~^ image[3][15])} + {7'd0,(kernel[0][4] ~^ image[3][16])} + {7'd0,(kernel[1][0] ~^ image[4][12])} + {7'd0,(kernel[1][1] ~^ image[4][13])} + {7'd0,(kernel[1][2] ~^ image[4][14])} + {7'd0,(kernel[1][3] ~^ image[4][15])} + {7'd0,(kernel[1][4] ~^ image[4][16])} + {7'd0,(kernel[2][0] ~^ image[5][12])} + {7'd0,(kernel[2][1] ~^ image[5][13])} + {7'd0,(kernel[2][2] ~^ image[5][14])} + {7'd0,(kernel[2][3] ~^ image[5][15])} + {7'd0,(kernel[2][4] ~^ image[5][16])} + {7'd0,(kernel[3][0] ~^ image[6][12])} + {7'd0,(kernel[3][1] ~^ image[6][13])} + {7'd0,(kernel[3][2] ~^ image[6][14])} + {7'd0,(kernel[3][3] ~^ image[6][15])} + {7'd0,(kernel[3][4] ~^ image[6][16])} + {7'd0,(kernel[4][0] ~^ image[7][12])} + {7'd0,(kernel[4][1] ~^ image[7][13])} + {7'd0,(kernel[4][2] ~^ image[7][14])} + {7'd0,(kernel[4][3] ~^ image[7][15])} + {7'd0,(kernel[4][4] ~^ image[7][16])};
assign out_fmap[3][13][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][13])} + {7'd0,(kernel[0][1] ~^ image[3][14])} + {7'd0,(kernel[0][2] ~^ image[3][15])} + {7'd0,(kernel[0][3] ~^ image[3][16])} + {7'd0,(kernel[0][4] ~^ image[3][17])} + {7'd0,(kernel[1][0] ~^ image[4][13])} + {7'd0,(kernel[1][1] ~^ image[4][14])} + {7'd0,(kernel[1][2] ~^ image[4][15])} + {7'd0,(kernel[1][3] ~^ image[4][16])} + {7'd0,(kernel[1][4] ~^ image[4][17])} + {7'd0,(kernel[2][0] ~^ image[5][13])} + {7'd0,(kernel[2][1] ~^ image[5][14])} + {7'd0,(kernel[2][2] ~^ image[5][15])} + {7'd0,(kernel[2][3] ~^ image[5][16])} + {7'd0,(kernel[2][4] ~^ image[5][17])} + {7'd0,(kernel[3][0] ~^ image[6][13])} + {7'd0,(kernel[3][1] ~^ image[6][14])} + {7'd0,(kernel[3][2] ~^ image[6][15])} + {7'd0,(kernel[3][3] ~^ image[6][16])} + {7'd0,(kernel[3][4] ~^ image[6][17])} + {7'd0,(kernel[4][0] ~^ image[7][13])} + {7'd0,(kernel[4][1] ~^ image[7][14])} + {7'd0,(kernel[4][2] ~^ image[7][15])} + {7'd0,(kernel[4][3] ~^ image[7][16])} + {7'd0,(kernel[4][4] ~^ image[7][17])};
assign out_fmap[3][14][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][14])} + {7'd0,(kernel[0][1] ~^ image[3][15])} + {7'd0,(kernel[0][2] ~^ image[3][16])} + {7'd0,(kernel[0][3] ~^ image[3][17])} + {7'd0,(kernel[0][4] ~^ image[3][18])} + {7'd0,(kernel[1][0] ~^ image[4][14])} + {7'd0,(kernel[1][1] ~^ image[4][15])} + {7'd0,(kernel[1][2] ~^ image[4][16])} + {7'd0,(kernel[1][3] ~^ image[4][17])} + {7'd0,(kernel[1][4] ~^ image[4][18])} + {7'd0,(kernel[2][0] ~^ image[5][14])} + {7'd0,(kernel[2][1] ~^ image[5][15])} + {7'd0,(kernel[2][2] ~^ image[5][16])} + {7'd0,(kernel[2][3] ~^ image[5][17])} + {7'd0,(kernel[2][4] ~^ image[5][18])} + {7'd0,(kernel[3][0] ~^ image[6][14])} + {7'd0,(kernel[3][1] ~^ image[6][15])} + {7'd0,(kernel[3][2] ~^ image[6][16])} + {7'd0,(kernel[3][3] ~^ image[6][17])} + {7'd0,(kernel[3][4] ~^ image[6][18])} + {7'd0,(kernel[4][0] ~^ image[7][14])} + {7'd0,(kernel[4][1] ~^ image[7][15])} + {7'd0,(kernel[4][2] ~^ image[7][16])} + {7'd0,(kernel[4][3] ~^ image[7][17])} + {7'd0,(kernel[4][4] ~^ image[7][18])};
assign out_fmap[3][15][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][15])} + {7'd0,(kernel[0][1] ~^ image[3][16])} + {7'd0,(kernel[0][2] ~^ image[3][17])} + {7'd0,(kernel[0][3] ~^ image[3][18])} + {7'd0,(kernel[0][4] ~^ image[3][19])} + {7'd0,(kernel[1][0] ~^ image[4][15])} + {7'd0,(kernel[1][1] ~^ image[4][16])} + {7'd0,(kernel[1][2] ~^ image[4][17])} + {7'd0,(kernel[1][3] ~^ image[4][18])} + {7'd0,(kernel[1][4] ~^ image[4][19])} + {7'd0,(kernel[2][0] ~^ image[5][15])} + {7'd0,(kernel[2][1] ~^ image[5][16])} + {7'd0,(kernel[2][2] ~^ image[5][17])} + {7'd0,(kernel[2][3] ~^ image[5][18])} + {7'd0,(kernel[2][4] ~^ image[5][19])} + {7'd0,(kernel[3][0] ~^ image[6][15])} + {7'd0,(kernel[3][1] ~^ image[6][16])} + {7'd0,(kernel[3][2] ~^ image[6][17])} + {7'd0,(kernel[3][3] ~^ image[6][18])} + {7'd0,(kernel[3][4] ~^ image[6][19])} + {7'd0,(kernel[4][0] ~^ image[7][15])} + {7'd0,(kernel[4][1] ~^ image[7][16])} + {7'd0,(kernel[4][2] ~^ image[7][17])} + {7'd0,(kernel[4][3] ~^ image[7][18])} + {7'd0,(kernel[4][4] ~^ image[7][19])};
assign out_fmap[3][16][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][16])} + {7'd0,(kernel[0][1] ~^ image[3][17])} + {7'd0,(kernel[0][2] ~^ image[3][18])} + {7'd0,(kernel[0][3] ~^ image[3][19])} + {7'd0,(kernel[0][4] ~^ image[3][20])} + {7'd0,(kernel[1][0] ~^ image[4][16])} + {7'd0,(kernel[1][1] ~^ image[4][17])} + {7'd0,(kernel[1][2] ~^ image[4][18])} + {7'd0,(kernel[1][3] ~^ image[4][19])} + {7'd0,(kernel[1][4] ~^ image[4][20])} + {7'd0,(kernel[2][0] ~^ image[5][16])} + {7'd0,(kernel[2][1] ~^ image[5][17])} + {7'd0,(kernel[2][2] ~^ image[5][18])} + {7'd0,(kernel[2][3] ~^ image[5][19])} + {7'd0,(kernel[2][4] ~^ image[5][20])} + {7'd0,(kernel[3][0] ~^ image[6][16])} + {7'd0,(kernel[3][1] ~^ image[6][17])} + {7'd0,(kernel[3][2] ~^ image[6][18])} + {7'd0,(kernel[3][3] ~^ image[6][19])} + {7'd0,(kernel[3][4] ~^ image[6][20])} + {7'd0,(kernel[4][0] ~^ image[7][16])} + {7'd0,(kernel[4][1] ~^ image[7][17])} + {7'd0,(kernel[4][2] ~^ image[7][18])} + {7'd0,(kernel[4][3] ~^ image[7][19])} + {7'd0,(kernel[4][4] ~^ image[7][20])};
assign out_fmap[3][17][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][17])} + {7'd0,(kernel[0][1] ~^ image[3][18])} + {7'd0,(kernel[0][2] ~^ image[3][19])} + {7'd0,(kernel[0][3] ~^ image[3][20])} + {7'd0,(kernel[0][4] ~^ image[3][21])} + {7'd0,(kernel[1][0] ~^ image[4][17])} + {7'd0,(kernel[1][1] ~^ image[4][18])} + {7'd0,(kernel[1][2] ~^ image[4][19])} + {7'd0,(kernel[1][3] ~^ image[4][20])} + {7'd0,(kernel[1][4] ~^ image[4][21])} + {7'd0,(kernel[2][0] ~^ image[5][17])} + {7'd0,(kernel[2][1] ~^ image[5][18])} + {7'd0,(kernel[2][2] ~^ image[5][19])} + {7'd0,(kernel[2][3] ~^ image[5][20])} + {7'd0,(kernel[2][4] ~^ image[5][21])} + {7'd0,(kernel[3][0] ~^ image[6][17])} + {7'd0,(kernel[3][1] ~^ image[6][18])} + {7'd0,(kernel[3][2] ~^ image[6][19])} + {7'd0,(kernel[3][3] ~^ image[6][20])} + {7'd0,(kernel[3][4] ~^ image[6][21])} + {7'd0,(kernel[4][0] ~^ image[7][17])} + {7'd0,(kernel[4][1] ~^ image[7][18])} + {7'd0,(kernel[4][2] ~^ image[7][19])} + {7'd0,(kernel[4][3] ~^ image[7][20])} + {7'd0,(kernel[4][4] ~^ image[7][21])};
assign out_fmap[3][18][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][18])} + {7'd0,(kernel[0][1] ~^ image[3][19])} + {7'd0,(kernel[0][2] ~^ image[3][20])} + {7'd0,(kernel[0][3] ~^ image[3][21])} + {7'd0,(kernel[0][4] ~^ image[3][22])} + {7'd0,(kernel[1][0] ~^ image[4][18])} + {7'd0,(kernel[1][1] ~^ image[4][19])} + {7'd0,(kernel[1][2] ~^ image[4][20])} + {7'd0,(kernel[1][3] ~^ image[4][21])} + {7'd0,(kernel[1][4] ~^ image[4][22])} + {7'd0,(kernel[2][0] ~^ image[5][18])} + {7'd0,(kernel[2][1] ~^ image[5][19])} + {7'd0,(kernel[2][2] ~^ image[5][20])} + {7'd0,(kernel[2][3] ~^ image[5][21])} + {7'd0,(kernel[2][4] ~^ image[5][22])} + {7'd0,(kernel[3][0] ~^ image[6][18])} + {7'd0,(kernel[3][1] ~^ image[6][19])} + {7'd0,(kernel[3][2] ~^ image[6][20])} + {7'd0,(kernel[3][3] ~^ image[6][21])} + {7'd0,(kernel[3][4] ~^ image[6][22])} + {7'd0,(kernel[4][0] ~^ image[7][18])} + {7'd0,(kernel[4][1] ~^ image[7][19])} + {7'd0,(kernel[4][2] ~^ image[7][20])} + {7'd0,(kernel[4][3] ~^ image[7][21])} + {7'd0,(kernel[4][4] ~^ image[7][22])};
assign out_fmap[3][19][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][19])} + {7'd0,(kernel[0][1] ~^ image[3][20])} + {7'd0,(kernel[0][2] ~^ image[3][21])} + {7'd0,(kernel[0][3] ~^ image[3][22])} + {7'd0,(kernel[0][4] ~^ image[3][23])} + {7'd0,(kernel[1][0] ~^ image[4][19])} + {7'd0,(kernel[1][1] ~^ image[4][20])} + {7'd0,(kernel[1][2] ~^ image[4][21])} + {7'd0,(kernel[1][3] ~^ image[4][22])} + {7'd0,(kernel[1][4] ~^ image[4][23])} + {7'd0,(kernel[2][0] ~^ image[5][19])} + {7'd0,(kernel[2][1] ~^ image[5][20])} + {7'd0,(kernel[2][2] ~^ image[5][21])} + {7'd0,(kernel[2][3] ~^ image[5][22])} + {7'd0,(kernel[2][4] ~^ image[5][23])} + {7'd0,(kernel[3][0] ~^ image[6][19])} + {7'd0,(kernel[3][1] ~^ image[6][20])} + {7'd0,(kernel[3][2] ~^ image[6][21])} + {7'd0,(kernel[3][3] ~^ image[6][22])} + {7'd0,(kernel[3][4] ~^ image[6][23])} + {7'd0,(kernel[4][0] ~^ image[7][19])} + {7'd0,(kernel[4][1] ~^ image[7][20])} + {7'd0,(kernel[4][2] ~^ image[7][21])} + {7'd0,(kernel[4][3] ~^ image[7][22])} + {7'd0,(kernel[4][4] ~^ image[7][23])};
assign out_fmap[3][20][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][20])} + {7'd0,(kernel[0][1] ~^ image[3][21])} + {7'd0,(kernel[0][2] ~^ image[3][22])} + {7'd0,(kernel[0][3] ~^ image[3][23])} + {7'd0,(kernel[0][4] ~^ image[3][24])} + {7'd0,(kernel[1][0] ~^ image[4][20])} + {7'd0,(kernel[1][1] ~^ image[4][21])} + {7'd0,(kernel[1][2] ~^ image[4][22])} + {7'd0,(kernel[1][3] ~^ image[4][23])} + {7'd0,(kernel[1][4] ~^ image[4][24])} + {7'd0,(kernel[2][0] ~^ image[5][20])} + {7'd0,(kernel[2][1] ~^ image[5][21])} + {7'd0,(kernel[2][2] ~^ image[5][22])} + {7'd0,(kernel[2][3] ~^ image[5][23])} + {7'd0,(kernel[2][4] ~^ image[5][24])} + {7'd0,(kernel[3][0] ~^ image[6][20])} + {7'd0,(kernel[3][1] ~^ image[6][21])} + {7'd0,(kernel[3][2] ~^ image[6][22])} + {7'd0,(kernel[3][3] ~^ image[6][23])} + {7'd0,(kernel[3][4] ~^ image[6][24])} + {7'd0,(kernel[4][0] ~^ image[7][20])} + {7'd0,(kernel[4][1] ~^ image[7][21])} + {7'd0,(kernel[4][2] ~^ image[7][22])} + {7'd0,(kernel[4][3] ~^ image[7][23])} + {7'd0,(kernel[4][4] ~^ image[7][24])};
assign out_fmap[3][21][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][21])} + {7'd0,(kernel[0][1] ~^ image[3][22])} + {7'd0,(kernel[0][2] ~^ image[3][23])} + {7'd0,(kernel[0][3] ~^ image[3][24])} + {7'd0,(kernel[0][4] ~^ image[3][25])} + {7'd0,(kernel[1][0] ~^ image[4][21])} + {7'd0,(kernel[1][1] ~^ image[4][22])} + {7'd0,(kernel[1][2] ~^ image[4][23])} + {7'd0,(kernel[1][3] ~^ image[4][24])} + {7'd0,(kernel[1][4] ~^ image[4][25])} + {7'd0,(kernel[2][0] ~^ image[5][21])} + {7'd0,(kernel[2][1] ~^ image[5][22])} + {7'd0,(kernel[2][2] ~^ image[5][23])} + {7'd0,(kernel[2][3] ~^ image[5][24])} + {7'd0,(kernel[2][4] ~^ image[5][25])} + {7'd0,(kernel[3][0] ~^ image[6][21])} + {7'd0,(kernel[3][1] ~^ image[6][22])} + {7'd0,(kernel[3][2] ~^ image[6][23])} + {7'd0,(kernel[3][3] ~^ image[6][24])} + {7'd0,(kernel[3][4] ~^ image[6][25])} + {7'd0,(kernel[4][0] ~^ image[7][21])} + {7'd0,(kernel[4][1] ~^ image[7][22])} + {7'd0,(kernel[4][2] ~^ image[7][23])} + {7'd0,(kernel[4][3] ~^ image[7][24])} + {7'd0,(kernel[4][4] ~^ image[7][25])};
assign out_fmap[3][22][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][22])} + {7'd0,(kernel[0][1] ~^ image[3][23])} + {7'd0,(kernel[0][2] ~^ image[3][24])} + {7'd0,(kernel[0][3] ~^ image[3][25])} + {7'd0,(kernel[0][4] ~^ image[3][26])} + {7'd0,(kernel[1][0] ~^ image[4][22])} + {7'd0,(kernel[1][1] ~^ image[4][23])} + {7'd0,(kernel[1][2] ~^ image[4][24])} + {7'd0,(kernel[1][3] ~^ image[4][25])} + {7'd0,(kernel[1][4] ~^ image[4][26])} + {7'd0,(kernel[2][0] ~^ image[5][22])} + {7'd0,(kernel[2][1] ~^ image[5][23])} + {7'd0,(kernel[2][2] ~^ image[5][24])} + {7'd0,(kernel[2][3] ~^ image[5][25])} + {7'd0,(kernel[2][4] ~^ image[5][26])} + {7'd0,(kernel[3][0] ~^ image[6][22])} + {7'd0,(kernel[3][1] ~^ image[6][23])} + {7'd0,(kernel[3][2] ~^ image[6][24])} + {7'd0,(kernel[3][3] ~^ image[6][25])} + {7'd0,(kernel[3][4] ~^ image[6][26])} + {7'd0,(kernel[4][0] ~^ image[7][22])} + {7'd0,(kernel[4][1] ~^ image[7][23])} + {7'd0,(kernel[4][2] ~^ image[7][24])} + {7'd0,(kernel[4][3] ~^ image[7][25])} + {7'd0,(kernel[4][4] ~^ image[7][26])};
assign out_fmap[3][23][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[3][23])} + {7'd0,(kernel[0][1] ~^ image[3][24])} + {7'd0,(kernel[0][2] ~^ image[3][25])} + {7'd0,(kernel[0][3] ~^ image[3][26])} + {7'd0,(kernel[0][4] ~^ image[3][27])} + {7'd0,(kernel[1][0] ~^ image[4][23])} + {7'd0,(kernel[1][1] ~^ image[4][24])} + {7'd0,(kernel[1][2] ~^ image[4][25])} + {7'd0,(kernel[1][3] ~^ image[4][26])} + {7'd0,(kernel[1][4] ~^ image[4][27])} + {7'd0,(kernel[2][0] ~^ image[5][23])} + {7'd0,(kernel[2][1] ~^ image[5][24])} + {7'd0,(kernel[2][2] ~^ image[5][25])} + {7'd0,(kernel[2][3] ~^ image[5][26])} + {7'd0,(kernel[2][4] ~^ image[5][27])} + {7'd0,(kernel[3][0] ~^ image[6][23])} + {7'd0,(kernel[3][1] ~^ image[6][24])} + {7'd0,(kernel[3][2] ~^ image[6][25])} + {7'd0,(kernel[3][3] ~^ image[6][26])} + {7'd0,(kernel[3][4] ~^ image[6][27])} + {7'd0,(kernel[4][0] ~^ image[7][23])} + {7'd0,(kernel[4][1] ~^ image[7][24])} + {7'd0,(kernel[4][2] ~^ image[7][25])} + {7'd0,(kernel[4][3] ~^ image[7][26])} + {7'd0,(kernel[4][4] ~^ image[7][27])};
assign out_fmap[4][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][0])} + {7'd0,(kernel[0][1] ~^ image[4][1])} + {7'd0,(kernel[0][2] ~^ image[4][2])} + {7'd0,(kernel[0][3] ~^ image[4][3])} + {7'd0,(kernel[0][4] ~^ image[4][4])} + {7'd0,(kernel[1][0] ~^ image[5][0])} + {7'd0,(kernel[1][1] ~^ image[5][1])} + {7'd0,(kernel[1][2] ~^ image[5][2])} + {7'd0,(kernel[1][3] ~^ image[5][3])} + {7'd0,(kernel[1][4] ~^ image[5][4])} + {7'd0,(kernel[2][0] ~^ image[6][0])} + {7'd0,(kernel[2][1] ~^ image[6][1])} + {7'd0,(kernel[2][2] ~^ image[6][2])} + {7'd0,(kernel[2][3] ~^ image[6][3])} + {7'd0,(kernel[2][4] ~^ image[6][4])} + {7'd0,(kernel[3][0] ~^ image[7][0])} + {7'd0,(kernel[3][1] ~^ image[7][1])} + {7'd0,(kernel[3][2] ~^ image[7][2])} + {7'd0,(kernel[3][3] ~^ image[7][3])} + {7'd0,(kernel[3][4] ~^ image[7][4])} + {7'd0,(kernel[4][0] ~^ image[8][0])} + {7'd0,(kernel[4][1] ~^ image[8][1])} + {7'd0,(kernel[4][2] ~^ image[8][2])} + {7'd0,(kernel[4][3] ~^ image[8][3])} + {7'd0,(kernel[4][4] ~^ image[8][4])};
assign out_fmap[4][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][1])} + {7'd0,(kernel[0][1] ~^ image[4][2])} + {7'd0,(kernel[0][2] ~^ image[4][3])} + {7'd0,(kernel[0][3] ~^ image[4][4])} + {7'd0,(kernel[0][4] ~^ image[4][5])} + {7'd0,(kernel[1][0] ~^ image[5][1])} + {7'd0,(kernel[1][1] ~^ image[5][2])} + {7'd0,(kernel[1][2] ~^ image[5][3])} + {7'd0,(kernel[1][3] ~^ image[5][4])} + {7'd0,(kernel[1][4] ~^ image[5][5])} + {7'd0,(kernel[2][0] ~^ image[6][1])} + {7'd0,(kernel[2][1] ~^ image[6][2])} + {7'd0,(kernel[2][2] ~^ image[6][3])} + {7'd0,(kernel[2][3] ~^ image[6][4])} + {7'd0,(kernel[2][4] ~^ image[6][5])} + {7'd0,(kernel[3][0] ~^ image[7][1])} + {7'd0,(kernel[3][1] ~^ image[7][2])} + {7'd0,(kernel[3][2] ~^ image[7][3])} + {7'd0,(kernel[3][3] ~^ image[7][4])} + {7'd0,(kernel[3][4] ~^ image[7][5])} + {7'd0,(kernel[4][0] ~^ image[8][1])} + {7'd0,(kernel[4][1] ~^ image[8][2])} + {7'd0,(kernel[4][2] ~^ image[8][3])} + {7'd0,(kernel[4][3] ~^ image[8][4])} + {7'd0,(kernel[4][4] ~^ image[8][5])};
assign out_fmap[4][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][2])} + {7'd0,(kernel[0][1] ~^ image[4][3])} + {7'd0,(kernel[0][2] ~^ image[4][4])} + {7'd0,(kernel[0][3] ~^ image[4][5])} + {7'd0,(kernel[0][4] ~^ image[4][6])} + {7'd0,(kernel[1][0] ~^ image[5][2])} + {7'd0,(kernel[1][1] ~^ image[5][3])} + {7'd0,(kernel[1][2] ~^ image[5][4])} + {7'd0,(kernel[1][3] ~^ image[5][5])} + {7'd0,(kernel[1][4] ~^ image[5][6])} + {7'd0,(kernel[2][0] ~^ image[6][2])} + {7'd0,(kernel[2][1] ~^ image[6][3])} + {7'd0,(kernel[2][2] ~^ image[6][4])} + {7'd0,(kernel[2][3] ~^ image[6][5])} + {7'd0,(kernel[2][4] ~^ image[6][6])} + {7'd0,(kernel[3][0] ~^ image[7][2])} + {7'd0,(kernel[3][1] ~^ image[7][3])} + {7'd0,(kernel[3][2] ~^ image[7][4])} + {7'd0,(kernel[3][3] ~^ image[7][5])} + {7'd0,(kernel[3][4] ~^ image[7][6])} + {7'd0,(kernel[4][0] ~^ image[8][2])} + {7'd0,(kernel[4][1] ~^ image[8][3])} + {7'd0,(kernel[4][2] ~^ image[8][4])} + {7'd0,(kernel[4][3] ~^ image[8][5])} + {7'd0,(kernel[4][4] ~^ image[8][6])};
assign out_fmap[4][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][3])} + {7'd0,(kernel[0][1] ~^ image[4][4])} + {7'd0,(kernel[0][2] ~^ image[4][5])} + {7'd0,(kernel[0][3] ~^ image[4][6])} + {7'd0,(kernel[0][4] ~^ image[4][7])} + {7'd0,(kernel[1][0] ~^ image[5][3])} + {7'd0,(kernel[1][1] ~^ image[5][4])} + {7'd0,(kernel[1][2] ~^ image[5][5])} + {7'd0,(kernel[1][3] ~^ image[5][6])} + {7'd0,(kernel[1][4] ~^ image[5][7])} + {7'd0,(kernel[2][0] ~^ image[6][3])} + {7'd0,(kernel[2][1] ~^ image[6][4])} + {7'd0,(kernel[2][2] ~^ image[6][5])} + {7'd0,(kernel[2][3] ~^ image[6][6])} + {7'd0,(kernel[2][4] ~^ image[6][7])} + {7'd0,(kernel[3][0] ~^ image[7][3])} + {7'd0,(kernel[3][1] ~^ image[7][4])} + {7'd0,(kernel[3][2] ~^ image[7][5])} + {7'd0,(kernel[3][3] ~^ image[7][6])} + {7'd0,(kernel[3][4] ~^ image[7][7])} + {7'd0,(kernel[4][0] ~^ image[8][3])} + {7'd0,(kernel[4][1] ~^ image[8][4])} + {7'd0,(kernel[4][2] ~^ image[8][5])} + {7'd0,(kernel[4][3] ~^ image[8][6])} + {7'd0,(kernel[4][4] ~^ image[8][7])};
assign out_fmap[4][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][4])} + {7'd0,(kernel[0][1] ~^ image[4][5])} + {7'd0,(kernel[0][2] ~^ image[4][6])} + {7'd0,(kernel[0][3] ~^ image[4][7])} + {7'd0,(kernel[0][4] ~^ image[4][8])} + {7'd0,(kernel[1][0] ~^ image[5][4])} + {7'd0,(kernel[1][1] ~^ image[5][5])} + {7'd0,(kernel[1][2] ~^ image[5][6])} + {7'd0,(kernel[1][3] ~^ image[5][7])} + {7'd0,(kernel[1][4] ~^ image[5][8])} + {7'd0,(kernel[2][0] ~^ image[6][4])} + {7'd0,(kernel[2][1] ~^ image[6][5])} + {7'd0,(kernel[2][2] ~^ image[6][6])} + {7'd0,(kernel[2][3] ~^ image[6][7])} + {7'd0,(kernel[2][4] ~^ image[6][8])} + {7'd0,(kernel[3][0] ~^ image[7][4])} + {7'd0,(kernel[3][1] ~^ image[7][5])} + {7'd0,(kernel[3][2] ~^ image[7][6])} + {7'd0,(kernel[3][3] ~^ image[7][7])} + {7'd0,(kernel[3][4] ~^ image[7][8])} + {7'd0,(kernel[4][0] ~^ image[8][4])} + {7'd0,(kernel[4][1] ~^ image[8][5])} + {7'd0,(kernel[4][2] ~^ image[8][6])} + {7'd0,(kernel[4][3] ~^ image[8][7])} + {7'd0,(kernel[4][4] ~^ image[8][8])};
assign out_fmap[4][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][5])} + {7'd0,(kernel[0][1] ~^ image[4][6])} + {7'd0,(kernel[0][2] ~^ image[4][7])} + {7'd0,(kernel[0][3] ~^ image[4][8])} + {7'd0,(kernel[0][4] ~^ image[4][9])} + {7'd0,(kernel[1][0] ~^ image[5][5])} + {7'd0,(kernel[1][1] ~^ image[5][6])} + {7'd0,(kernel[1][2] ~^ image[5][7])} + {7'd0,(kernel[1][3] ~^ image[5][8])} + {7'd0,(kernel[1][4] ~^ image[5][9])} + {7'd0,(kernel[2][0] ~^ image[6][5])} + {7'd0,(kernel[2][1] ~^ image[6][6])} + {7'd0,(kernel[2][2] ~^ image[6][7])} + {7'd0,(kernel[2][3] ~^ image[6][8])} + {7'd0,(kernel[2][4] ~^ image[6][9])} + {7'd0,(kernel[3][0] ~^ image[7][5])} + {7'd0,(kernel[3][1] ~^ image[7][6])} + {7'd0,(kernel[3][2] ~^ image[7][7])} + {7'd0,(kernel[3][3] ~^ image[7][8])} + {7'd0,(kernel[3][4] ~^ image[7][9])} + {7'd0,(kernel[4][0] ~^ image[8][5])} + {7'd0,(kernel[4][1] ~^ image[8][6])} + {7'd0,(kernel[4][2] ~^ image[8][7])} + {7'd0,(kernel[4][3] ~^ image[8][8])} + {7'd0,(kernel[4][4] ~^ image[8][9])};
assign out_fmap[4][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][6])} + {7'd0,(kernel[0][1] ~^ image[4][7])} + {7'd0,(kernel[0][2] ~^ image[4][8])} + {7'd0,(kernel[0][3] ~^ image[4][9])} + {7'd0,(kernel[0][4] ~^ image[4][10])} + {7'd0,(kernel[1][0] ~^ image[5][6])} + {7'd0,(kernel[1][1] ~^ image[5][7])} + {7'd0,(kernel[1][2] ~^ image[5][8])} + {7'd0,(kernel[1][3] ~^ image[5][9])} + {7'd0,(kernel[1][4] ~^ image[5][10])} + {7'd0,(kernel[2][0] ~^ image[6][6])} + {7'd0,(kernel[2][1] ~^ image[6][7])} + {7'd0,(kernel[2][2] ~^ image[6][8])} + {7'd0,(kernel[2][3] ~^ image[6][9])} + {7'd0,(kernel[2][4] ~^ image[6][10])} + {7'd0,(kernel[3][0] ~^ image[7][6])} + {7'd0,(kernel[3][1] ~^ image[7][7])} + {7'd0,(kernel[3][2] ~^ image[7][8])} + {7'd0,(kernel[3][3] ~^ image[7][9])} + {7'd0,(kernel[3][4] ~^ image[7][10])} + {7'd0,(kernel[4][0] ~^ image[8][6])} + {7'd0,(kernel[4][1] ~^ image[8][7])} + {7'd0,(kernel[4][2] ~^ image[8][8])} + {7'd0,(kernel[4][3] ~^ image[8][9])} + {7'd0,(kernel[4][4] ~^ image[8][10])};
assign out_fmap[4][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][7])} + {7'd0,(kernel[0][1] ~^ image[4][8])} + {7'd0,(kernel[0][2] ~^ image[4][9])} + {7'd0,(kernel[0][3] ~^ image[4][10])} + {7'd0,(kernel[0][4] ~^ image[4][11])} + {7'd0,(kernel[1][0] ~^ image[5][7])} + {7'd0,(kernel[1][1] ~^ image[5][8])} + {7'd0,(kernel[1][2] ~^ image[5][9])} + {7'd0,(kernel[1][3] ~^ image[5][10])} + {7'd0,(kernel[1][4] ~^ image[5][11])} + {7'd0,(kernel[2][0] ~^ image[6][7])} + {7'd0,(kernel[2][1] ~^ image[6][8])} + {7'd0,(kernel[2][2] ~^ image[6][9])} + {7'd0,(kernel[2][3] ~^ image[6][10])} + {7'd0,(kernel[2][4] ~^ image[6][11])} + {7'd0,(kernel[3][0] ~^ image[7][7])} + {7'd0,(kernel[3][1] ~^ image[7][8])} + {7'd0,(kernel[3][2] ~^ image[7][9])} + {7'd0,(kernel[3][3] ~^ image[7][10])} + {7'd0,(kernel[3][4] ~^ image[7][11])} + {7'd0,(kernel[4][0] ~^ image[8][7])} + {7'd0,(kernel[4][1] ~^ image[8][8])} + {7'd0,(kernel[4][2] ~^ image[8][9])} + {7'd0,(kernel[4][3] ~^ image[8][10])} + {7'd0,(kernel[4][4] ~^ image[8][11])};
assign out_fmap[4][8][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][8])} + {7'd0,(kernel[0][1] ~^ image[4][9])} + {7'd0,(kernel[0][2] ~^ image[4][10])} + {7'd0,(kernel[0][3] ~^ image[4][11])} + {7'd0,(kernel[0][4] ~^ image[4][12])} + {7'd0,(kernel[1][0] ~^ image[5][8])} + {7'd0,(kernel[1][1] ~^ image[5][9])} + {7'd0,(kernel[1][2] ~^ image[5][10])} + {7'd0,(kernel[1][3] ~^ image[5][11])} + {7'd0,(kernel[1][4] ~^ image[5][12])} + {7'd0,(kernel[2][0] ~^ image[6][8])} + {7'd0,(kernel[2][1] ~^ image[6][9])} + {7'd0,(kernel[2][2] ~^ image[6][10])} + {7'd0,(kernel[2][3] ~^ image[6][11])} + {7'd0,(kernel[2][4] ~^ image[6][12])} + {7'd0,(kernel[3][0] ~^ image[7][8])} + {7'd0,(kernel[3][1] ~^ image[7][9])} + {7'd0,(kernel[3][2] ~^ image[7][10])} + {7'd0,(kernel[3][3] ~^ image[7][11])} + {7'd0,(kernel[3][4] ~^ image[7][12])} + {7'd0,(kernel[4][0] ~^ image[8][8])} + {7'd0,(kernel[4][1] ~^ image[8][9])} + {7'd0,(kernel[4][2] ~^ image[8][10])} + {7'd0,(kernel[4][3] ~^ image[8][11])} + {7'd0,(kernel[4][4] ~^ image[8][12])};
assign out_fmap[4][9][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][9])} + {7'd0,(kernel[0][1] ~^ image[4][10])} + {7'd0,(kernel[0][2] ~^ image[4][11])} + {7'd0,(kernel[0][3] ~^ image[4][12])} + {7'd0,(kernel[0][4] ~^ image[4][13])} + {7'd0,(kernel[1][0] ~^ image[5][9])} + {7'd0,(kernel[1][1] ~^ image[5][10])} + {7'd0,(kernel[1][2] ~^ image[5][11])} + {7'd0,(kernel[1][3] ~^ image[5][12])} + {7'd0,(kernel[1][4] ~^ image[5][13])} + {7'd0,(kernel[2][0] ~^ image[6][9])} + {7'd0,(kernel[2][1] ~^ image[6][10])} + {7'd0,(kernel[2][2] ~^ image[6][11])} + {7'd0,(kernel[2][3] ~^ image[6][12])} + {7'd0,(kernel[2][4] ~^ image[6][13])} + {7'd0,(kernel[3][0] ~^ image[7][9])} + {7'd0,(kernel[3][1] ~^ image[7][10])} + {7'd0,(kernel[3][2] ~^ image[7][11])} + {7'd0,(kernel[3][3] ~^ image[7][12])} + {7'd0,(kernel[3][4] ~^ image[7][13])} + {7'd0,(kernel[4][0] ~^ image[8][9])} + {7'd0,(kernel[4][1] ~^ image[8][10])} + {7'd0,(kernel[4][2] ~^ image[8][11])} + {7'd0,(kernel[4][3] ~^ image[8][12])} + {7'd0,(kernel[4][4] ~^ image[8][13])};
assign out_fmap[4][10][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][10])} + {7'd0,(kernel[0][1] ~^ image[4][11])} + {7'd0,(kernel[0][2] ~^ image[4][12])} + {7'd0,(kernel[0][3] ~^ image[4][13])} + {7'd0,(kernel[0][4] ~^ image[4][14])} + {7'd0,(kernel[1][0] ~^ image[5][10])} + {7'd0,(kernel[1][1] ~^ image[5][11])} + {7'd0,(kernel[1][2] ~^ image[5][12])} + {7'd0,(kernel[1][3] ~^ image[5][13])} + {7'd0,(kernel[1][4] ~^ image[5][14])} + {7'd0,(kernel[2][0] ~^ image[6][10])} + {7'd0,(kernel[2][1] ~^ image[6][11])} + {7'd0,(kernel[2][2] ~^ image[6][12])} + {7'd0,(kernel[2][3] ~^ image[6][13])} + {7'd0,(kernel[2][4] ~^ image[6][14])} + {7'd0,(kernel[3][0] ~^ image[7][10])} + {7'd0,(kernel[3][1] ~^ image[7][11])} + {7'd0,(kernel[3][2] ~^ image[7][12])} + {7'd0,(kernel[3][3] ~^ image[7][13])} + {7'd0,(kernel[3][4] ~^ image[7][14])} + {7'd0,(kernel[4][0] ~^ image[8][10])} + {7'd0,(kernel[4][1] ~^ image[8][11])} + {7'd0,(kernel[4][2] ~^ image[8][12])} + {7'd0,(kernel[4][3] ~^ image[8][13])} + {7'd0,(kernel[4][4] ~^ image[8][14])};
assign out_fmap[4][11][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][11])} + {7'd0,(kernel[0][1] ~^ image[4][12])} + {7'd0,(kernel[0][2] ~^ image[4][13])} + {7'd0,(kernel[0][3] ~^ image[4][14])} + {7'd0,(kernel[0][4] ~^ image[4][15])} + {7'd0,(kernel[1][0] ~^ image[5][11])} + {7'd0,(kernel[1][1] ~^ image[5][12])} + {7'd0,(kernel[1][2] ~^ image[5][13])} + {7'd0,(kernel[1][3] ~^ image[5][14])} + {7'd0,(kernel[1][4] ~^ image[5][15])} + {7'd0,(kernel[2][0] ~^ image[6][11])} + {7'd0,(kernel[2][1] ~^ image[6][12])} + {7'd0,(kernel[2][2] ~^ image[6][13])} + {7'd0,(kernel[2][3] ~^ image[6][14])} + {7'd0,(kernel[2][4] ~^ image[6][15])} + {7'd0,(kernel[3][0] ~^ image[7][11])} + {7'd0,(kernel[3][1] ~^ image[7][12])} + {7'd0,(kernel[3][2] ~^ image[7][13])} + {7'd0,(kernel[3][3] ~^ image[7][14])} + {7'd0,(kernel[3][4] ~^ image[7][15])} + {7'd0,(kernel[4][0] ~^ image[8][11])} + {7'd0,(kernel[4][1] ~^ image[8][12])} + {7'd0,(kernel[4][2] ~^ image[8][13])} + {7'd0,(kernel[4][3] ~^ image[8][14])} + {7'd0,(kernel[4][4] ~^ image[8][15])};
assign out_fmap[4][12][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][12])} + {7'd0,(kernel[0][1] ~^ image[4][13])} + {7'd0,(kernel[0][2] ~^ image[4][14])} + {7'd0,(kernel[0][3] ~^ image[4][15])} + {7'd0,(kernel[0][4] ~^ image[4][16])} + {7'd0,(kernel[1][0] ~^ image[5][12])} + {7'd0,(kernel[1][1] ~^ image[5][13])} + {7'd0,(kernel[1][2] ~^ image[5][14])} + {7'd0,(kernel[1][3] ~^ image[5][15])} + {7'd0,(kernel[1][4] ~^ image[5][16])} + {7'd0,(kernel[2][0] ~^ image[6][12])} + {7'd0,(kernel[2][1] ~^ image[6][13])} + {7'd0,(kernel[2][2] ~^ image[6][14])} + {7'd0,(kernel[2][3] ~^ image[6][15])} + {7'd0,(kernel[2][4] ~^ image[6][16])} + {7'd0,(kernel[3][0] ~^ image[7][12])} + {7'd0,(kernel[3][1] ~^ image[7][13])} + {7'd0,(kernel[3][2] ~^ image[7][14])} + {7'd0,(kernel[3][3] ~^ image[7][15])} + {7'd0,(kernel[3][4] ~^ image[7][16])} + {7'd0,(kernel[4][0] ~^ image[8][12])} + {7'd0,(kernel[4][1] ~^ image[8][13])} + {7'd0,(kernel[4][2] ~^ image[8][14])} + {7'd0,(kernel[4][3] ~^ image[8][15])} + {7'd0,(kernel[4][4] ~^ image[8][16])};
assign out_fmap[4][13][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][13])} + {7'd0,(kernel[0][1] ~^ image[4][14])} + {7'd0,(kernel[0][2] ~^ image[4][15])} + {7'd0,(kernel[0][3] ~^ image[4][16])} + {7'd0,(kernel[0][4] ~^ image[4][17])} + {7'd0,(kernel[1][0] ~^ image[5][13])} + {7'd0,(kernel[1][1] ~^ image[5][14])} + {7'd0,(kernel[1][2] ~^ image[5][15])} + {7'd0,(kernel[1][3] ~^ image[5][16])} + {7'd0,(kernel[1][4] ~^ image[5][17])} + {7'd0,(kernel[2][0] ~^ image[6][13])} + {7'd0,(kernel[2][1] ~^ image[6][14])} + {7'd0,(kernel[2][2] ~^ image[6][15])} + {7'd0,(kernel[2][3] ~^ image[6][16])} + {7'd0,(kernel[2][4] ~^ image[6][17])} + {7'd0,(kernel[3][0] ~^ image[7][13])} + {7'd0,(kernel[3][1] ~^ image[7][14])} + {7'd0,(kernel[3][2] ~^ image[7][15])} + {7'd0,(kernel[3][3] ~^ image[7][16])} + {7'd0,(kernel[3][4] ~^ image[7][17])} + {7'd0,(kernel[4][0] ~^ image[8][13])} + {7'd0,(kernel[4][1] ~^ image[8][14])} + {7'd0,(kernel[4][2] ~^ image[8][15])} + {7'd0,(kernel[4][3] ~^ image[8][16])} + {7'd0,(kernel[4][4] ~^ image[8][17])};
assign out_fmap[4][14][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][14])} + {7'd0,(kernel[0][1] ~^ image[4][15])} + {7'd0,(kernel[0][2] ~^ image[4][16])} + {7'd0,(kernel[0][3] ~^ image[4][17])} + {7'd0,(kernel[0][4] ~^ image[4][18])} + {7'd0,(kernel[1][0] ~^ image[5][14])} + {7'd0,(kernel[1][1] ~^ image[5][15])} + {7'd0,(kernel[1][2] ~^ image[5][16])} + {7'd0,(kernel[1][3] ~^ image[5][17])} + {7'd0,(kernel[1][4] ~^ image[5][18])} + {7'd0,(kernel[2][0] ~^ image[6][14])} + {7'd0,(kernel[2][1] ~^ image[6][15])} + {7'd0,(kernel[2][2] ~^ image[6][16])} + {7'd0,(kernel[2][3] ~^ image[6][17])} + {7'd0,(kernel[2][4] ~^ image[6][18])} + {7'd0,(kernel[3][0] ~^ image[7][14])} + {7'd0,(kernel[3][1] ~^ image[7][15])} + {7'd0,(kernel[3][2] ~^ image[7][16])} + {7'd0,(kernel[3][3] ~^ image[7][17])} + {7'd0,(kernel[3][4] ~^ image[7][18])} + {7'd0,(kernel[4][0] ~^ image[8][14])} + {7'd0,(kernel[4][1] ~^ image[8][15])} + {7'd0,(kernel[4][2] ~^ image[8][16])} + {7'd0,(kernel[4][3] ~^ image[8][17])} + {7'd0,(kernel[4][4] ~^ image[8][18])};
assign out_fmap[4][15][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][15])} + {7'd0,(kernel[0][1] ~^ image[4][16])} + {7'd0,(kernel[0][2] ~^ image[4][17])} + {7'd0,(kernel[0][3] ~^ image[4][18])} + {7'd0,(kernel[0][4] ~^ image[4][19])} + {7'd0,(kernel[1][0] ~^ image[5][15])} + {7'd0,(kernel[1][1] ~^ image[5][16])} + {7'd0,(kernel[1][2] ~^ image[5][17])} + {7'd0,(kernel[1][3] ~^ image[5][18])} + {7'd0,(kernel[1][4] ~^ image[5][19])} + {7'd0,(kernel[2][0] ~^ image[6][15])} + {7'd0,(kernel[2][1] ~^ image[6][16])} + {7'd0,(kernel[2][2] ~^ image[6][17])} + {7'd0,(kernel[2][3] ~^ image[6][18])} + {7'd0,(kernel[2][4] ~^ image[6][19])} + {7'd0,(kernel[3][0] ~^ image[7][15])} + {7'd0,(kernel[3][1] ~^ image[7][16])} + {7'd0,(kernel[3][2] ~^ image[7][17])} + {7'd0,(kernel[3][3] ~^ image[7][18])} + {7'd0,(kernel[3][4] ~^ image[7][19])} + {7'd0,(kernel[4][0] ~^ image[8][15])} + {7'd0,(kernel[4][1] ~^ image[8][16])} + {7'd0,(kernel[4][2] ~^ image[8][17])} + {7'd0,(kernel[4][3] ~^ image[8][18])} + {7'd0,(kernel[4][4] ~^ image[8][19])};
assign out_fmap[4][16][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][16])} + {7'd0,(kernel[0][1] ~^ image[4][17])} + {7'd0,(kernel[0][2] ~^ image[4][18])} + {7'd0,(kernel[0][3] ~^ image[4][19])} + {7'd0,(kernel[0][4] ~^ image[4][20])} + {7'd0,(kernel[1][0] ~^ image[5][16])} + {7'd0,(kernel[1][1] ~^ image[5][17])} + {7'd0,(kernel[1][2] ~^ image[5][18])} + {7'd0,(kernel[1][3] ~^ image[5][19])} + {7'd0,(kernel[1][4] ~^ image[5][20])} + {7'd0,(kernel[2][0] ~^ image[6][16])} + {7'd0,(kernel[2][1] ~^ image[6][17])} + {7'd0,(kernel[2][2] ~^ image[6][18])} + {7'd0,(kernel[2][3] ~^ image[6][19])} + {7'd0,(kernel[2][4] ~^ image[6][20])} + {7'd0,(kernel[3][0] ~^ image[7][16])} + {7'd0,(kernel[3][1] ~^ image[7][17])} + {7'd0,(kernel[3][2] ~^ image[7][18])} + {7'd0,(kernel[3][3] ~^ image[7][19])} + {7'd0,(kernel[3][4] ~^ image[7][20])} + {7'd0,(kernel[4][0] ~^ image[8][16])} + {7'd0,(kernel[4][1] ~^ image[8][17])} + {7'd0,(kernel[4][2] ~^ image[8][18])} + {7'd0,(kernel[4][3] ~^ image[8][19])} + {7'd0,(kernel[4][4] ~^ image[8][20])};
assign out_fmap[4][17][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][17])} + {7'd0,(kernel[0][1] ~^ image[4][18])} + {7'd0,(kernel[0][2] ~^ image[4][19])} + {7'd0,(kernel[0][3] ~^ image[4][20])} + {7'd0,(kernel[0][4] ~^ image[4][21])} + {7'd0,(kernel[1][0] ~^ image[5][17])} + {7'd0,(kernel[1][1] ~^ image[5][18])} + {7'd0,(kernel[1][2] ~^ image[5][19])} + {7'd0,(kernel[1][3] ~^ image[5][20])} + {7'd0,(kernel[1][4] ~^ image[5][21])} + {7'd0,(kernel[2][0] ~^ image[6][17])} + {7'd0,(kernel[2][1] ~^ image[6][18])} + {7'd0,(kernel[2][2] ~^ image[6][19])} + {7'd0,(kernel[2][3] ~^ image[6][20])} + {7'd0,(kernel[2][4] ~^ image[6][21])} + {7'd0,(kernel[3][0] ~^ image[7][17])} + {7'd0,(kernel[3][1] ~^ image[7][18])} + {7'd0,(kernel[3][2] ~^ image[7][19])} + {7'd0,(kernel[3][3] ~^ image[7][20])} + {7'd0,(kernel[3][4] ~^ image[7][21])} + {7'd0,(kernel[4][0] ~^ image[8][17])} + {7'd0,(kernel[4][1] ~^ image[8][18])} + {7'd0,(kernel[4][2] ~^ image[8][19])} + {7'd0,(kernel[4][3] ~^ image[8][20])} + {7'd0,(kernel[4][4] ~^ image[8][21])};
assign out_fmap[4][18][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][18])} + {7'd0,(kernel[0][1] ~^ image[4][19])} + {7'd0,(kernel[0][2] ~^ image[4][20])} + {7'd0,(kernel[0][3] ~^ image[4][21])} + {7'd0,(kernel[0][4] ~^ image[4][22])} + {7'd0,(kernel[1][0] ~^ image[5][18])} + {7'd0,(kernel[1][1] ~^ image[5][19])} + {7'd0,(kernel[1][2] ~^ image[5][20])} + {7'd0,(kernel[1][3] ~^ image[5][21])} + {7'd0,(kernel[1][4] ~^ image[5][22])} + {7'd0,(kernel[2][0] ~^ image[6][18])} + {7'd0,(kernel[2][1] ~^ image[6][19])} + {7'd0,(kernel[2][2] ~^ image[6][20])} + {7'd0,(kernel[2][3] ~^ image[6][21])} + {7'd0,(kernel[2][4] ~^ image[6][22])} + {7'd0,(kernel[3][0] ~^ image[7][18])} + {7'd0,(kernel[3][1] ~^ image[7][19])} + {7'd0,(kernel[3][2] ~^ image[7][20])} + {7'd0,(kernel[3][3] ~^ image[7][21])} + {7'd0,(kernel[3][4] ~^ image[7][22])} + {7'd0,(kernel[4][0] ~^ image[8][18])} + {7'd0,(kernel[4][1] ~^ image[8][19])} + {7'd0,(kernel[4][2] ~^ image[8][20])} + {7'd0,(kernel[4][3] ~^ image[8][21])} + {7'd0,(kernel[4][4] ~^ image[8][22])};
assign out_fmap[4][19][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][19])} + {7'd0,(kernel[0][1] ~^ image[4][20])} + {7'd0,(kernel[0][2] ~^ image[4][21])} + {7'd0,(kernel[0][3] ~^ image[4][22])} + {7'd0,(kernel[0][4] ~^ image[4][23])} + {7'd0,(kernel[1][0] ~^ image[5][19])} + {7'd0,(kernel[1][1] ~^ image[5][20])} + {7'd0,(kernel[1][2] ~^ image[5][21])} + {7'd0,(kernel[1][3] ~^ image[5][22])} + {7'd0,(kernel[1][4] ~^ image[5][23])} + {7'd0,(kernel[2][0] ~^ image[6][19])} + {7'd0,(kernel[2][1] ~^ image[6][20])} + {7'd0,(kernel[2][2] ~^ image[6][21])} + {7'd0,(kernel[2][3] ~^ image[6][22])} + {7'd0,(kernel[2][4] ~^ image[6][23])} + {7'd0,(kernel[3][0] ~^ image[7][19])} + {7'd0,(kernel[3][1] ~^ image[7][20])} + {7'd0,(kernel[3][2] ~^ image[7][21])} + {7'd0,(kernel[3][3] ~^ image[7][22])} + {7'd0,(kernel[3][4] ~^ image[7][23])} + {7'd0,(kernel[4][0] ~^ image[8][19])} + {7'd0,(kernel[4][1] ~^ image[8][20])} + {7'd0,(kernel[4][2] ~^ image[8][21])} + {7'd0,(kernel[4][3] ~^ image[8][22])} + {7'd0,(kernel[4][4] ~^ image[8][23])};
assign out_fmap[4][20][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][20])} + {7'd0,(kernel[0][1] ~^ image[4][21])} + {7'd0,(kernel[0][2] ~^ image[4][22])} + {7'd0,(kernel[0][3] ~^ image[4][23])} + {7'd0,(kernel[0][4] ~^ image[4][24])} + {7'd0,(kernel[1][0] ~^ image[5][20])} + {7'd0,(kernel[1][1] ~^ image[5][21])} + {7'd0,(kernel[1][2] ~^ image[5][22])} + {7'd0,(kernel[1][3] ~^ image[5][23])} + {7'd0,(kernel[1][4] ~^ image[5][24])} + {7'd0,(kernel[2][0] ~^ image[6][20])} + {7'd0,(kernel[2][1] ~^ image[6][21])} + {7'd0,(kernel[2][2] ~^ image[6][22])} + {7'd0,(kernel[2][3] ~^ image[6][23])} + {7'd0,(kernel[2][4] ~^ image[6][24])} + {7'd0,(kernel[3][0] ~^ image[7][20])} + {7'd0,(kernel[3][1] ~^ image[7][21])} + {7'd0,(kernel[3][2] ~^ image[7][22])} + {7'd0,(kernel[3][3] ~^ image[7][23])} + {7'd0,(kernel[3][4] ~^ image[7][24])} + {7'd0,(kernel[4][0] ~^ image[8][20])} + {7'd0,(kernel[4][1] ~^ image[8][21])} + {7'd0,(kernel[4][2] ~^ image[8][22])} + {7'd0,(kernel[4][3] ~^ image[8][23])} + {7'd0,(kernel[4][4] ~^ image[8][24])};
assign out_fmap[4][21][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][21])} + {7'd0,(kernel[0][1] ~^ image[4][22])} + {7'd0,(kernel[0][2] ~^ image[4][23])} + {7'd0,(kernel[0][3] ~^ image[4][24])} + {7'd0,(kernel[0][4] ~^ image[4][25])} + {7'd0,(kernel[1][0] ~^ image[5][21])} + {7'd0,(kernel[1][1] ~^ image[5][22])} + {7'd0,(kernel[1][2] ~^ image[5][23])} + {7'd0,(kernel[1][3] ~^ image[5][24])} + {7'd0,(kernel[1][4] ~^ image[5][25])} + {7'd0,(kernel[2][0] ~^ image[6][21])} + {7'd0,(kernel[2][1] ~^ image[6][22])} + {7'd0,(kernel[2][2] ~^ image[6][23])} + {7'd0,(kernel[2][3] ~^ image[6][24])} + {7'd0,(kernel[2][4] ~^ image[6][25])} + {7'd0,(kernel[3][0] ~^ image[7][21])} + {7'd0,(kernel[3][1] ~^ image[7][22])} + {7'd0,(kernel[3][2] ~^ image[7][23])} + {7'd0,(kernel[3][3] ~^ image[7][24])} + {7'd0,(kernel[3][4] ~^ image[7][25])} + {7'd0,(kernel[4][0] ~^ image[8][21])} + {7'd0,(kernel[4][1] ~^ image[8][22])} + {7'd0,(kernel[4][2] ~^ image[8][23])} + {7'd0,(kernel[4][3] ~^ image[8][24])} + {7'd0,(kernel[4][4] ~^ image[8][25])};
assign out_fmap[4][22][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][22])} + {7'd0,(kernel[0][1] ~^ image[4][23])} + {7'd0,(kernel[0][2] ~^ image[4][24])} + {7'd0,(kernel[0][3] ~^ image[4][25])} + {7'd0,(kernel[0][4] ~^ image[4][26])} + {7'd0,(kernel[1][0] ~^ image[5][22])} + {7'd0,(kernel[1][1] ~^ image[5][23])} + {7'd0,(kernel[1][2] ~^ image[5][24])} + {7'd0,(kernel[1][3] ~^ image[5][25])} + {7'd0,(kernel[1][4] ~^ image[5][26])} + {7'd0,(kernel[2][0] ~^ image[6][22])} + {7'd0,(kernel[2][1] ~^ image[6][23])} + {7'd0,(kernel[2][2] ~^ image[6][24])} + {7'd0,(kernel[2][3] ~^ image[6][25])} + {7'd0,(kernel[2][4] ~^ image[6][26])} + {7'd0,(kernel[3][0] ~^ image[7][22])} + {7'd0,(kernel[3][1] ~^ image[7][23])} + {7'd0,(kernel[3][2] ~^ image[7][24])} + {7'd0,(kernel[3][3] ~^ image[7][25])} + {7'd0,(kernel[3][4] ~^ image[7][26])} + {7'd0,(kernel[4][0] ~^ image[8][22])} + {7'd0,(kernel[4][1] ~^ image[8][23])} + {7'd0,(kernel[4][2] ~^ image[8][24])} + {7'd0,(kernel[4][3] ~^ image[8][25])} + {7'd0,(kernel[4][4] ~^ image[8][26])};
assign out_fmap[4][23][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[4][23])} + {7'd0,(kernel[0][1] ~^ image[4][24])} + {7'd0,(kernel[0][2] ~^ image[4][25])} + {7'd0,(kernel[0][3] ~^ image[4][26])} + {7'd0,(kernel[0][4] ~^ image[4][27])} + {7'd0,(kernel[1][0] ~^ image[5][23])} + {7'd0,(kernel[1][1] ~^ image[5][24])} + {7'd0,(kernel[1][2] ~^ image[5][25])} + {7'd0,(kernel[1][3] ~^ image[5][26])} + {7'd0,(kernel[1][4] ~^ image[5][27])} + {7'd0,(kernel[2][0] ~^ image[6][23])} + {7'd0,(kernel[2][1] ~^ image[6][24])} + {7'd0,(kernel[2][2] ~^ image[6][25])} + {7'd0,(kernel[2][3] ~^ image[6][26])} + {7'd0,(kernel[2][4] ~^ image[6][27])} + {7'd0,(kernel[3][0] ~^ image[7][23])} + {7'd0,(kernel[3][1] ~^ image[7][24])} + {7'd0,(kernel[3][2] ~^ image[7][25])} + {7'd0,(kernel[3][3] ~^ image[7][26])} + {7'd0,(kernel[3][4] ~^ image[7][27])} + {7'd0,(kernel[4][0] ~^ image[8][23])} + {7'd0,(kernel[4][1] ~^ image[8][24])} + {7'd0,(kernel[4][2] ~^ image[8][25])} + {7'd0,(kernel[4][3] ~^ image[8][26])} + {7'd0,(kernel[4][4] ~^ image[8][27])};
assign out_fmap[5][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][0])} + {7'd0,(kernel[0][1] ~^ image[5][1])} + {7'd0,(kernel[0][2] ~^ image[5][2])} + {7'd0,(kernel[0][3] ~^ image[5][3])} + {7'd0,(kernel[0][4] ~^ image[5][4])} + {7'd0,(kernel[1][0] ~^ image[6][0])} + {7'd0,(kernel[1][1] ~^ image[6][1])} + {7'd0,(kernel[1][2] ~^ image[6][2])} + {7'd0,(kernel[1][3] ~^ image[6][3])} + {7'd0,(kernel[1][4] ~^ image[6][4])} + {7'd0,(kernel[2][0] ~^ image[7][0])} + {7'd0,(kernel[2][1] ~^ image[7][1])} + {7'd0,(kernel[2][2] ~^ image[7][2])} + {7'd0,(kernel[2][3] ~^ image[7][3])} + {7'd0,(kernel[2][4] ~^ image[7][4])} + {7'd0,(kernel[3][0] ~^ image[8][0])} + {7'd0,(kernel[3][1] ~^ image[8][1])} + {7'd0,(kernel[3][2] ~^ image[8][2])} + {7'd0,(kernel[3][3] ~^ image[8][3])} + {7'd0,(kernel[3][4] ~^ image[8][4])} + {7'd0,(kernel[4][0] ~^ image[9][0])} + {7'd0,(kernel[4][1] ~^ image[9][1])} + {7'd0,(kernel[4][2] ~^ image[9][2])} + {7'd0,(kernel[4][3] ~^ image[9][3])} + {7'd0,(kernel[4][4] ~^ image[9][4])};
assign out_fmap[5][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][1])} + {7'd0,(kernel[0][1] ~^ image[5][2])} + {7'd0,(kernel[0][2] ~^ image[5][3])} + {7'd0,(kernel[0][3] ~^ image[5][4])} + {7'd0,(kernel[0][4] ~^ image[5][5])} + {7'd0,(kernel[1][0] ~^ image[6][1])} + {7'd0,(kernel[1][1] ~^ image[6][2])} + {7'd0,(kernel[1][2] ~^ image[6][3])} + {7'd0,(kernel[1][3] ~^ image[6][4])} + {7'd0,(kernel[1][4] ~^ image[6][5])} + {7'd0,(kernel[2][0] ~^ image[7][1])} + {7'd0,(kernel[2][1] ~^ image[7][2])} + {7'd0,(kernel[2][2] ~^ image[7][3])} + {7'd0,(kernel[2][3] ~^ image[7][4])} + {7'd0,(kernel[2][4] ~^ image[7][5])} + {7'd0,(kernel[3][0] ~^ image[8][1])} + {7'd0,(kernel[3][1] ~^ image[8][2])} + {7'd0,(kernel[3][2] ~^ image[8][3])} + {7'd0,(kernel[3][3] ~^ image[8][4])} + {7'd0,(kernel[3][4] ~^ image[8][5])} + {7'd0,(kernel[4][0] ~^ image[9][1])} + {7'd0,(kernel[4][1] ~^ image[9][2])} + {7'd0,(kernel[4][2] ~^ image[9][3])} + {7'd0,(kernel[4][3] ~^ image[9][4])} + {7'd0,(kernel[4][4] ~^ image[9][5])};
assign out_fmap[5][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][2])} + {7'd0,(kernel[0][1] ~^ image[5][3])} + {7'd0,(kernel[0][2] ~^ image[5][4])} + {7'd0,(kernel[0][3] ~^ image[5][5])} + {7'd0,(kernel[0][4] ~^ image[5][6])} + {7'd0,(kernel[1][0] ~^ image[6][2])} + {7'd0,(kernel[1][1] ~^ image[6][3])} + {7'd0,(kernel[1][2] ~^ image[6][4])} + {7'd0,(kernel[1][3] ~^ image[6][5])} + {7'd0,(kernel[1][4] ~^ image[6][6])} + {7'd0,(kernel[2][0] ~^ image[7][2])} + {7'd0,(kernel[2][1] ~^ image[7][3])} + {7'd0,(kernel[2][2] ~^ image[7][4])} + {7'd0,(kernel[2][3] ~^ image[7][5])} + {7'd0,(kernel[2][4] ~^ image[7][6])} + {7'd0,(kernel[3][0] ~^ image[8][2])} + {7'd0,(kernel[3][1] ~^ image[8][3])} + {7'd0,(kernel[3][2] ~^ image[8][4])} + {7'd0,(kernel[3][3] ~^ image[8][5])} + {7'd0,(kernel[3][4] ~^ image[8][6])} + {7'd0,(kernel[4][0] ~^ image[9][2])} + {7'd0,(kernel[4][1] ~^ image[9][3])} + {7'd0,(kernel[4][2] ~^ image[9][4])} + {7'd0,(kernel[4][3] ~^ image[9][5])} + {7'd0,(kernel[4][4] ~^ image[9][6])};
assign out_fmap[5][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][3])} + {7'd0,(kernel[0][1] ~^ image[5][4])} + {7'd0,(kernel[0][2] ~^ image[5][5])} + {7'd0,(kernel[0][3] ~^ image[5][6])} + {7'd0,(kernel[0][4] ~^ image[5][7])} + {7'd0,(kernel[1][0] ~^ image[6][3])} + {7'd0,(kernel[1][1] ~^ image[6][4])} + {7'd0,(kernel[1][2] ~^ image[6][5])} + {7'd0,(kernel[1][3] ~^ image[6][6])} + {7'd0,(kernel[1][4] ~^ image[6][7])} + {7'd0,(kernel[2][0] ~^ image[7][3])} + {7'd0,(kernel[2][1] ~^ image[7][4])} + {7'd0,(kernel[2][2] ~^ image[7][5])} + {7'd0,(kernel[2][3] ~^ image[7][6])} + {7'd0,(kernel[2][4] ~^ image[7][7])} + {7'd0,(kernel[3][0] ~^ image[8][3])} + {7'd0,(kernel[3][1] ~^ image[8][4])} + {7'd0,(kernel[3][2] ~^ image[8][5])} + {7'd0,(kernel[3][3] ~^ image[8][6])} + {7'd0,(kernel[3][4] ~^ image[8][7])} + {7'd0,(kernel[4][0] ~^ image[9][3])} + {7'd0,(kernel[4][1] ~^ image[9][4])} + {7'd0,(kernel[4][2] ~^ image[9][5])} + {7'd0,(kernel[4][3] ~^ image[9][6])} + {7'd0,(kernel[4][4] ~^ image[9][7])};
assign out_fmap[5][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][4])} + {7'd0,(kernel[0][1] ~^ image[5][5])} + {7'd0,(kernel[0][2] ~^ image[5][6])} + {7'd0,(kernel[0][3] ~^ image[5][7])} + {7'd0,(kernel[0][4] ~^ image[5][8])} + {7'd0,(kernel[1][0] ~^ image[6][4])} + {7'd0,(kernel[1][1] ~^ image[6][5])} + {7'd0,(kernel[1][2] ~^ image[6][6])} + {7'd0,(kernel[1][3] ~^ image[6][7])} + {7'd0,(kernel[1][4] ~^ image[6][8])} + {7'd0,(kernel[2][0] ~^ image[7][4])} + {7'd0,(kernel[2][1] ~^ image[7][5])} + {7'd0,(kernel[2][2] ~^ image[7][6])} + {7'd0,(kernel[2][3] ~^ image[7][7])} + {7'd0,(kernel[2][4] ~^ image[7][8])} + {7'd0,(kernel[3][0] ~^ image[8][4])} + {7'd0,(kernel[3][1] ~^ image[8][5])} + {7'd0,(kernel[3][2] ~^ image[8][6])} + {7'd0,(kernel[3][3] ~^ image[8][7])} + {7'd0,(kernel[3][4] ~^ image[8][8])} + {7'd0,(kernel[4][0] ~^ image[9][4])} + {7'd0,(kernel[4][1] ~^ image[9][5])} + {7'd0,(kernel[4][2] ~^ image[9][6])} + {7'd0,(kernel[4][3] ~^ image[9][7])} + {7'd0,(kernel[4][4] ~^ image[9][8])};
assign out_fmap[5][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][5])} + {7'd0,(kernel[0][1] ~^ image[5][6])} + {7'd0,(kernel[0][2] ~^ image[5][7])} + {7'd0,(kernel[0][3] ~^ image[5][8])} + {7'd0,(kernel[0][4] ~^ image[5][9])} + {7'd0,(kernel[1][0] ~^ image[6][5])} + {7'd0,(kernel[1][1] ~^ image[6][6])} + {7'd0,(kernel[1][2] ~^ image[6][7])} + {7'd0,(kernel[1][3] ~^ image[6][8])} + {7'd0,(kernel[1][4] ~^ image[6][9])} + {7'd0,(kernel[2][0] ~^ image[7][5])} + {7'd0,(kernel[2][1] ~^ image[7][6])} + {7'd0,(kernel[2][2] ~^ image[7][7])} + {7'd0,(kernel[2][3] ~^ image[7][8])} + {7'd0,(kernel[2][4] ~^ image[7][9])} + {7'd0,(kernel[3][0] ~^ image[8][5])} + {7'd0,(kernel[3][1] ~^ image[8][6])} + {7'd0,(kernel[3][2] ~^ image[8][7])} + {7'd0,(kernel[3][3] ~^ image[8][8])} + {7'd0,(kernel[3][4] ~^ image[8][9])} + {7'd0,(kernel[4][0] ~^ image[9][5])} + {7'd0,(kernel[4][1] ~^ image[9][6])} + {7'd0,(kernel[4][2] ~^ image[9][7])} + {7'd0,(kernel[4][3] ~^ image[9][8])} + {7'd0,(kernel[4][4] ~^ image[9][9])};
assign out_fmap[5][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][6])} + {7'd0,(kernel[0][1] ~^ image[5][7])} + {7'd0,(kernel[0][2] ~^ image[5][8])} + {7'd0,(kernel[0][3] ~^ image[5][9])} + {7'd0,(kernel[0][4] ~^ image[5][10])} + {7'd0,(kernel[1][0] ~^ image[6][6])} + {7'd0,(kernel[1][1] ~^ image[6][7])} + {7'd0,(kernel[1][2] ~^ image[6][8])} + {7'd0,(kernel[1][3] ~^ image[6][9])} + {7'd0,(kernel[1][4] ~^ image[6][10])} + {7'd0,(kernel[2][0] ~^ image[7][6])} + {7'd0,(kernel[2][1] ~^ image[7][7])} + {7'd0,(kernel[2][2] ~^ image[7][8])} + {7'd0,(kernel[2][3] ~^ image[7][9])} + {7'd0,(kernel[2][4] ~^ image[7][10])} + {7'd0,(kernel[3][0] ~^ image[8][6])} + {7'd0,(kernel[3][1] ~^ image[8][7])} + {7'd0,(kernel[3][2] ~^ image[8][8])} + {7'd0,(kernel[3][3] ~^ image[8][9])} + {7'd0,(kernel[3][4] ~^ image[8][10])} + {7'd0,(kernel[4][0] ~^ image[9][6])} + {7'd0,(kernel[4][1] ~^ image[9][7])} + {7'd0,(kernel[4][2] ~^ image[9][8])} + {7'd0,(kernel[4][3] ~^ image[9][9])} + {7'd0,(kernel[4][4] ~^ image[9][10])};
assign out_fmap[5][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][7])} + {7'd0,(kernel[0][1] ~^ image[5][8])} + {7'd0,(kernel[0][2] ~^ image[5][9])} + {7'd0,(kernel[0][3] ~^ image[5][10])} + {7'd0,(kernel[0][4] ~^ image[5][11])} + {7'd0,(kernel[1][0] ~^ image[6][7])} + {7'd0,(kernel[1][1] ~^ image[6][8])} + {7'd0,(kernel[1][2] ~^ image[6][9])} + {7'd0,(kernel[1][3] ~^ image[6][10])} + {7'd0,(kernel[1][4] ~^ image[6][11])} + {7'd0,(kernel[2][0] ~^ image[7][7])} + {7'd0,(kernel[2][1] ~^ image[7][8])} + {7'd0,(kernel[2][2] ~^ image[7][9])} + {7'd0,(kernel[2][3] ~^ image[7][10])} + {7'd0,(kernel[2][4] ~^ image[7][11])} + {7'd0,(kernel[3][0] ~^ image[8][7])} + {7'd0,(kernel[3][1] ~^ image[8][8])} + {7'd0,(kernel[3][2] ~^ image[8][9])} + {7'd0,(kernel[3][3] ~^ image[8][10])} + {7'd0,(kernel[3][4] ~^ image[8][11])} + {7'd0,(kernel[4][0] ~^ image[9][7])} + {7'd0,(kernel[4][1] ~^ image[9][8])} + {7'd0,(kernel[4][2] ~^ image[9][9])} + {7'd0,(kernel[4][3] ~^ image[9][10])} + {7'd0,(kernel[4][4] ~^ image[9][11])};
assign out_fmap[5][8][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][8])} + {7'd0,(kernel[0][1] ~^ image[5][9])} + {7'd0,(kernel[0][2] ~^ image[5][10])} + {7'd0,(kernel[0][3] ~^ image[5][11])} + {7'd0,(kernel[0][4] ~^ image[5][12])} + {7'd0,(kernel[1][0] ~^ image[6][8])} + {7'd0,(kernel[1][1] ~^ image[6][9])} + {7'd0,(kernel[1][2] ~^ image[6][10])} + {7'd0,(kernel[1][3] ~^ image[6][11])} + {7'd0,(kernel[1][4] ~^ image[6][12])} + {7'd0,(kernel[2][0] ~^ image[7][8])} + {7'd0,(kernel[2][1] ~^ image[7][9])} + {7'd0,(kernel[2][2] ~^ image[7][10])} + {7'd0,(kernel[2][3] ~^ image[7][11])} + {7'd0,(kernel[2][4] ~^ image[7][12])} + {7'd0,(kernel[3][0] ~^ image[8][8])} + {7'd0,(kernel[3][1] ~^ image[8][9])} + {7'd0,(kernel[3][2] ~^ image[8][10])} + {7'd0,(kernel[3][3] ~^ image[8][11])} + {7'd0,(kernel[3][4] ~^ image[8][12])} + {7'd0,(kernel[4][0] ~^ image[9][8])} + {7'd0,(kernel[4][1] ~^ image[9][9])} + {7'd0,(kernel[4][2] ~^ image[9][10])} + {7'd0,(kernel[4][3] ~^ image[9][11])} + {7'd0,(kernel[4][4] ~^ image[9][12])};
assign out_fmap[5][9][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][9])} + {7'd0,(kernel[0][1] ~^ image[5][10])} + {7'd0,(kernel[0][2] ~^ image[5][11])} + {7'd0,(kernel[0][3] ~^ image[5][12])} + {7'd0,(kernel[0][4] ~^ image[5][13])} + {7'd0,(kernel[1][0] ~^ image[6][9])} + {7'd0,(kernel[1][1] ~^ image[6][10])} + {7'd0,(kernel[1][2] ~^ image[6][11])} + {7'd0,(kernel[1][3] ~^ image[6][12])} + {7'd0,(kernel[1][4] ~^ image[6][13])} + {7'd0,(kernel[2][0] ~^ image[7][9])} + {7'd0,(kernel[2][1] ~^ image[7][10])} + {7'd0,(kernel[2][2] ~^ image[7][11])} + {7'd0,(kernel[2][3] ~^ image[7][12])} + {7'd0,(kernel[2][4] ~^ image[7][13])} + {7'd0,(kernel[3][0] ~^ image[8][9])} + {7'd0,(kernel[3][1] ~^ image[8][10])} + {7'd0,(kernel[3][2] ~^ image[8][11])} + {7'd0,(kernel[3][3] ~^ image[8][12])} + {7'd0,(kernel[3][4] ~^ image[8][13])} + {7'd0,(kernel[4][0] ~^ image[9][9])} + {7'd0,(kernel[4][1] ~^ image[9][10])} + {7'd0,(kernel[4][2] ~^ image[9][11])} + {7'd0,(kernel[4][3] ~^ image[9][12])} + {7'd0,(kernel[4][4] ~^ image[9][13])};
assign out_fmap[5][10][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][10])} + {7'd0,(kernel[0][1] ~^ image[5][11])} + {7'd0,(kernel[0][2] ~^ image[5][12])} + {7'd0,(kernel[0][3] ~^ image[5][13])} + {7'd0,(kernel[0][4] ~^ image[5][14])} + {7'd0,(kernel[1][0] ~^ image[6][10])} + {7'd0,(kernel[1][1] ~^ image[6][11])} + {7'd0,(kernel[1][2] ~^ image[6][12])} + {7'd0,(kernel[1][3] ~^ image[6][13])} + {7'd0,(kernel[1][4] ~^ image[6][14])} + {7'd0,(kernel[2][0] ~^ image[7][10])} + {7'd0,(kernel[2][1] ~^ image[7][11])} + {7'd0,(kernel[2][2] ~^ image[7][12])} + {7'd0,(kernel[2][3] ~^ image[7][13])} + {7'd0,(kernel[2][4] ~^ image[7][14])} + {7'd0,(kernel[3][0] ~^ image[8][10])} + {7'd0,(kernel[3][1] ~^ image[8][11])} + {7'd0,(kernel[3][2] ~^ image[8][12])} + {7'd0,(kernel[3][3] ~^ image[8][13])} + {7'd0,(kernel[3][4] ~^ image[8][14])} + {7'd0,(kernel[4][0] ~^ image[9][10])} + {7'd0,(kernel[4][1] ~^ image[9][11])} + {7'd0,(kernel[4][2] ~^ image[9][12])} + {7'd0,(kernel[4][3] ~^ image[9][13])} + {7'd0,(kernel[4][4] ~^ image[9][14])};
assign out_fmap[5][11][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][11])} + {7'd0,(kernel[0][1] ~^ image[5][12])} + {7'd0,(kernel[0][2] ~^ image[5][13])} + {7'd0,(kernel[0][3] ~^ image[5][14])} + {7'd0,(kernel[0][4] ~^ image[5][15])} + {7'd0,(kernel[1][0] ~^ image[6][11])} + {7'd0,(kernel[1][1] ~^ image[6][12])} + {7'd0,(kernel[1][2] ~^ image[6][13])} + {7'd0,(kernel[1][3] ~^ image[6][14])} + {7'd0,(kernel[1][4] ~^ image[6][15])} + {7'd0,(kernel[2][0] ~^ image[7][11])} + {7'd0,(kernel[2][1] ~^ image[7][12])} + {7'd0,(kernel[2][2] ~^ image[7][13])} + {7'd0,(kernel[2][3] ~^ image[7][14])} + {7'd0,(kernel[2][4] ~^ image[7][15])} + {7'd0,(kernel[3][0] ~^ image[8][11])} + {7'd0,(kernel[3][1] ~^ image[8][12])} + {7'd0,(kernel[3][2] ~^ image[8][13])} + {7'd0,(kernel[3][3] ~^ image[8][14])} + {7'd0,(kernel[3][4] ~^ image[8][15])} + {7'd0,(kernel[4][0] ~^ image[9][11])} + {7'd0,(kernel[4][1] ~^ image[9][12])} + {7'd0,(kernel[4][2] ~^ image[9][13])} + {7'd0,(kernel[4][3] ~^ image[9][14])} + {7'd0,(kernel[4][4] ~^ image[9][15])};
assign out_fmap[5][12][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][12])} + {7'd0,(kernel[0][1] ~^ image[5][13])} + {7'd0,(kernel[0][2] ~^ image[5][14])} + {7'd0,(kernel[0][3] ~^ image[5][15])} + {7'd0,(kernel[0][4] ~^ image[5][16])} + {7'd0,(kernel[1][0] ~^ image[6][12])} + {7'd0,(kernel[1][1] ~^ image[6][13])} + {7'd0,(kernel[1][2] ~^ image[6][14])} + {7'd0,(kernel[1][3] ~^ image[6][15])} + {7'd0,(kernel[1][4] ~^ image[6][16])} + {7'd0,(kernel[2][0] ~^ image[7][12])} + {7'd0,(kernel[2][1] ~^ image[7][13])} + {7'd0,(kernel[2][2] ~^ image[7][14])} + {7'd0,(kernel[2][3] ~^ image[7][15])} + {7'd0,(kernel[2][4] ~^ image[7][16])} + {7'd0,(kernel[3][0] ~^ image[8][12])} + {7'd0,(kernel[3][1] ~^ image[8][13])} + {7'd0,(kernel[3][2] ~^ image[8][14])} + {7'd0,(kernel[3][3] ~^ image[8][15])} + {7'd0,(kernel[3][4] ~^ image[8][16])} + {7'd0,(kernel[4][0] ~^ image[9][12])} + {7'd0,(kernel[4][1] ~^ image[9][13])} + {7'd0,(kernel[4][2] ~^ image[9][14])} + {7'd0,(kernel[4][3] ~^ image[9][15])} + {7'd0,(kernel[4][4] ~^ image[9][16])};
assign out_fmap[5][13][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][13])} + {7'd0,(kernel[0][1] ~^ image[5][14])} + {7'd0,(kernel[0][2] ~^ image[5][15])} + {7'd0,(kernel[0][3] ~^ image[5][16])} + {7'd0,(kernel[0][4] ~^ image[5][17])} + {7'd0,(kernel[1][0] ~^ image[6][13])} + {7'd0,(kernel[1][1] ~^ image[6][14])} + {7'd0,(kernel[1][2] ~^ image[6][15])} + {7'd0,(kernel[1][3] ~^ image[6][16])} + {7'd0,(kernel[1][4] ~^ image[6][17])} + {7'd0,(kernel[2][0] ~^ image[7][13])} + {7'd0,(kernel[2][1] ~^ image[7][14])} + {7'd0,(kernel[2][2] ~^ image[7][15])} + {7'd0,(kernel[2][3] ~^ image[7][16])} + {7'd0,(kernel[2][4] ~^ image[7][17])} + {7'd0,(kernel[3][0] ~^ image[8][13])} + {7'd0,(kernel[3][1] ~^ image[8][14])} + {7'd0,(kernel[3][2] ~^ image[8][15])} + {7'd0,(kernel[3][3] ~^ image[8][16])} + {7'd0,(kernel[3][4] ~^ image[8][17])} + {7'd0,(kernel[4][0] ~^ image[9][13])} + {7'd0,(kernel[4][1] ~^ image[9][14])} + {7'd0,(kernel[4][2] ~^ image[9][15])} + {7'd0,(kernel[4][3] ~^ image[9][16])} + {7'd0,(kernel[4][4] ~^ image[9][17])};
assign out_fmap[5][14][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][14])} + {7'd0,(kernel[0][1] ~^ image[5][15])} + {7'd0,(kernel[0][2] ~^ image[5][16])} + {7'd0,(kernel[0][3] ~^ image[5][17])} + {7'd0,(kernel[0][4] ~^ image[5][18])} + {7'd0,(kernel[1][0] ~^ image[6][14])} + {7'd0,(kernel[1][1] ~^ image[6][15])} + {7'd0,(kernel[1][2] ~^ image[6][16])} + {7'd0,(kernel[1][3] ~^ image[6][17])} + {7'd0,(kernel[1][4] ~^ image[6][18])} + {7'd0,(kernel[2][0] ~^ image[7][14])} + {7'd0,(kernel[2][1] ~^ image[7][15])} + {7'd0,(kernel[2][2] ~^ image[7][16])} + {7'd0,(kernel[2][3] ~^ image[7][17])} + {7'd0,(kernel[2][4] ~^ image[7][18])} + {7'd0,(kernel[3][0] ~^ image[8][14])} + {7'd0,(kernel[3][1] ~^ image[8][15])} + {7'd0,(kernel[3][2] ~^ image[8][16])} + {7'd0,(kernel[3][3] ~^ image[8][17])} + {7'd0,(kernel[3][4] ~^ image[8][18])} + {7'd0,(kernel[4][0] ~^ image[9][14])} + {7'd0,(kernel[4][1] ~^ image[9][15])} + {7'd0,(kernel[4][2] ~^ image[9][16])} + {7'd0,(kernel[4][3] ~^ image[9][17])} + {7'd0,(kernel[4][4] ~^ image[9][18])};
assign out_fmap[5][15][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][15])} + {7'd0,(kernel[0][1] ~^ image[5][16])} + {7'd0,(kernel[0][2] ~^ image[5][17])} + {7'd0,(kernel[0][3] ~^ image[5][18])} + {7'd0,(kernel[0][4] ~^ image[5][19])} + {7'd0,(kernel[1][0] ~^ image[6][15])} + {7'd0,(kernel[1][1] ~^ image[6][16])} + {7'd0,(kernel[1][2] ~^ image[6][17])} + {7'd0,(kernel[1][3] ~^ image[6][18])} + {7'd0,(kernel[1][4] ~^ image[6][19])} + {7'd0,(kernel[2][0] ~^ image[7][15])} + {7'd0,(kernel[2][1] ~^ image[7][16])} + {7'd0,(kernel[2][2] ~^ image[7][17])} + {7'd0,(kernel[2][3] ~^ image[7][18])} + {7'd0,(kernel[2][4] ~^ image[7][19])} + {7'd0,(kernel[3][0] ~^ image[8][15])} + {7'd0,(kernel[3][1] ~^ image[8][16])} + {7'd0,(kernel[3][2] ~^ image[8][17])} + {7'd0,(kernel[3][3] ~^ image[8][18])} + {7'd0,(kernel[3][4] ~^ image[8][19])} + {7'd0,(kernel[4][0] ~^ image[9][15])} + {7'd0,(kernel[4][1] ~^ image[9][16])} + {7'd0,(kernel[4][2] ~^ image[9][17])} + {7'd0,(kernel[4][3] ~^ image[9][18])} + {7'd0,(kernel[4][4] ~^ image[9][19])};
assign out_fmap[5][16][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][16])} + {7'd0,(kernel[0][1] ~^ image[5][17])} + {7'd0,(kernel[0][2] ~^ image[5][18])} + {7'd0,(kernel[0][3] ~^ image[5][19])} + {7'd0,(kernel[0][4] ~^ image[5][20])} + {7'd0,(kernel[1][0] ~^ image[6][16])} + {7'd0,(kernel[1][1] ~^ image[6][17])} + {7'd0,(kernel[1][2] ~^ image[6][18])} + {7'd0,(kernel[1][3] ~^ image[6][19])} + {7'd0,(kernel[1][4] ~^ image[6][20])} + {7'd0,(kernel[2][0] ~^ image[7][16])} + {7'd0,(kernel[2][1] ~^ image[7][17])} + {7'd0,(kernel[2][2] ~^ image[7][18])} + {7'd0,(kernel[2][3] ~^ image[7][19])} + {7'd0,(kernel[2][4] ~^ image[7][20])} + {7'd0,(kernel[3][0] ~^ image[8][16])} + {7'd0,(kernel[3][1] ~^ image[8][17])} + {7'd0,(kernel[3][2] ~^ image[8][18])} + {7'd0,(kernel[3][3] ~^ image[8][19])} + {7'd0,(kernel[3][4] ~^ image[8][20])} + {7'd0,(kernel[4][0] ~^ image[9][16])} + {7'd0,(kernel[4][1] ~^ image[9][17])} + {7'd0,(kernel[4][2] ~^ image[9][18])} + {7'd0,(kernel[4][3] ~^ image[9][19])} + {7'd0,(kernel[4][4] ~^ image[9][20])};
assign out_fmap[5][17][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][17])} + {7'd0,(kernel[0][1] ~^ image[5][18])} + {7'd0,(kernel[0][2] ~^ image[5][19])} + {7'd0,(kernel[0][3] ~^ image[5][20])} + {7'd0,(kernel[0][4] ~^ image[5][21])} + {7'd0,(kernel[1][0] ~^ image[6][17])} + {7'd0,(kernel[1][1] ~^ image[6][18])} + {7'd0,(kernel[1][2] ~^ image[6][19])} + {7'd0,(kernel[1][3] ~^ image[6][20])} + {7'd0,(kernel[1][4] ~^ image[6][21])} + {7'd0,(kernel[2][0] ~^ image[7][17])} + {7'd0,(kernel[2][1] ~^ image[7][18])} + {7'd0,(kernel[2][2] ~^ image[7][19])} + {7'd0,(kernel[2][3] ~^ image[7][20])} + {7'd0,(kernel[2][4] ~^ image[7][21])} + {7'd0,(kernel[3][0] ~^ image[8][17])} + {7'd0,(kernel[3][1] ~^ image[8][18])} + {7'd0,(kernel[3][2] ~^ image[8][19])} + {7'd0,(kernel[3][3] ~^ image[8][20])} + {7'd0,(kernel[3][4] ~^ image[8][21])} + {7'd0,(kernel[4][0] ~^ image[9][17])} + {7'd0,(kernel[4][1] ~^ image[9][18])} + {7'd0,(kernel[4][2] ~^ image[9][19])} + {7'd0,(kernel[4][3] ~^ image[9][20])} + {7'd0,(kernel[4][4] ~^ image[9][21])};
assign out_fmap[5][18][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][18])} + {7'd0,(kernel[0][1] ~^ image[5][19])} + {7'd0,(kernel[0][2] ~^ image[5][20])} + {7'd0,(kernel[0][3] ~^ image[5][21])} + {7'd0,(kernel[0][4] ~^ image[5][22])} + {7'd0,(kernel[1][0] ~^ image[6][18])} + {7'd0,(kernel[1][1] ~^ image[6][19])} + {7'd0,(kernel[1][2] ~^ image[6][20])} + {7'd0,(kernel[1][3] ~^ image[6][21])} + {7'd0,(kernel[1][4] ~^ image[6][22])} + {7'd0,(kernel[2][0] ~^ image[7][18])} + {7'd0,(kernel[2][1] ~^ image[7][19])} + {7'd0,(kernel[2][2] ~^ image[7][20])} + {7'd0,(kernel[2][3] ~^ image[7][21])} + {7'd0,(kernel[2][4] ~^ image[7][22])} + {7'd0,(kernel[3][0] ~^ image[8][18])} + {7'd0,(kernel[3][1] ~^ image[8][19])} + {7'd0,(kernel[3][2] ~^ image[8][20])} + {7'd0,(kernel[3][3] ~^ image[8][21])} + {7'd0,(kernel[3][4] ~^ image[8][22])} + {7'd0,(kernel[4][0] ~^ image[9][18])} + {7'd0,(kernel[4][1] ~^ image[9][19])} + {7'd0,(kernel[4][2] ~^ image[9][20])} + {7'd0,(kernel[4][3] ~^ image[9][21])} + {7'd0,(kernel[4][4] ~^ image[9][22])};
assign out_fmap[5][19][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][19])} + {7'd0,(kernel[0][1] ~^ image[5][20])} + {7'd0,(kernel[0][2] ~^ image[5][21])} + {7'd0,(kernel[0][3] ~^ image[5][22])} + {7'd0,(kernel[0][4] ~^ image[5][23])} + {7'd0,(kernel[1][0] ~^ image[6][19])} + {7'd0,(kernel[1][1] ~^ image[6][20])} + {7'd0,(kernel[1][2] ~^ image[6][21])} + {7'd0,(kernel[1][3] ~^ image[6][22])} + {7'd0,(kernel[1][4] ~^ image[6][23])} + {7'd0,(kernel[2][0] ~^ image[7][19])} + {7'd0,(kernel[2][1] ~^ image[7][20])} + {7'd0,(kernel[2][2] ~^ image[7][21])} + {7'd0,(kernel[2][3] ~^ image[7][22])} + {7'd0,(kernel[2][4] ~^ image[7][23])} + {7'd0,(kernel[3][0] ~^ image[8][19])} + {7'd0,(kernel[3][1] ~^ image[8][20])} + {7'd0,(kernel[3][2] ~^ image[8][21])} + {7'd0,(kernel[3][3] ~^ image[8][22])} + {7'd0,(kernel[3][4] ~^ image[8][23])} + {7'd0,(kernel[4][0] ~^ image[9][19])} + {7'd0,(kernel[4][1] ~^ image[9][20])} + {7'd0,(kernel[4][2] ~^ image[9][21])} + {7'd0,(kernel[4][3] ~^ image[9][22])} + {7'd0,(kernel[4][4] ~^ image[9][23])};
assign out_fmap[5][20][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][20])} + {7'd0,(kernel[0][1] ~^ image[5][21])} + {7'd0,(kernel[0][2] ~^ image[5][22])} + {7'd0,(kernel[0][3] ~^ image[5][23])} + {7'd0,(kernel[0][4] ~^ image[5][24])} + {7'd0,(kernel[1][0] ~^ image[6][20])} + {7'd0,(kernel[1][1] ~^ image[6][21])} + {7'd0,(kernel[1][2] ~^ image[6][22])} + {7'd0,(kernel[1][3] ~^ image[6][23])} + {7'd0,(kernel[1][4] ~^ image[6][24])} + {7'd0,(kernel[2][0] ~^ image[7][20])} + {7'd0,(kernel[2][1] ~^ image[7][21])} + {7'd0,(kernel[2][2] ~^ image[7][22])} + {7'd0,(kernel[2][3] ~^ image[7][23])} + {7'd0,(kernel[2][4] ~^ image[7][24])} + {7'd0,(kernel[3][0] ~^ image[8][20])} + {7'd0,(kernel[3][1] ~^ image[8][21])} + {7'd0,(kernel[3][2] ~^ image[8][22])} + {7'd0,(kernel[3][3] ~^ image[8][23])} + {7'd0,(kernel[3][4] ~^ image[8][24])} + {7'd0,(kernel[4][0] ~^ image[9][20])} + {7'd0,(kernel[4][1] ~^ image[9][21])} + {7'd0,(kernel[4][2] ~^ image[9][22])} + {7'd0,(kernel[4][3] ~^ image[9][23])} + {7'd0,(kernel[4][4] ~^ image[9][24])};
assign out_fmap[5][21][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][21])} + {7'd0,(kernel[0][1] ~^ image[5][22])} + {7'd0,(kernel[0][2] ~^ image[5][23])} + {7'd0,(kernel[0][3] ~^ image[5][24])} + {7'd0,(kernel[0][4] ~^ image[5][25])} + {7'd0,(kernel[1][0] ~^ image[6][21])} + {7'd0,(kernel[1][1] ~^ image[6][22])} + {7'd0,(kernel[1][2] ~^ image[6][23])} + {7'd0,(kernel[1][3] ~^ image[6][24])} + {7'd0,(kernel[1][4] ~^ image[6][25])} + {7'd0,(kernel[2][0] ~^ image[7][21])} + {7'd0,(kernel[2][1] ~^ image[7][22])} + {7'd0,(kernel[2][2] ~^ image[7][23])} + {7'd0,(kernel[2][3] ~^ image[7][24])} + {7'd0,(kernel[2][4] ~^ image[7][25])} + {7'd0,(kernel[3][0] ~^ image[8][21])} + {7'd0,(kernel[3][1] ~^ image[8][22])} + {7'd0,(kernel[3][2] ~^ image[8][23])} + {7'd0,(kernel[3][3] ~^ image[8][24])} + {7'd0,(kernel[3][4] ~^ image[8][25])} + {7'd0,(kernel[4][0] ~^ image[9][21])} + {7'd0,(kernel[4][1] ~^ image[9][22])} + {7'd0,(kernel[4][2] ~^ image[9][23])} + {7'd0,(kernel[4][3] ~^ image[9][24])} + {7'd0,(kernel[4][4] ~^ image[9][25])};
assign out_fmap[5][22][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][22])} + {7'd0,(kernel[0][1] ~^ image[5][23])} + {7'd0,(kernel[0][2] ~^ image[5][24])} + {7'd0,(kernel[0][3] ~^ image[5][25])} + {7'd0,(kernel[0][4] ~^ image[5][26])} + {7'd0,(kernel[1][0] ~^ image[6][22])} + {7'd0,(kernel[1][1] ~^ image[6][23])} + {7'd0,(kernel[1][2] ~^ image[6][24])} + {7'd0,(kernel[1][3] ~^ image[6][25])} + {7'd0,(kernel[1][4] ~^ image[6][26])} + {7'd0,(kernel[2][0] ~^ image[7][22])} + {7'd0,(kernel[2][1] ~^ image[7][23])} + {7'd0,(kernel[2][2] ~^ image[7][24])} + {7'd0,(kernel[2][3] ~^ image[7][25])} + {7'd0,(kernel[2][4] ~^ image[7][26])} + {7'd0,(kernel[3][0] ~^ image[8][22])} + {7'd0,(kernel[3][1] ~^ image[8][23])} + {7'd0,(kernel[3][2] ~^ image[8][24])} + {7'd0,(kernel[3][3] ~^ image[8][25])} + {7'd0,(kernel[3][4] ~^ image[8][26])} + {7'd0,(kernel[4][0] ~^ image[9][22])} + {7'd0,(kernel[4][1] ~^ image[9][23])} + {7'd0,(kernel[4][2] ~^ image[9][24])} + {7'd0,(kernel[4][3] ~^ image[9][25])} + {7'd0,(kernel[4][4] ~^ image[9][26])};
assign out_fmap[5][23][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[5][23])} + {7'd0,(kernel[0][1] ~^ image[5][24])} + {7'd0,(kernel[0][2] ~^ image[5][25])} + {7'd0,(kernel[0][3] ~^ image[5][26])} + {7'd0,(kernel[0][4] ~^ image[5][27])} + {7'd0,(kernel[1][0] ~^ image[6][23])} + {7'd0,(kernel[1][1] ~^ image[6][24])} + {7'd0,(kernel[1][2] ~^ image[6][25])} + {7'd0,(kernel[1][3] ~^ image[6][26])} + {7'd0,(kernel[1][4] ~^ image[6][27])} + {7'd0,(kernel[2][0] ~^ image[7][23])} + {7'd0,(kernel[2][1] ~^ image[7][24])} + {7'd0,(kernel[2][2] ~^ image[7][25])} + {7'd0,(kernel[2][3] ~^ image[7][26])} + {7'd0,(kernel[2][4] ~^ image[7][27])} + {7'd0,(kernel[3][0] ~^ image[8][23])} + {7'd0,(kernel[3][1] ~^ image[8][24])} + {7'd0,(kernel[3][2] ~^ image[8][25])} + {7'd0,(kernel[3][3] ~^ image[8][26])} + {7'd0,(kernel[3][4] ~^ image[8][27])} + {7'd0,(kernel[4][0] ~^ image[9][23])} + {7'd0,(kernel[4][1] ~^ image[9][24])} + {7'd0,(kernel[4][2] ~^ image[9][25])} + {7'd0,(kernel[4][3] ~^ image[9][26])} + {7'd0,(kernel[4][4] ~^ image[9][27])};
assign out_fmap[6][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][0])} + {7'd0,(kernel[0][1] ~^ image[6][1])} + {7'd0,(kernel[0][2] ~^ image[6][2])} + {7'd0,(kernel[0][3] ~^ image[6][3])} + {7'd0,(kernel[0][4] ~^ image[6][4])} + {7'd0,(kernel[1][0] ~^ image[7][0])} + {7'd0,(kernel[1][1] ~^ image[7][1])} + {7'd0,(kernel[1][2] ~^ image[7][2])} + {7'd0,(kernel[1][3] ~^ image[7][3])} + {7'd0,(kernel[1][4] ~^ image[7][4])} + {7'd0,(kernel[2][0] ~^ image[8][0])} + {7'd0,(kernel[2][1] ~^ image[8][1])} + {7'd0,(kernel[2][2] ~^ image[8][2])} + {7'd0,(kernel[2][3] ~^ image[8][3])} + {7'd0,(kernel[2][4] ~^ image[8][4])} + {7'd0,(kernel[3][0] ~^ image[9][0])} + {7'd0,(kernel[3][1] ~^ image[9][1])} + {7'd0,(kernel[3][2] ~^ image[9][2])} + {7'd0,(kernel[3][3] ~^ image[9][3])} + {7'd0,(kernel[3][4] ~^ image[9][4])} + {7'd0,(kernel[4][0] ~^ image[10][0])} + {7'd0,(kernel[4][1] ~^ image[10][1])} + {7'd0,(kernel[4][2] ~^ image[10][2])} + {7'd0,(kernel[4][3] ~^ image[10][3])} + {7'd0,(kernel[4][4] ~^ image[10][4])};
assign out_fmap[6][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][1])} + {7'd0,(kernel[0][1] ~^ image[6][2])} + {7'd0,(kernel[0][2] ~^ image[6][3])} + {7'd0,(kernel[0][3] ~^ image[6][4])} + {7'd0,(kernel[0][4] ~^ image[6][5])} + {7'd0,(kernel[1][0] ~^ image[7][1])} + {7'd0,(kernel[1][1] ~^ image[7][2])} + {7'd0,(kernel[1][2] ~^ image[7][3])} + {7'd0,(kernel[1][3] ~^ image[7][4])} + {7'd0,(kernel[1][4] ~^ image[7][5])} + {7'd0,(kernel[2][0] ~^ image[8][1])} + {7'd0,(kernel[2][1] ~^ image[8][2])} + {7'd0,(kernel[2][2] ~^ image[8][3])} + {7'd0,(kernel[2][3] ~^ image[8][4])} + {7'd0,(kernel[2][4] ~^ image[8][5])} + {7'd0,(kernel[3][0] ~^ image[9][1])} + {7'd0,(kernel[3][1] ~^ image[9][2])} + {7'd0,(kernel[3][2] ~^ image[9][3])} + {7'd0,(kernel[3][3] ~^ image[9][4])} + {7'd0,(kernel[3][4] ~^ image[9][5])} + {7'd0,(kernel[4][0] ~^ image[10][1])} + {7'd0,(kernel[4][1] ~^ image[10][2])} + {7'd0,(kernel[4][2] ~^ image[10][3])} + {7'd0,(kernel[4][3] ~^ image[10][4])} + {7'd0,(kernel[4][4] ~^ image[10][5])};
assign out_fmap[6][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][2])} + {7'd0,(kernel[0][1] ~^ image[6][3])} + {7'd0,(kernel[0][2] ~^ image[6][4])} + {7'd0,(kernel[0][3] ~^ image[6][5])} + {7'd0,(kernel[0][4] ~^ image[6][6])} + {7'd0,(kernel[1][0] ~^ image[7][2])} + {7'd0,(kernel[1][1] ~^ image[7][3])} + {7'd0,(kernel[1][2] ~^ image[7][4])} + {7'd0,(kernel[1][3] ~^ image[7][5])} + {7'd0,(kernel[1][4] ~^ image[7][6])} + {7'd0,(kernel[2][0] ~^ image[8][2])} + {7'd0,(kernel[2][1] ~^ image[8][3])} + {7'd0,(kernel[2][2] ~^ image[8][4])} + {7'd0,(kernel[2][3] ~^ image[8][5])} + {7'd0,(kernel[2][4] ~^ image[8][6])} + {7'd0,(kernel[3][0] ~^ image[9][2])} + {7'd0,(kernel[3][1] ~^ image[9][3])} + {7'd0,(kernel[3][2] ~^ image[9][4])} + {7'd0,(kernel[3][3] ~^ image[9][5])} + {7'd0,(kernel[3][4] ~^ image[9][6])} + {7'd0,(kernel[4][0] ~^ image[10][2])} + {7'd0,(kernel[4][1] ~^ image[10][3])} + {7'd0,(kernel[4][2] ~^ image[10][4])} + {7'd0,(kernel[4][3] ~^ image[10][5])} + {7'd0,(kernel[4][4] ~^ image[10][6])};
assign out_fmap[6][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][3])} + {7'd0,(kernel[0][1] ~^ image[6][4])} + {7'd0,(kernel[0][2] ~^ image[6][5])} + {7'd0,(kernel[0][3] ~^ image[6][6])} + {7'd0,(kernel[0][4] ~^ image[6][7])} + {7'd0,(kernel[1][0] ~^ image[7][3])} + {7'd0,(kernel[1][1] ~^ image[7][4])} + {7'd0,(kernel[1][2] ~^ image[7][5])} + {7'd0,(kernel[1][3] ~^ image[7][6])} + {7'd0,(kernel[1][4] ~^ image[7][7])} + {7'd0,(kernel[2][0] ~^ image[8][3])} + {7'd0,(kernel[2][1] ~^ image[8][4])} + {7'd0,(kernel[2][2] ~^ image[8][5])} + {7'd0,(kernel[2][3] ~^ image[8][6])} + {7'd0,(kernel[2][4] ~^ image[8][7])} + {7'd0,(kernel[3][0] ~^ image[9][3])} + {7'd0,(kernel[3][1] ~^ image[9][4])} + {7'd0,(kernel[3][2] ~^ image[9][5])} + {7'd0,(kernel[3][3] ~^ image[9][6])} + {7'd0,(kernel[3][4] ~^ image[9][7])} + {7'd0,(kernel[4][0] ~^ image[10][3])} + {7'd0,(kernel[4][1] ~^ image[10][4])} + {7'd0,(kernel[4][2] ~^ image[10][5])} + {7'd0,(kernel[4][3] ~^ image[10][6])} + {7'd0,(kernel[4][4] ~^ image[10][7])};
assign out_fmap[6][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][4])} + {7'd0,(kernel[0][1] ~^ image[6][5])} + {7'd0,(kernel[0][2] ~^ image[6][6])} + {7'd0,(kernel[0][3] ~^ image[6][7])} + {7'd0,(kernel[0][4] ~^ image[6][8])} + {7'd0,(kernel[1][0] ~^ image[7][4])} + {7'd0,(kernel[1][1] ~^ image[7][5])} + {7'd0,(kernel[1][2] ~^ image[7][6])} + {7'd0,(kernel[1][3] ~^ image[7][7])} + {7'd0,(kernel[1][4] ~^ image[7][8])} + {7'd0,(kernel[2][0] ~^ image[8][4])} + {7'd0,(kernel[2][1] ~^ image[8][5])} + {7'd0,(kernel[2][2] ~^ image[8][6])} + {7'd0,(kernel[2][3] ~^ image[8][7])} + {7'd0,(kernel[2][4] ~^ image[8][8])} + {7'd0,(kernel[3][0] ~^ image[9][4])} + {7'd0,(kernel[3][1] ~^ image[9][5])} + {7'd0,(kernel[3][2] ~^ image[9][6])} + {7'd0,(kernel[3][3] ~^ image[9][7])} + {7'd0,(kernel[3][4] ~^ image[9][8])} + {7'd0,(kernel[4][0] ~^ image[10][4])} + {7'd0,(kernel[4][1] ~^ image[10][5])} + {7'd0,(kernel[4][2] ~^ image[10][6])} + {7'd0,(kernel[4][3] ~^ image[10][7])} + {7'd0,(kernel[4][4] ~^ image[10][8])};
assign out_fmap[6][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][5])} + {7'd0,(kernel[0][1] ~^ image[6][6])} + {7'd0,(kernel[0][2] ~^ image[6][7])} + {7'd0,(kernel[0][3] ~^ image[6][8])} + {7'd0,(kernel[0][4] ~^ image[6][9])} + {7'd0,(kernel[1][0] ~^ image[7][5])} + {7'd0,(kernel[1][1] ~^ image[7][6])} + {7'd0,(kernel[1][2] ~^ image[7][7])} + {7'd0,(kernel[1][3] ~^ image[7][8])} + {7'd0,(kernel[1][4] ~^ image[7][9])} + {7'd0,(kernel[2][0] ~^ image[8][5])} + {7'd0,(kernel[2][1] ~^ image[8][6])} + {7'd0,(kernel[2][2] ~^ image[8][7])} + {7'd0,(kernel[2][3] ~^ image[8][8])} + {7'd0,(kernel[2][4] ~^ image[8][9])} + {7'd0,(kernel[3][0] ~^ image[9][5])} + {7'd0,(kernel[3][1] ~^ image[9][6])} + {7'd0,(kernel[3][2] ~^ image[9][7])} + {7'd0,(kernel[3][3] ~^ image[9][8])} + {7'd0,(kernel[3][4] ~^ image[9][9])} + {7'd0,(kernel[4][0] ~^ image[10][5])} + {7'd0,(kernel[4][1] ~^ image[10][6])} + {7'd0,(kernel[4][2] ~^ image[10][7])} + {7'd0,(kernel[4][3] ~^ image[10][8])} + {7'd0,(kernel[4][4] ~^ image[10][9])};
assign out_fmap[6][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][6])} + {7'd0,(kernel[0][1] ~^ image[6][7])} + {7'd0,(kernel[0][2] ~^ image[6][8])} + {7'd0,(kernel[0][3] ~^ image[6][9])} + {7'd0,(kernel[0][4] ~^ image[6][10])} + {7'd0,(kernel[1][0] ~^ image[7][6])} + {7'd0,(kernel[1][1] ~^ image[7][7])} + {7'd0,(kernel[1][2] ~^ image[7][8])} + {7'd0,(kernel[1][3] ~^ image[7][9])} + {7'd0,(kernel[1][4] ~^ image[7][10])} + {7'd0,(kernel[2][0] ~^ image[8][6])} + {7'd0,(kernel[2][1] ~^ image[8][7])} + {7'd0,(kernel[2][2] ~^ image[8][8])} + {7'd0,(kernel[2][3] ~^ image[8][9])} + {7'd0,(kernel[2][4] ~^ image[8][10])} + {7'd0,(kernel[3][0] ~^ image[9][6])} + {7'd0,(kernel[3][1] ~^ image[9][7])} + {7'd0,(kernel[3][2] ~^ image[9][8])} + {7'd0,(kernel[3][3] ~^ image[9][9])} + {7'd0,(kernel[3][4] ~^ image[9][10])} + {7'd0,(kernel[4][0] ~^ image[10][6])} + {7'd0,(kernel[4][1] ~^ image[10][7])} + {7'd0,(kernel[4][2] ~^ image[10][8])} + {7'd0,(kernel[4][3] ~^ image[10][9])} + {7'd0,(kernel[4][4] ~^ image[10][10])};
assign out_fmap[6][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][7])} + {7'd0,(kernel[0][1] ~^ image[6][8])} + {7'd0,(kernel[0][2] ~^ image[6][9])} + {7'd0,(kernel[0][3] ~^ image[6][10])} + {7'd0,(kernel[0][4] ~^ image[6][11])} + {7'd0,(kernel[1][0] ~^ image[7][7])} + {7'd0,(kernel[1][1] ~^ image[7][8])} + {7'd0,(kernel[1][2] ~^ image[7][9])} + {7'd0,(kernel[1][3] ~^ image[7][10])} + {7'd0,(kernel[1][4] ~^ image[7][11])} + {7'd0,(kernel[2][0] ~^ image[8][7])} + {7'd0,(kernel[2][1] ~^ image[8][8])} + {7'd0,(kernel[2][2] ~^ image[8][9])} + {7'd0,(kernel[2][3] ~^ image[8][10])} + {7'd0,(kernel[2][4] ~^ image[8][11])} + {7'd0,(kernel[3][0] ~^ image[9][7])} + {7'd0,(kernel[3][1] ~^ image[9][8])} + {7'd0,(kernel[3][2] ~^ image[9][9])} + {7'd0,(kernel[3][3] ~^ image[9][10])} + {7'd0,(kernel[3][4] ~^ image[9][11])} + {7'd0,(kernel[4][0] ~^ image[10][7])} + {7'd0,(kernel[4][1] ~^ image[10][8])} + {7'd0,(kernel[4][2] ~^ image[10][9])} + {7'd0,(kernel[4][3] ~^ image[10][10])} + {7'd0,(kernel[4][4] ~^ image[10][11])};
assign out_fmap[6][8][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][8])} + {7'd0,(kernel[0][1] ~^ image[6][9])} + {7'd0,(kernel[0][2] ~^ image[6][10])} + {7'd0,(kernel[0][3] ~^ image[6][11])} + {7'd0,(kernel[0][4] ~^ image[6][12])} + {7'd0,(kernel[1][0] ~^ image[7][8])} + {7'd0,(kernel[1][1] ~^ image[7][9])} + {7'd0,(kernel[1][2] ~^ image[7][10])} + {7'd0,(kernel[1][3] ~^ image[7][11])} + {7'd0,(kernel[1][4] ~^ image[7][12])} + {7'd0,(kernel[2][0] ~^ image[8][8])} + {7'd0,(kernel[2][1] ~^ image[8][9])} + {7'd0,(kernel[2][2] ~^ image[8][10])} + {7'd0,(kernel[2][3] ~^ image[8][11])} + {7'd0,(kernel[2][4] ~^ image[8][12])} + {7'd0,(kernel[3][0] ~^ image[9][8])} + {7'd0,(kernel[3][1] ~^ image[9][9])} + {7'd0,(kernel[3][2] ~^ image[9][10])} + {7'd0,(kernel[3][3] ~^ image[9][11])} + {7'd0,(kernel[3][4] ~^ image[9][12])} + {7'd0,(kernel[4][0] ~^ image[10][8])} + {7'd0,(kernel[4][1] ~^ image[10][9])} + {7'd0,(kernel[4][2] ~^ image[10][10])} + {7'd0,(kernel[4][3] ~^ image[10][11])} + {7'd0,(kernel[4][4] ~^ image[10][12])};
assign out_fmap[6][9][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][9])} + {7'd0,(kernel[0][1] ~^ image[6][10])} + {7'd0,(kernel[0][2] ~^ image[6][11])} + {7'd0,(kernel[0][3] ~^ image[6][12])} + {7'd0,(kernel[0][4] ~^ image[6][13])} + {7'd0,(kernel[1][0] ~^ image[7][9])} + {7'd0,(kernel[1][1] ~^ image[7][10])} + {7'd0,(kernel[1][2] ~^ image[7][11])} + {7'd0,(kernel[1][3] ~^ image[7][12])} + {7'd0,(kernel[1][4] ~^ image[7][13])} + {7'd0,(kernel[2][0] ~^ image[8][9])} + {7'd0,(kernel[2][1] ~^ image[8][10])} + {7'd0,(kernel[2][2] ~^ image[8][11])} + {7'd0,(kernel[2][3] ~^ image[8][12])} + {7'd0,(kernel[2][4] ~^ image[8][13])} + {7'd0,(kernel[3][0] ~^ image[9][9])} + {7'd0,(kernel[3][1] ~^ image[9][10])} + {7'd0,(kernel[3][2] ~^ image[9][11])} + {7'd0,(kernel[3][3] ~^ image[9][12])} + {7'd0,(kernel[3][4] ~^ image[9][13])} + {7'd0,(kernel[4][0] ~^ image[10][9])} + {7'd0,(kernel[4][1] ~^ image[10][10])} + {7'd0,(kernel[4][2] ~^ image[10][11])} + {7'd0,(kernel[4][3] ~^ image[10][12])} + {7'd0,(kernel[4][4] ~^ image[10][13])};
assign out_fmap[6][10][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][10])} + {7'd0,(kernel[0][1] ~^ image[6][11])} + {7'd0,(kernel[0][2] ~^ image[6][12])} + {7'd0,(kernel[0][3] ~^ image[6][13])} + {7'd0,(kernel[0][4] ~^ image[6][14])} + {7'd0,(kernel[1][0] ~^ image[7][10])} + {7'd0,(kernel[1][1] ~^ image[7][11])} + {7'd0,(kernel[1][2] ~^ image[7][12])} + {7'd0,(kernel[1][3] ~^ image[7][13])} + {7'd0,(kernel[1][4] ~^ image[7][14])} + {7'd0,(kernel[2][0] ~^ image[8][10])} + {7'd0,(kernel[2][1] ~^ image[8][11])} + {7'd0,(kernel[2][2] ~^ image[8][12])} + {7'd0,(kernel[2][3] ~^ image[8][13])} + {7'd0,(kernel[2][4] ~^ image[8][14])} + {7'd0,(kernel[3][0] ~^ image[9][10])} + {7'd0,(kernel[3][1] ~^ image[9][11])} + {7'd0,(kernel[3][2] ~^ image[9][12])} + {7'd0,(kernel[3][3] ~^ image[9][13])} + {7'd0,(kernel[3][4] ~^ image[9][14])} + {7'd0,(kernel[4][0] ~^ image[10][10])} + {7'd0,(kernel[4][1] ~^ image[10][11])} + {7'd0,(kernel[4][2] ~^ image[10][12])} + {7'd0,(kernel[4][3] ~^ image[10][13])} + {7'd0,(kernel[4][4] ~^ image[10][14])};
assign out_fmap[6][11][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][11])} + {7'd0,(kernel[0][1] ~^ image[6][12])} + {7'd0,(kernel[0][2] ~^ image[6][13])} + {7'd0,(kernel[0][3] ~^ image[6][14])} + {7'd0,(kernel[0][4] ~^ image[6][15])} + {7'd0,(kernel[1][0] ~^ image[7][11])} + {7'd0,(kernel[1][1] ~^ image[7][12])} + {7'd0,(kernel[1][2] ~^ image[7][13])} + {7'd0,(kernel[1][3] ~^ image[7][14])} + {7'd0,(kernel[1][4] ~^ image[7][15])} + {7'd0,(kernel[2][0] ~^ image[8][11])} + {7'd0,(kernel[2][1] ~^ image[8][12])} + {7'd0,(kernel[2][2] ~^ image[8][13])} + {7'd0,(kernel[2][3] ~^ image[8][14])} + {7'd0,(kernel[2][4] ~^ image[8][15])} + {7'd0,(kernel[3][0] ~^ image[9][11])} + {7'd0,(kernel[3][1] ~^ image[9][12])} + {7'd0,(kernel[3][2] ~^ image[9][13])} + {7'd0,(kernel[3][3] ~^ image[9][14])} + {7'd0,(kernel[3][4] ~^ image[9][15])} + {7'd0,(kernel[4][0] ~^ image[10][11])} + {7'd0,(kernel[4][1] ~^ image[10][12])} + {7'd0,(kernel[4][2] ~^ image[10][13])} + {7'd0,(kernel[4][3] ~^ image[10][14])} + {7'd0,(kernel[4][4] ~^ image[10][15])};
assign out_fmap[6][12][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][12])} + {7'd0,(kernel[0][1] ~^ image[6][13])} + {7'd0,(kernel[0][2] ~^ image[6][14])} + {7'd0,(kernel[0][3] ~^ image[6][15])} + {7'd0,(kernel[0][4] ~^ image[6][16])} + {7'd0,(kernel[1][0] ~^ image[7][12])} + {7'd0,(kernel[1][1] ~^ image[7][13])} + {7'd0,(kernel[1][2] ~^ image[7][14])} + {7'd0,(kernel[1][3] ~^ image[7][15])} + {7'd0,(kernel[1][4] ~^ image[7][16])} + {7'd0,(kernel[2][0] ~^ image[8][12])} + {7'd0,(kernel[2][1] ~^ image[8][13])} + {7'd0,(kernel[2][2] ~^ image[8][14])} + {7'd0,(kernel[2][3] ~^ image[8][15])} + {7'd0,(kernel[2][4] ~^ image[8][16])} + {7'd0,(kernel[3][0] ~^ image[9][12])} + {7'd0,(kernel[3][1] ~^ image[9][13])} + {7'd0,(kernel[3][2] ~^ image[9][14])} + {7'd0,(kernel[3][3] ~^ image[9][15])} + {7'd0,(kernel[3][4] ~^ image[9][16])} + {7'd0,(kernel[4][0] ~^ image[10][12])} + {7'd0,(kernel[4][1] ~^ image[10][13])} + {7'd0,(kernel[4][2] ~^ image[10][14])} + {7'd0,(kernel[4][3] ~^ image[10][15])} + {7'd0,(kernel[4][4] ~^ image[10][16])};
assign out_fmap[6][13][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][13])} + {7'd0,(kernel[0][1] ~^ image[6][14])} + {7'd0,(kernel[0][2] ~^ image[6][15])} + {7'd0,(kernel[0][3] ~^ image[6][16])} + {7'd0,(kernel[0][4] ~^ image[6][17])} + {7'd0,(kernel[1][0] ~^ image[7][13])} + {7'd0,(kernel[1][1] ~^ image[7][14])} + {7'd0,(kernel[1][2] ~^ image[7][15])} + {7'd0,(kernel[1][3] ~^ image[7][16])} + {7'd0,(kernel[1][4] ~^ image[7][17])} + {7'd0,(kernel[2][0] ~^ image[8][13])} + {7'd0,(kernel[2][1] ~^ image[8][14])} + {7'd0,(kernel[2][2] ~^ image[8][15])} + {7'd0,(kernel[2][3] ~^ image[8][16])} + {7'd0,(kernel[2][4] ~^ image[8][17])} + {7'd0,(kernel[3][0] ~^ image[9][13])} + {7'd0,(kernel[3][1] ~^ image[9][14])} + {7'd0,(kernel[3][2] ~^ image[9][15])} + {7'd0,(kernel[3][3] ~^ image[9][16])} + {7'd0,(kernel[3][4] ~^ image[9][17])} + {7'd0,(kernel[4][0] ~^ image[10][13])} + {7'd0,(kernel[4][1] ~^ image[10][14])} + {7'd0,(kernel[4][2] ~^ image[10][15])} + {7'd0,(kernel[4][3] ~^ image[10][16])} + {7'd0,(kernel[4][4] ~^ image[10][17])};
assign out_fmap[6][14][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][14])} + {7'd0,(kernel[0][1] ~^ image[6][15])} + {7'd0,(kernel[0][2] ~^ image[6][16])} + {7'd0,(kernel[0][3] ~^ image[6][17])} + {7'd0,(kernel[0][4] ~^ image[6][18])} + {7'd0,(kernel[1][0] ~^ image[7][14])} + {7'd0,(kernel[1][1] ~^ image[7][15])} + {7'd0,(kernel[1][2] ~^ image[7][16])} + {7'd0,(kernel[1][3] ~^ image[7][17])} + {7'd0,(kernel[1][4] ~^ image[7][18])} + {7'd0,(kernel[2][0] ~^ image[8][14])} + {7'd0,(kernel[2][1] ~^ image[8][15])} + {7'd0,(kernel[2][2] ~^ image[8][16])} + {7'd0,(kernel[2][3] ~^ image[8][17])} + {7'd0,(kernel[2][4] ~^ image[8][18])} + {7'd0,(kernel[3][0] ~^ image[9][14])} + {7'd0,(kernel[3][1] ~^ image[9][15])} + {7'd0,(kernel[3][2] ~^ image[9][16])} + {7'd0,(kernel[3][3] ~^ image[9][17])} + {7'd0,(kernel[3][4] ~^ image[9][18])} + {7'd0,(kernel[4][0] ~^ image[10][14])} + {7'd0,(kernel[4][1] ~^ image[10][15])} + {7'd0,(kernel[4][2] ~^ image[10][16])} + {7'd0,(kernel[4][3] ~^ image[10][17])} + {7'd0,(kernel[4][4] ~^ image[10][18])};
assign out_fmap[6][15][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][15])} + {7'd0,(kernel[0][1] ~^ image[6][16])} + {7'd0,(kernel[0][2] ~^ image[6][17])} + {7'd0,(kernel[0][3] ~^ image[6][18])} + {7'd0,(kernel[0][4] ~^ image[6][19])} + {7'd0,(kernel[1][0] ~^ image[7][15])} + {7'd0,(kernel[1][1] ~^ image[7][16])} + {7'd0,(kernel[1][2] ~^ image[7][17])} + {7'd0,(kernel[1][3] ~^ image[7][18])} + {7'd0,(kernel[1][4] ~^ image[7][19])} + {7'd0,(kernel[2][0] ~^ image[8][15])} + {7'd0,(kernel[2][1] ~^ image[8][16])} + {7'd0,(kernel[2][2] ~^ image[8][17])} + {7'd0,(kernel[2][3] ~^ image[8][18])} + {7'd0,(kernel[2][4] ~^ image[8][19])} + {7'd0,(kernel[3][0] ~^ image[9][15])} + {7'd0,(kernel[3][1] ~^ image[9][16])} + {7'd0,(kernel[3][2] ~^ image[9][17])} + {7'd0,(kernel[3][3] ~^ image[9][18])} + {7'd0,(kernel[3][4] ~^ image[9][19])} + {7'd0,(kernel[4][0] ~^ image[10][15])} + {7'd0,(kernel[4][1] ~^ image[10][16])} + {7'd0,(kernel[4][2] ~^ image[10][17])} + {7'd0,(kernel[4][3] ~^ image[10][18])} + {7'd0,(kernel[4][4] ~^ image[10][19])};
assign out_fmap[6][16][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][16])} + {7'd0,(kernel[0][1] ~^ image[6][17])} + {7'd0,(kernel[0][2] ~^ image[6][18])} + {7'd0,(kernel[0][3] ~^ image[6][19])} + {7'd0,(kernel[0][4] ~^ image[6][20])} + {7'd0,(kernel[1][0] ~^ image[7][16])} + {7'd0,(kernel[1][1] ~^ image[7][17])} + {7'd0,(kernel[1][2] ~^ image[7][18])} + {7'd0,(kernel[1][3] ~^ image[7][19])} + {7'd0,(kernel[1][4] ~^ image[7][20])} + {7'd0,(kernel[2][0] ~^ image[8][16])} + {7'd0,(kernel[2][1] ~^ image[8][17])} + {7'd0,(kernel[2][2] ~^ image[8][18])} + {7'd0,(kernel[2][3] ~^ image[8][19])} + {7'd0,(kernel[2][4] ~^ image[8][20])} + {7'd0,(kernel[3][0] ~^ image[9][16])} + {7'd0,(kernel[3][1] ~^ image[9][17])} + {7'd0,(kernel[3][2] ~^ image[9][18])} + {7'd0,(kernel[3][3] ~^ image[9][19])} + {7'd0,(kernel[3][4] ~^ image[9][20])} + {7'd0,(kernel[4][0] ~^ image[10][16])} + {7'd0,(kernel[4][1] ~^ image[10][17])} + {7'd0,(kernel[4][2] ~^ image[10][18])} + {7'd0,(kernel[4][3] ~^ image[10][19])} + {7'd0,(kernel[4][4] ~^ image[10][20])};
assign out_fmap[6][17][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][17])} + {7'd0,(kernel[0][1] ~^ image[6][18])} + {7'd0,(kernel[0][2] ~^ image[6][19])} + {7'd0,(kernel[0][3] ~^ image[6][20])} + {7'd0,(kernel[0][4] ~^ image[6][21])} + {7'd0,(kernel[1][0] ~^ image[7][17])} + {7'd0,(kernel[1][1] ~^ image[7][18])} + {7'd0,(kernel[1][2] ~^ image[7][19])} + {7'd0,(kernel[1][3] ~^ image[7][20])} + {7'd0,(kernel[1][4] ~^ image[7][21])} + {7'd0,(kernel[2][0] ~^ image[8][17])} + {7'd0,(kernel[2][1] ~^ image[8][18])} + {7'd0,(kernel[2][2] ~^ image[8][19])} + {7'd0,(kernel[2][3] ~^ image[8][20])} + {7'd0,(kernel[2][4] ~^ image[8][21])} + {7'd0,(kernel[3][0] ~^ image[9][17])} + {7'd0,(kernel[3][1] ~^ image[9][18])} + {7'd0,(kernel[3][2] ~^ image[9][19])} + {7'd0,(kernel[3][3] ~^ image[9][20])} + {7'd0,(kernel[3][4] ~^ image[9][21])} + {7'd0,(kernel[4][0] ~^ image[10][17])} + {7'd0,(kernel[4][1] ~^ image[10][18])} + {7'd0,(kernel[4][2] ~^ image[10][19])} + {7'd0,(kernel[4][3] ~^ image[10][20])} + {7'd0,(kernel[4][4] ~^ image[10][21])};
assign out_fmap[6][18][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][18])} + {7'd0,(kernel[0][1] ~^ image[6][19])} + {7'd0,(kernel[0][2] ~^ image[6][20])} + {7'd0,(kernel[0][3] ~^ image[6][21])} + {7'd0,(kernel[0][4] ~^ image[6][22])} + {7'd0,(kernel[1][0] ~^ image[7][18])} + {7'd0,(kernel[1][1] ~^ image[7][19])} + {7'd0,(kernel[1][2] ~^ image[7][20])} + {7'd0,(kernel[1][3] ~^ image[7][21])} + {7'd0,(kernel[1][4] ~^ image[7][22])} + {7'd0,(kernel[2][0] ~^ image[8][18])} + {7'd0,(kernel[2][1] ~^ image[8][19])} + {7'd0,(kernel[2][2] ~^ image[8][20])} + {7'd0,(kernel[2][3] ~^ image[8][21])} + {7'd0,(kernel[2][4] ~^ image[8][22])} + {7'd0,(kernel[3][0] ~^ image[9][18])} + {7'd0,(kernel[3][1] ~^ image[9][19])} + {7'd0,(kernel[3][2] ~^ image[9][20])} + {7'd0,(kernel[3][3] ~^ image[9][21])} + {7'd0,(kernel[3][4] ~^ image[9][22])} + {7'd0,(kernel[4][0] ~^ image[10][18])} + {7'd0,(kernel[4][1] ~^ image[10][19])} + {7'd0,(kernel[4][2] ~^ image[10][20])} + {7'd0,(kernel[4][3] ~^ image[10][21])} + {7'd0,(kernel[4][4] ~^ image[10][22])};
assign out_fmap[6][19][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][19])} + {7'd0,(kernel[0][1] ~^ image[6][20])} + {7'd0,(kernel[0][2] ~^ image[6][21])} + {7'd0,(kernel[0][3] ~^ image[6][22])} + {7'd0,(kernel[0][4] ~^ image[6][23])} + {7'd0,(kernel[1][0] ~^ image[7][19])} + {7'd0,(kernel[1][1] ~^ image[7][20])} + {7'd0,(kernel[1][2] ~^ image[7][21])} + {7'd0,(kernel[1][3] ~^ image[7][22])} + {7'd0,(kernel[1][4] ~^ image[7][23])} + {7'd0,(kernel[2][0] ~^ image[8][19])} + {7'd0,(kernel[2][1] ~^ image[8][20])} + {7'd0,(kernel[2][2] ~^ image[8][21])} + {7'd0,(kernel[2][3] ~^ image[8][22])} + {7'd0,(kernel[2][4] ~^ image[8][23])} + {7'd0,(kernel[3][0] ~^ image[9][19])} + {7'd0,(kernel[3][1] ~^ image[9][20])} + {7'd0,(kernel[3][2] ~^ image[9][21])} + {7'd0,(kernel[3][3] ~^ image[9][22])} + {7'd0,(kernel[3][4] ~^ image[9][23])} + {7'd0,(kernel[4][0] ~^ image[10][19])} + {7'd0,(kernel[4][1] ~^ image[10][20])} + {7'd0,(kernel[4][2] ~^ image[10][21])} + {7'd0,(kernel[4][3] ~^ image[10][22])} + {7'd0,(kernel[4][4] ~^ image[10][23])};
assign out_fmap[6][20][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][20])} + {7'd0,(kernel[0][1] ~^ image[6][21])} + {7'd0,(kernel[0][2] ~^ image[6][22])} + {7'd0,(kernel[0][3] ~^ image[6][23])} + {7'd0,(kernel[0][4] ~^ image[6][24])} + {7'd0,(kernel[1][0] ~^ image[7][20])} + {7'd0,(kernel[1][1] ~^ image[7][21])} + {7'd0,(kernel[1][2] ~^ image[7][22])} + {7'd0,(kernel[1][3] ~^ image[7][23])} + {7'd0,(kernel[1][4] ~^ image[7][24])} + {7'd0,(kernel[2][0] ~^ image[8][20])} + {7'd0,(kernel[2][1] ~^ image[8][21])} + {7'd0,(kernel[2][2] ~^ image[8][22])} + {7'd0,(kernel[2][3] ~^ image[8][23])} + {7'd0,(kernel[2][4] ~^ image[8][24])} + {7'd0,(kernel[3][0] ~^ image[9][20])} + {7'd0,(kernel[3][1] ~^ image[9][21])} + {7'd0,(kernel[3][2] ~^ image[9][22])} + {7'd0,(kernel[3][3] ~^ image[9][23])} + {7'd0,(kernel[3][4] ~^ image[9][24])} + {7'd0,(kernel[4][0] ~^ image[10][20])} + {7'd0,(kernel[4][1] ~^ image[10][21])} + {7'd0,(kernel[4][2] ~^ image[10][22])} + {7'd0,(kernel[4][3] ~^ image[10][23])} + {7'd0,(kernel[4][4] ~^ image[10][24])};
assign out_fmap[6][21][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][21])} + {7'd0,(kernel[0][1] ~^ image[6][22])} + {7'd0,(kernel[0][2] ~^ image[6][23])} + {7'd0,(kernel[0][3] ~^ image[6][24])} + {7'd0,(kernel[0][4] ~^ image[6][25])} + {7'd0,(kernel[1][0] ~^ image[7][21])} + {7'd0,(kernel[1][1] ~^ image[7][22])} + {7'd0,(kernel[1][2] ~^ image[7][23])} + {7'd0,(kernel[1][3] ~^ image[7][24])} + {7'd0,(kernel[1][4] ~^ image[7][25])} + {7'd0,(kernel[2][0] ~^ image[8][21])} + {7'd0,(kernel[2][1] ~^ image[8][22])} + {7'd0,(kernel[2][2] ~^ image[8][23])} + {7'd0,(kernel[2][3] ~^ image[8][24])} + {7'd0,(kernel[2][4] ~^ image[8][25])} + {7'd0,(kernel[3][0] ~^ image[9][21])} + {7'd0,(kernel[3][1] ~^ image[9][22])} + {7'd0,(kernel[3][2] ~^ image[9][23])} + {7'd0,(kernel[3][3] ~^ image[9][24])} + {7'd0,(kernel[3][4] ~^ image[9][25])} + {7'd0,(kernel[4][0] ~^ image[10][21])} + {7'd0,(kernel[4][1] ~^ image[10][22])} + {7'd0,(kernel[4][2] ~^ image[10][23])} + {7'd0,(kernel[4][3] ~^ image[10][24])} + {7'd0,(kernel[4][4] ~^ image[10][25])};
assign out_fmap[6][22][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][22])} + {7'd0,(kernel[0][1] ~^ image[6][23])} + {7'd0,(kernel[0][2] ~^ image[6][24])} + {7'd0,(kernel[0][3] ~^ image[6][25])} + {7'd0,(kernel[0][4] ~^ image[6][26])} + {7'd0,(kernel[1][0] ~^ image[7][22])} + {7'd0,(kernel[1][1] ~^ image[7][23])} + {7'd0,(kernel[1][2] ~^ image[7][24])} + {7'd0,(kernel[1][3] ~^ image[7][25])} + {7'd0,(kernel[1][4] ~^ image[7][26])} + {7'd0,(kernel[2][0] ~^ image[8][22])} + {7'd0,(kernel[2][1] ~^ image[8][23])} + {7'd0,(kernel[2][2] ~^ image[8][24])} + {7'd0,(kernel[2][3] ~^ image[8][25])} + {7'd0,(kernel[2][4] ~^ image[8][26])} + {7'd0,(kernel[3][0] ~^ image[9][22])} + {7'd0,(kernel[3][1] ~^ image[9][23])} + {7'd0,(kernel[3][2] ~^ image[9][24])} + {7'd0,(kernel[3][3] ~^ image[9][25])} + {7'd0,(kernel[3][4] ~^ image[9][26])} + {7'd0,(kernel[4][0] ~^ image[10][22])} + {7'd0,(kernel[4][1] ~^ image[10][23])} + {7'd0,(kernel[4][2] ~^ image[10][24])} + {7'd0,(kernel[4][3] ~^ image[10][25])} + {7'd0,(kernel[4][4] ~^ image[10][26])};
assign out_fmap[6][23][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[6][23])} + {7'd0,(kernel[0][1] ~^ image[6][24])} + {7'd0,(kernel[0][2] ~^ image[6][25])} + {7'd0,(kernel[0][3] ~^ image[6][26])} + {7'd0,(kernel[0][4] ~^ image[6][27])} + {7'd0,(kernel[1][0] ~^ image[7][23])} + {7'd0,(kernel[1][1] ~^ image[7][24])} + {7'd0,(kernel[1][2] ~^ image[7][25])} + {7'd0,(kernel[1][3] ~^ image[7][26])} + {7'd0,(kernel[1][4] ~^ image[7][27])} + {7'd0,(kernel[2][0] ~^ image[8][23])} + {7'd0,(kernel[2][1] ~^ image[8][24])} + {7'd0,(kernel[2][2] ~^ image[8][25])} + {7'd0,(kernel[2][3] ~^ image[8][26])} + {7'd0,(kernel[2][4] ~^ image[8][27])} + {7'd0,(kernel[3][0] ~^ image[9][23])} + {7'd0,(kernel[3][1] ~^ image[9][24])} + {7'd0,(kernel[3][2] ~^ image[9][25])} + {7'd0,(kernel[3][3] ~^ image[9][26])} + {7'd0,(kernel[3][4] ~^ image[9][27])} + {7'd0,(kernel[4][0] ~^ image[10][23])} + {7'd0,(kernel[4][1] ~^ image[10][24])} + {7'd0,(kernel[4][2] ~^ image[10][25])} + {7'd0,(kernel[4][3] ~^ image[10][26])} + {7'd0,(kernel[4][4] ~^ image[10][27])};
assign out_fmap[7][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][0])} + {7'd0,(kernel[0][1] ~^ image[7][1])} + {7'd0,(kernel[0][2] ~^ image[7][2])} + {7'd0,(kernel[0][3] ~^ image[7][3])} + {7'd0,(kernel[0][4] ~^ image[7][4])} + {7'd0,(kernel[1][0] ~^ image[8][0])} + {7'd0,(kernel[1][1] ~^ image[8][1])} + {7'd0,(kernel[1][2] ~^ image[8][2])} + {7'd0,(kernel[1][3] ~^ image[8][3])} + {7'd0,(kernel[1][4] ~^ image[8][4])} + {7'd0,(kernel[2][0] ~^ image[9][0])} + {7'd0,(kernel[2][1] ~^ image[9][1])} + {7'd0,(kernel[2][2] ~^ image[9][2])} + {7'd0,(kernel[2][3] ~^ image[9][3])} + {7'd0,(kernel[2][4] ~^ image[9][4])} + {7'd0,(kernel[3][0] ~^ image[10][0])} + {7'd0,(kernel[3][1] ~^ image[10][1])} + {7'd0,(kernel[3][2] ~^ image[10][2])} + {7'd0,(kernel[3][3] ~^ image[10][3])} + {7'd0,(kernel[3][4] ~^ image[10][4])} + {7'd0,(kernel[4][0] ~^ image[11][0])} + {7'd0,(kernel[4][1] ~^ image[11][1])} + {7'd0,(kernel[4][2] ~^ image[11][2])} + {7'd0,(kernel[4][3] ~^ image[11][3])} + {7'd0,(kernel[4][4] ~^ image[11][4])};
assign out_fmap[7][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][1])} + {7'd0,(kernel[0][1] ~^ image[7][2])} + {7'd0,(kernel[0][2] ~^ image[7][3])} + {7'd0,(kernel[0][3] ~^ image[7][4])} + {7'd0,(kernel[0][4] ~^ image[7][5])} + {7'd0,(kernel[1][0] ~^ image[8][1])} + {7'd0,(kernel[1][1] ~^ image[8][2])} + {7'd0,(kernel[1][2] ~^ image[8][3])} + {7'd0,(kernel[1][3] ~^ image[8][4])} + {7'd0,(kernel[1][4] ~^ image[8][5])} + {7'd0,(kernel[2][0] ~^ image[9][1])} + {7'd0,(kernel[2][1] ~^ image[9][2])} + {7'd0,(kernel[2][2] ~^ image[9][3])} + {7'd0,(kernel[2][3] ~^ image[9][4])} + {7'd0,(kernel[2][4] ~^ image[9][5])} + {7'd0,(kernel[3][0] ~^ image[10][1])} + {7'd0,(kernel[3][1] ~^ image[10][2])} + {7'd0,(kernel[3][2] ~^ image[10][3])} + {7'd0,(kernel[3][3] ~^ image[10][4])} + {7'd0,(kernel[3][4] ~^ image[10][5])} + {7'd0,(kernel[4][0] ~^ image[11][1])} + {7'd0,(kernel[4][1] ~^ image[11][2])} + {7'd0,(kernel[4][2] ~^ image[11][3])} + {7'd0,(kernel[4][3] ~^ image[11][4])} + {7'd0,(kernel[4][4] ~^ image[11][5])};
assign out_fmap[7][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][2])} + {7'd0,(kernel[0][1] ~^ image[7][3])} + {7'd0,(kernel[0][2] ~^ image[7][4])} + {7'd0,(kernel[0][3] ~^ image[7][5])} + {7'd0,(kernel[0][4] ~^ image[7][6])} + {7'd0,(kernel[1][0] ~^ image[8][2])} + {7'd0,(kernel[1][1] ~^ image[8][3])} + {7'd0,(kernel[1][2] ~^ image[8][4])} + {7'd0,(kernel[1][3] ~^ image[8][5])} + {7'd0,(kernel[1][4] ~^ image[8][6])} + {7'd0,(kernel[2][0] ~^ image[9][2])} + {7'd0,(kernel[2][1] ~^ image[9][3])} + {7'd0,(kernel[2][2] ~^ image[9][4])} + {7'd0,(kernel[2][3] ~^ image[9][5])} + {7'd0,(kernel[2][4] ~^ image[9][6])} + {7'd0,(kernel[3][0] ~^ image[10][2])} + {7'd0,(kernel[3][1] ~^ image[10][3])} + {7'd0,(kernel[3][2] ~^ image[10][4])} + {7'd0,(kernel[3][3] ~^ image[10][5])} + {7'd0,(kernel[3][4] ~^ image[10][6])} + {7'd0,(kernel[4][0] ~^ image[11][2])} + {7'd0,(kernel[4][1] ~^ image[11][3])} + {7'd0,(kernel[4][2] ~^ image[11][4])} + {7'd0,(kernel[4][3] ~^ image[11][5])} + {7'd0,(kernel[4][4] ~^ image[11][6])};
assign out_fmap[7][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][3])} + {7'd0,(kernel[0][1] ~^ image[7][4])} + {7'd0,(kernel[0][2] ~^ image[7][5])} + {7'd0,(kernel[0][3] ~^ image[7][6])} + {7'd0,(kernel[0][4] ~^ image[7][7])} + {7'd0,(kernel[1][0] ~^ image[8][3])} + {7'd0,(kernel[1][1] ~^ image[8][4])} + {7'd0,(kernel[1][2] ~^ image[8][5])} + {7'd0,(kernel[1][3] ~^ image[8][6])} + {7'd0,(kernel[1][4] ~^ image[8][7])} + {7'd0,(kernel[2][0] ~^ image[9][3])} + {7'd0,(kernel[2][1] ~^ image[9][4])} + {7'd0,(kernel[2][2] ~^ image[9][5])} + {7'd0,(kernel[2][3] ~^ image[9][6])} + {7'd0,(kernel[2][4] ~^ image[9][7])} + {7'd0,(kernel[3][0] ~^ image[10][3])} + {7'd0,(kernel[3][1] ~^ image[10][4])} + {7'd0,(kernel[3][2] ~^ image[10][5])} + {7'd0,(kernel[3][3] ~^ image[10][6])} + {7'd0,(kernel[3][4] ~^ image[10][7])} + {7'd0,(kernel[4][0] ~^ image[11][3])} + {7'd0,(kernel[4][1] ~^ image[11][4])} + {7'd0,(kernel[4][2] ~^ image[11][5])} + {7'd0,(kernel[4][3] ~^ image[11][6])} + {7'd0,(kernel[4][4] ~^ image[11][7])};
assign out_fmap[7][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][4])} + {7'd0,(kernel[0][1] ~^ image[7][5])} + {7'd0,(kernel[0][2] ~^ image[7][6])} + {7'd0,(kernel[0][3] ~^ image[7][7])} + {7'd0,(kernel[0][4] ~^ image[7][8])} + {7'd0,(kernel[1][0] ~^ image[8][4])} + {7'd0,(kernel[1][1] ~^ image[8][5])} + {7'd0,(kernel[1][2] ~^ image[8][6])} + {7'd0,(kernel[1][3] ~^ image[8][7])} + {7'd0,(kernel[1][4] ~^ image[8][8])} + {7'd0,(kernel[2][0] ~^ image[9][4])} + {7'd0,(kernel[2][1] ~^ image[9][5])} + {7'd0,(kernel[2][2] ~^ image[9][6])} + {7'd0,(kernel[2][3] ~^ image[9][7])} + {7'd0,(kernel[2][4] ~^ image[9][8])} + {7'd0,(kernel[3][0] ~^ image[10][4])} + {7'd0,(kernel[3][1] ~^ image[10][5])} + {7'd0,(kernel[3][2] ~^ image[10][6])} + {7'd0,(kernel[3][3] ~^ image[10][7])} + {7'd0,(kernel[3][4] ~^ image[10][8])} + {7'd0,(kernel[4][0] ~^ image[11][4])} + {7'd0,(kernel[4][1] ~^ image[11][5])} + {7'd0,(kernel[4][2] ~^ image[11][6])} + {7'd0,(kernel[4][3] ~^ image[11][7])} + {7'd0,(kernel[4][4] ~^ image[11][8])};
assign out_fmap[7][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][5])} + {7'd0,(kernel[0][1] ~^ image[7][6])} + {7'd0,(kernel[0][2] ~^ image[7][7])} + {7'd0,(kernel[0][3] ~^ image[7][8])} + {7'd0,(kernel[0][4] ~^ image[7][9])} + {7'd0,(kernel[1][0] ~^ image[8][5])} + {7'd0,(kernel[1][1] ~^ image[8][6])} + {7'd0,(kernel[1][2] ~^ image[8][7])} + {7'd0,(kernel[1][3] ~^ image[8][8])} + {7'd0,(kernel[1][4] ~^ image[8][9])} + {7'd0,(kernel[2][0] ~^ image[9][5])} + {7'd0,(kernel[2][1] ~^ image[9][6])} + {7'd0,(kernel[2][2] ~^ image[9][7])} + {7'd0,(kernel[2][3] ~^ image[9][8])} + {7'd0,(kernel[2][4] ~^ image[9][9])} + {7'd0,(kernel[3][0] ~^ image[10][5])} + {7'd0,(kernel[3][1] ~^ image[10][6])} + {7'd0,(kernel[3][2] ~^ image[10][7])} + {7'd0,(kernel[3][3] ~^ image[10][8])} + {7'd0,(kernel[3][4] ~^ image[10][9])} + {7'd0,(kernel[4][0] ~^ image[11][5])} + {7'd0,(kernel[4][1] ~^ image[11][6])} + {7'd0,(kernel[4][2] ~^ image[11][7])} + {7'd0,(kernel[4][3] ~^ image[11][8])} + {7'd0,(kernel[4][4] ~^ image[11][9])};
assign out_fmap[7][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][6])} + {7'd0,(kernel[0][1] ~^ image[7][7])} + {7'd0,(kernel[0][2] ~^ image[7][8])} + {7'd0,(kernel[0][3] ~^ image[7][9])} + {7'd0,(kernel[0][4] ~^ image[7][10])} + {7'd0,(kernel[1][0] ~^ image[8][6])} + {7'd0,(kernel[1][1] ~^ image[8][7])} + {7'd0,(kernel[1][2] ~^ image[8][8])} + {7'd0,(kernel[1][3] ~^ image[8][9])} + {7'd0,(kernel[1][4] ~^ image[8][10])} + {7'd0,(kernel[2][0] ~^ image[9][6])} + {7'd0,(kernel[2][1] ~^ image[9][7])} + {7'd0,(kernel[2][2] ~^ image[9][8])} + {7'd0,(kernel[2][3] ~^ image[9][9])} + {7'd0,(kernel[2][4] ~^ image[9][10])} + {7'd0,(kernel[3][0] ~^ image[10][6])} + {7'd0,(kernel[3][1] ~^ image[10][7])} + {7'd0,(kernel[3][2] ~^ image[10][8])} + {7'd0,(kernel[3][3] ~^ image[10][9])} + {7'd0,(kernel[3][4] ~^ image[10][10])} + {7'd0,(kernel[4][0] ~^ image[11][6])} + {7'd0,(kernel[4][1] ~^ image[11][7])} + {7'd0,(kernel[4][2] ~^ image[11][8])} + {7'd0,(kernel[4][3] ~^ image[11][9])} + {7'd0,(kernel[4][4] ~^ image[11][10])};
assign out_fmap[7][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][7])} + {7'd0,(kernel[0][1] ~^ image[7][8])} + {7'd0,(kernel[0][2] ~^ image[7][9])} + {7'd0,(kernel[0][3] ~^ image[7][10])} + {7'd0,(kernel[0][4] ~^ image[7][11])} + {7'd0,(kernel[1][0] ~^ image[8][7])} + {7'd0,(kernel[1][1] ~^ image[8][8])} + {7'd0,(kernel[1][2] ~^ image[8][9])} + {7'd0,(kernel[1][3] ~^ image[8][10])} + {7'd0,(kernel[1][4] ~^ image[8][11])} + {7'd0,(kernel[2][0] ~^ image[9][7])} + {7'd0,(kernel[2][1] ~^ image[9][8])} + {7'd0,(kernel[2][2] ~^ image[9][9])} + {7'd0,(kernel[2][3] ~^ image[9][10])} + {7'd0,(kernel[2][4] ~^ image[9][11])} + {7'd0,(kernel[3][0] ~^ image[10][7])} + {7'd0,(kernel[3][1] ~^ image[10][8])} + {7'd0,(kernel[3][2] ~^ image[10][9])} + {7'd0,(kernel[3][3] ~^ image[10][10])} + {7'd0,(kernel[3][4] ~^ image[10][11])} + {7'd0,(kernel[4][0] ~^ image[11][7])} + {7'd0,(kernel[4][1] ~^ image[11][8])} + {7'd0,(kernel[4][2] ~^ image[11][9])} + {7'd0,(kernel[4][3] ~^ image[11][10])} + {7'd0,(kernel[4][4] ~^ image[11][11])};
assign out_fmap[7][8][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][8])} + {7'd0,(kernel[0][1] ~^ image[7][9])} + {7'd0,(kernel[0][2] ~^ image[7][10])} + {7'd0,(kernel[0][3] ~^ image[7][11])} + {7'd0,(kernel[0][4] ~^ image[7][12])} + {7'd0,(kernel[1][0] ~^ image[8][8])} + {7'd0,(kernel[1][1] ~^ image[8][9])} + {7'd0,(kernel[1][2] ~^ image[8][10])} + {7'd0,(kernel[1][3] ~^ image[8][11])} + {7'd0,(kernel[1][4] ~^ image[8][12])} + {7'd0,(kernel[2][0] ~^ image[9][8])} + {7'd0,(kernel[2][1] ~^ image[9][9])} + {7'd0,(kernel[2][2] ~^ image[9][10])} + {7'd0,(kernel[2][3] ~^ image[9][11])} + {7'd0,(kernel[2][4] ~^ image[9][12])} + {7'd0,(kernel[3][0] ~^ image[10][8])} + {7'd0,(kernel[3][1] ~^ image[10][9])} + {7'd0,(kernel[3][2] ~^ image[10][10])} + {7'd0,(kernel[3][3] ~^ image[10][11])} + {7'd0,(kernel[3][4] ~^ image[10][12])} + {7'd0,(kernel[4][0] ~^ image[11][8])} + {7'd0,(kernel[4][1] ~^ image[11][9])} + {7'd0,(kernel[4][2] ~^ image[11][10])} + {7'd0,(kernel[4][3] ~^ image[11][11])} + {7'd0,(kernel[4][4] ~^ image[11][12])};
assign out_fmap[7][9][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][9])} + {7'd0,(kernel[0][1] ~^ image[7][10])} + {7'd0,(kernel[0][2] ~^ image[7][11])} + {7'd0,(kernel[0][3] ~^ image[7][12])} + {7'd0,(kernel[0][4] ~^ image[7][13])} + {7'd0,(kernel[1][0] ~^ image[8][9])} + {7'd0,(kernel[1][1] ~^ image[8][10])} + {7'd0,(kernel[1][2] ~^ image[8][11])} + {7'd0,(kernel[1][3] ~^ image[8][12])} + {7'd0,(kernel[1][4] ~^ image[8][13])} + {7'd0,(kernel[2][0] ~^ image[9][9])} + {7'd0,(kernel[2][1] ~^ image[9][10])} + {7'd0,(kernel[2][2] ~^ image[9][11])} + {7'd0,(kernel[2][3] ~^ image[9][12])} + {7'd0,(kernel[2][4] ~^ image[9][13])} + {7'd0,(kernel[3][0] ~^ image[10][9])} + {7'd0,(kernel[3][1] ~^ image[10][10])} + {7'd0,(kernel[3][2] ~^ image[10][11])} + {7'd0,(kernel[3][3] ~^ image[10][12])} + {7'd0,(kernel[3][4] ~^ image[10][13])} + {7'd0,(kernel[4][0] ~^ image[11][9])} + {7'd0,(kernel[4][1] ~^ image[11][10])} + {7'd0,(kernel[4][2] ~^ image[11][11])} + {7'd0,(kernel[4][3] ~^ image[11][12])} + {7'd0,(kernel[4][4] ~^ image[11][13])};
assign out_fmap[7][10][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][10])} + {7'd0,(kernel[0][1] ~^ image[7][11])} + {7'd0,(kernel[0][2] ~^ image[7][12])} + {7'd0,(kernel[0][3] ~^ image[7][13])} + {7'd0,(kernel[0][4] ~^ image[7][14])} + {7'd0,(kernel[1][0] ~^ image[8][10])} + {7'd0,(kernel[1][1] ~^ image[8][11])} + {7'd0,(kernel[1][2] ~^ image[8][12])} + {7'd0,(kernel[1][3] ~^ image[8][13])} + {7'd0,(kernel[1][4] ~^ image[8][14])} + {7'd0,(kernel[2][0] ~^ image[9][10])} + {7'd0,(kernel[2][1] ~^ image[9][11])} + {7'd0,(kernel[2][2] ~^ image[9][12])} + {7'd0,(kernel[2][3] ~^ image[9][13])} + {7'd0,(kernel[2][4] ~^ image[9][14])} + {7'd0,(kernel[3][0] ~^ image[10][10])} + {7'd0,(kernel[3][1] ~^ image[10][11])} + {7'd0,(kernel[3][2] ~^ image[10][12])} + {7'd0,(kernel[3][3] ~^ image[10][13])} + {7'd0,(kernel[3][4] ~^ image[10][14])} + {7'd0,(kernel[4][0] ~^ image[11][10])} + {7'd0,(kernel[4][1] ~^ image[11][11])} + {7'd0,(kernel[4][2] ~^ image[11][12])} + {7'd0,(kernel[4][3] ~^ image[11][13])} + {7'd0,(kernel[4][4] ~^ image[11][14])};
assign out_fmap[7][11][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][11])} + {7'd0,(kernel[0][1] ~^ image[7][12])} + {7'd0,(kernel[0][2] ~^ image[7][13])} + {7'd0,(kernel[0][3] ~^ image[7][14])} + {7'd0,(kernel[0][4] ~^ image[7][15])} + {7'd0,(kernel[1][0] ~^ image[8][11])} + {7'd0,(kernel[1][1] ~^ image[8][12])} + {7'd0,(kernel[1][2] ~^ image[8][13])} + {7'd0,(kernel[1][3] ~^ image[8][14])} + {7'd0,(kernel[1][4] ~^ image[8][15])} + {7'd0,(kernel[2][0] ~^ image[9][11])} + {7'd0,(kernel[2][1] ~^ image[9][12])} + {7'd0,(kernel[2][2] ~^ image[9][13])} + {7'd0,(kernel[2][3] ~^ image[9][14])} + {7'd0,(kernel[2][4] ~^ image[9][15])} + {7'd0,(kernel[3][0] ~^ image[10][11])} + {7'd0,(kernel[3][1] ~^ image[10][12])} + {7'd0,(kernel[3][2] ~^ image[10][13])} + {7'd0,(kernel[3][3] ~^ image[10][14])} + {7'd0,(kernel[3][4] ~^ image[10][15])} + {7'd0,(kernel[4][0] ~^ image[11][11])} + {7'd0,(kernel[4][1] ~^ image[11][12])} + {7'd0,(kernel[4][2] ~^ image[11][13])} + {7'd0,(kernel[4][3] ~^ image[11][14])} + {7'd0,(kernel[4][4] ~^ image[11][15])};
assign out_fmap[7][12][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][12])} + {7'd0,(kernel[0][1] ~^ image[7][13])} + {7'd0,(kernel[0][2] ~^ image[7][14])} + {7'd0,(kernel[0][3] ~^ image[7][15])} + {7'd0,(kernel[0][4] ~^ image[7][16])} + {7'd0,(kernel[1][0] ~^ image[8][12])} + {7'd0,(kernel[1][1] ~^ image[8][13])} + {7'd0,(kernel[1][2] ~^ image[8][14])} + {7'd0,(kernel[1][3] ~^ image[8][15])} + {7'd0,(kernel[1][4] ~^ image[8][16])} + {7'd0,(kernel[2][0] ~^ image[9][12])} + {7'd0,(kernel[2][1] ~^ image[9][13])} + {7'd0,(kernel[2][2] ~^ image[9][14])} + {7'd0,(kernel[2][3] ~^ image[9][15])} + {7'd0,(kernel[2][4] ~^ image[9][16])} + {7'd0,(kernel[3][0] ~^ image[10][12])} + {7'd0,(kernel[3][1] ~^ image[10][13])} + {7'd0,(kernel[3][2] ~^ image[10][14])} + {7'd0,(kernel[3][3] ~^ image[10][15])} + {7'd0,(kernel[3][4] ~^ image[10][16])} + {7'd0,(kernel[4][0] ~^ image[11][12])} + {7'd0,(kernel[4][1] ~^ image[11][13])} + {7'd0,(kernel[4][2] ~^ image[11][14])} + {7'd0,(kernel[4][3] ~^ image[11][15])} + {7'd0,(kernel[4][4] ~^ image[11][16])};
assign out_fmap[7][13][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][13])} + {7'd0,(kernel[0][1] ~^ image[7][14])} + {7'd0,(kernel[0][2] ~^ image[7][15])} + {7'd0,(kernel[0][3] ~^ image[7][16])} + {7'd0,(kernel[0][4] ~^ image[7][17])} + {7'd0,(kernel[1][0] ~^ image[8][13])} + {7'd0,(kernel[1][1] ~^ image[8][14])} + {7'd0,(kernel[1][2] ~^ image[8][15])} + {7'd0,(kernel[1][3] ~^ image[8][16])} + {7'd0,(kernel[1][4] ~^ image[8][17])} + {7'd0,(kernel[2][0] ~^ image[9][13])} + {7'd0,(kernel[2][1] ~^ image[9][14])} + {7'd0,(kernel[2][2] ~^ image[9][15])} + {7'd0,(kernel[2][3] ~^ image[9][16])} + {7'd0,(kernel[2][4] ~^ image[9][17])} + {7'd0,(kernel[3][0] ~^ image[10][13])} + {7'd0,(kernel[3][1] ~^ image[10][14])} + {7'd0,(kernel[3][2] ~^ image[10][15])} + {7'd0,(kernel[3][3] ~^ image[10][16])} + {7'd0,(kernel[3][4] ~^ image[10][17])} + {7'd0,(kernel[4][0] ~^ image[11][13])} + {7'd0,(kernel[4][1] ~^ image[11][14])} + {7'd0,(kernel[4][2] ~^ image[11][15])} + {7'd0,(kernel[4][3] ~^ image[11][16])} + {7'd0,(kernel[4][4] ~^ image[11][17])};
assign out_fmap[7][14][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][14])} + {7'd0,(kernel[0][1] ~^ image[7][15])} + {7'd0,(kernel[0][2] ~^ image[7][16])} + {7'd0,(kernel[0][3] ~^ image[7][17])} + {7'd0,(kernel[0][4] ~^ image[7][18])} + {7'd0,(kernel[1][0] ~^ image[8][14])} + {7'd0,(kernel[1][1] ~^ image[8][15])} + {7'd0,(kernel[1][2] ~^ image[8][16])} + {7'd0,(kernel[1][3] ~^ image[8][17])} + {7'd0,(kernel[1][4] ~^ image[8][18])} + {7'd0,(kernel[2][0] ~^ image[9][14])} + {7'd0,(kernel[2][1] ~^ image[9][15])} + {7'd0,(kernel[2][2] ~^ image[9][16])} + {7'd0,(kernel[2][3] ~^ image[9][17])} + {7'd0,(kernel[2][4] ~^ image[9][18])} + {7'd0,(kernel[3][0] ~^ image[10][14])} + {7'd0,(kernel[3][1] ~^ image[10][15])} + {7'd0,(kernel[3][2] ~^ image[10][16])} + {7'd0,(kernel[3][3] ~^ image[10][17])} + {7'd0,(kernel[3][4] ~^ image[10][18])} + {7'd0,(kernel[4][0] ~^ image[11][14])} + {7'd0,(kernel[4][1] ~^ image[11][15])} + {7'd0,(kernel[4][2] ~^ image[11][16])} + {7'd0,(kernel[4][3] ~^ image[11][17])} + {7'd0,(kernel[4][4] ~^ image[11][18])};
assign out_fmap[7][15][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][15])} + {7'd0,(kernel[0][1] ~^ image[7][16])} + {7'd0,(kernel[0][2] ~^ image[7][17])} + {7'd0,(kernel[0][3] ~^ image[7][18])} + {7'd0,(kernel[0][4] ~^ image[7][19])} + {7'd0,(kernel[1][0] ~^ image[8][15])} + {7'd0,(kernel[1][1] ~^ image[8][16])} + {7'd0,(kernel[1][2] ~^ image[8][17])} + {7'd0,(kernel[1][3] ~^ image[8][18])} + {7'd0,(kernel[1][4] ~^ image[8][19])} + {7'd0,(kernel[2][0] ~^ image[9][15])} + {7'd0,(kernel[2][1] ~^ image[9][16])} + {7'd0,(kernel[2][2] ~^ image[9][17])} + {7'd0,(kernel[2][3] ~^ image[9][18])} + {7'd0,(kernel[2][4] ~^ image[9][19])} + {7'd0,(kernel[3][0] ~^ image[10][15])} + {7'd0,(kernel[3][1] ~^ image[10][16])} + {7'd0,(kernel[3][2] ~^ image[10][17])} + {7'd0,(kernel[3][3] ~^ image[10][18])} + {7'd0,(kernel[3][4] ~^ image[10][19])} + {7'd0,(kernel[4][0] ~^ image[11][15])} + {7'd0,(kernel[4][1] ~^ image[11][16])} + {7'd0,(kernel[4][2] ~^ image[11][17])} + {7'd0,(kernel[4][3] ~^ image[11][18])} + {7'd0,(kernel[4][4] ~^ image[11][19])};
assign out_fmap[7][16][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][16])} + {7'd0,(kernel[0][1] ~^ image[7][17])} + {7'd0,(kernel[0][2] ~^ image[7][18])} + {7'd0,(kernel[0][3] ~^ image[7][19])} + {7'd0,(kernel[0][4] ~^ image[7][20])} + {7'd0,(kernel[1][0] ~^ image[8][16])} + {7'd0,(kernel[1][1] ~^ image[8][17])} + {7'd0,(kernel[1][2] ~^ image[8][18])} + {7'd0,(kernel[1][3] ~^ image[8][19])} + {7'd0,(kernel[1][4] ~^ image[8][20])} + {7'd0,(kernel[2][0] ~^ image[9][16])} + {7'd0,(kernel[2][1] ~^ image[9][17])} + {7'd0,(kernel[2][2] ~^ image[9][18])} + {7'd0,(kernel[2][3] ~^ image[9][19])} + {7'd0,(kernel[2][4] ~^ image[9][20])} + {7'd0,(kernel[3][0] ~^ image[10][16])} + {7'd0,(kernel[3][1] ~^ image[10][17])} + {7'd0,(kernel[3][2] ~^ image[10][18])} + {7'd0,(kernel[3][3] ~^ image[10][19])} + {7'd0,(kernel[3][4] ~^ image[10][20])} + {7'd0,(kernel[4][0] ~^ image[11][16])} + {7'd0,(kernel[4][1] ~^ image[11][17])} + {7'd0,(kernel[4][2] ~^ image[11][18])} + {7'd0,(kernel[4][3] ~^ image[11][19])} + {7'd0,(kernel[4][4] ~^ image[11][20])};
assign out_fmap[7][17][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][17])} + {7'd0,(kernel[0][1] ~^ image[7][18])} + {7'd0,(kernel[0][2] ~^ image[7][19])} + {7'd0,(kernel[0][3] ~^ image[7][20])} + {7'd0,(kernel[0][4] ~^ image[7][21])} + {7'd0,(kernel[1][0] ~^ image[8][17])} + {7'd0,(kernel[1][1] ~^ image[8][18])} + {7'd0,(kernel[1][2] ~^ image[8][19])} + {7'd0,(kernel[1][3] ~^ image[8][20])} + {7'd0,(kernel[1][4] ~^ image[8][21])} + {7'd0,(kernel[2][0] ~^ image[9][17])} + {7'd0,(kernel[2][1] ~^ image[9][18])} + {7'd0,(kernel[2][2] ~^ image[9][19])} + {7'd0,(kernel[2][3] ~^ image[9][20])} + {7'd0,(kernel[2][4] ~^ image[9][21])} + {7'd0,(kernel[3][0] ~^ image[10][17])} + {7'd0,(kernel[3][1] ~^ image[10][18])} + {7'd0,(kernel[3][2] ~^ image[10][19])} + {7'd0,(kernel[3][3] ~^ image[10][20])} + {7'd0,(kernel[3][4] ~^ image[10][21])} + {7'd0,(kernel[4][0] ~^ image[11][17])} + {7'd0,(kernel[4][1] ~^ image[11][18])} + {7'd0,(kernel[4][2] ~^ image[11][19])} + {7'd0,(kernel[4][3] ~^ image[11][20])} + {7'd0,(kernel[4][4] ~^ image[11][21])};
assign out_fmap[7][18][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][18])} + {7'd0,(kernel[0][1] ~^ image[7][19])} + {7'd0,(kernel[0][2] ~^ image[7][20])} + {7'd0,(kernel[0][3] ~^ image[7][21])} + {7'd0,(kernel[0][4] ~^ image[7][22])} + {7'd0,(kernel[1][0] ~^ image[8][18])} + {7'd0,(kernel[1][1] ~^ image[8][19])} + {7'd0,(kernel[1][2] ~^ image[8][20])} + {7'd0,(kernel[1][3] ~^ image[8][21])} + {7'd0,(kernel[1][4] ~^ image[8][22])} + {7'd0,(kernel[2][0] ~^ image[9][18])} + {7'd0,(kernel[2][1] ~^ image[9][19])} + {7'd0,(kernel[2][2] ~^ image[9][20])} + {7'd0,(kernel[2][3] ~^ image[9][21])} + {7'd0,(kernel[2][4] ~^ image[9][22])} + {7'd0,(kernel[3][0] ~^ image[10][18])} + {7'd0,(kernel[3][1] ~^ image[10][19])} + {7'd0,(kernel[3][2] ~^ image[10][20])} + {7'd0,(kernel[3][3] ~^ image[10][21])} + {7'd0,(kernel[3][4] ~^ image[10][22])} + {7'd0,(kernel[4][0] ~^ image[11][18])} + {7'd0,(kernel[4][1] ~^ image[11][19])} + {7'd0,(kernel[4][2] ~^ image[11][20])} + {7'd0,(kernel[4][3] ~^ image[11][21])} + {7'd0,(kernel[4][4] ~^ image[11][22])};
assign out_fmap[7][19][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][19])} + {7'd0,(kernel[0][1] ~^ image[7][20])} + {7'd0,(kernel[0][2] ~^ image[7][21])} + {7'd0,(kernel[0][3] ~^ image[7][22])} + {7'd0,(kernel[0][4] ~^ image[7][23])} + {7'd0,(kernel[1][0] ~^ image[8][19])} + {7'd0,(kernel[1][1] ~^ image[8][20])} + {7'd0,(kernel[1][2] ~^ image[8][21])} + {7'd0,(kernel[1][3] ~^ image[8][22])} + {7'd0,(kernel[1][4] ~^ image[8][23])} + {7'd0,(kernel[2][0] ~^ image[9][19])} + {7'd0,(kernel[2][1] ~^ image[9][20])} + {7'd0,(kernel[2][2] ~^ image[9][21])} + {7'd0,(kernel[2][3] ~^ image[9][22])} + {7'd0,(kernel[2][4] ~^ image[9][23])} + {7'd0,(kernel[3][0] ~^ image[10][19])} + {7'd0,(kernel[3][1] ~^ image[10][20])} + {7'd0,(kernel[3][2] ~^ image[10][21])} + {7'd0,(kernel[3][3] ~^ image[10][22])} + {7'd0,(kernel[3][4] ~^ image[10][23])} + {7'd0,(kernel[4][0] ~^ image[11][19])} + {7'd0,(kernel[4][1] ~^ image[11][20])} + {7'd0,(kernel[4][2] ~^ image[11][21])} + {7'd0,(kernel[4][3] ~^ image[11][22])} + {7'd0,(kernel[4][4] ~^ image[11][23])};
assign out_fmap[7][20][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][20])} + {7'd0,(kernel[0][1] ~^ image[7][21])} + {7'd0,(kernel[0][2] ~^ image[7][22])} + {7'd0,(kernel[0][3] ~^ image[7][23])} + {7'd0,(kernel[0][4] ~^ image[7][24])} + {7'd0,(kernel[1][0] ~^ image[8][20])} + {7'd0,(kernel[1][1] ~^ image[8][21])} + {7'd0,(kernel[1][2] ~^ image[8][22])} + {7'd0,(kernel[1][3] ~^ image[8][23])} + {7'd0,(kernel[1][4] ~^ image[8][24])} + {7'd0,(kernel[2][0] ~^ image[9][20])} + {7'd0,(kernel[2][1] ~^ image[9][21])} + {7'd0,(kernel[2][2] ~^ image[9][22])} + {7'd0,(kernel[2][3] ~^ image[9][23])} + {7'd0,(kernel[2][4] ~^ image[9][24])} + {7'd0,(kernel[3][0] ~^ image[10][20])} + {7'd0,(kernel[3][1] ~^ image[10][21])} + {7'd0,(kernel[3][2] ~^ image[10][22])} + {7'd0,(kernel[3][3] ~^ image[10][23])} + {7'd0,(kernel[3][4] ~^ image[10][24])} + {7'd0,(kernel[4][0] ~^ image[11][20])} + {7'd0,(kernel[4][1] ~^ image[11][21])} + {7'd0,(kernel[4][2] ~^ image[11][22])} + {7'd0,(kernel[4][3] ~^ image[11][23])} + {7'd0,(kernel[4][4] ~^ image[11][24])};
assign out_fmap[7][21][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][21])} + {7'd0,(kernel[0][1] ~^ image[7][22])} + {7'd0,(kernel[0][2] ~^ image[7][23])} + {7'd0,(kernel[0][3] ~^ image[7][24])} + {7'd0,(kernel[0][4] ~^ image[7][25])} + {7'd0,(kernel[1][0] ~^ image[8][21])} + {7'd0,(kernel[1][1] ~^ image[8][22])} + {7'd0,(kernel[1][2] ~^ image[8][23])} + {7'd0,(kernel[1][3] ~^ image[8][24])} + {7'd0,(kernel[1][4] ~^ image[8][25])} + {7'd0,(kernel[2][0] ~^ image[9][21])} + {7'd0,(kernel[2][1] ~^ image[9][22])} + {7'd0,(kernel[2][2] ~^ image[9][23])} + {7'd0,(kernel[2][3] ~^ image[9][24])} + {7'd0,(kernel[2][4] ~^ image[9][25])} + {7'd0,(kernel[3][0] ~^ image[10][21])} + {7'd0,(kernel[3][1] ~^ image[10][22])} + {7'd0,(kernel[3][2] ~^ image[10][23])} + {7'd0,(kernel[3][3] ~^ image[10][24])} + {7'd0,(kernel[3][4] ~^ image[10][25])} + {7'd0,(kernel[4][0] ~^ image[11][21])} + {7'd0,(kernel[4][1] ~^ image[11][22])} + {7'd0,(kernel[4][2] ~^ image[11][23])} + {7'd0,(kernel[4][3] ~^ image[11][24])} + {7'd0,(kernel[4][4] ~^ image[11][25])};
assign out_fmap[7][22][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][22])} + {7'd0,(kernel[0][1] ~^ image[7][23])} + {7'd0,(kernel[0][2] ~^ image[7][24])} + {7'd0,(kernel[0][3] ~^ image[7][25])} + {7'd0,(kernel[0][4] ~^ image[7][26])} + {7'd0,(kernel[1][0] ~^ image[8][22])} + {7'd0,(kernel[1][1] ~^ image[8][23])} + {7'd0,(kernel[1][2] ~^ image[8][24])} + {7'd0,(kernel[1][3] ~^ image[8][25])} + {7'd0,(kernel[1][4] ~^ image[8][26])} + {7'd0,(kernel[2][0] ~^ image[9][22])} + {7'd0,(kernel[2][1] ~^ image[9][23])} + {7'd0,(kernel[2][2] ~^ image[9][24])} + {7'd0,(kernel[2][3] ~^ image[9][25])} + {7'd0,(kernel[2][4] ~^ image[9][26])} + {7'd0,(kernel[3][0] ~^ image[10][22])} + {7'd0,(kernel[3][1] ~^ image[10][23])} + {7'd0,(kernel[3][2] ~^ image[10][24])} + {7'd0,(kernel[3][3] ~^ image[10][25])} + {7'd0,(kernel[3][4] ~^ image[10][26])} + {7'd0,(kernel[4][0] ~^ image[11][22])} + {7'd0,(kernel[4][1] ~^ image[11][23])} + {7'd0,(kernel[4][2] ~^ image[11][24])} + {7'd0,(kernel[4][3] ~^ image[11][25])} + {7'd0,(kernel[4][4] ~^ image[11][26])};
assign out_fmap[7][23][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[7][23])} + {7'd0,(kernel[0][1] ~^ image[7][24])} + {7'd0,(kernel[0][2] ~^ image[7][25])} + {7'd0,(kernel[0][3] ~^ image[7][26])} + {7'd0,(kernel[0][4] ~^ image[7][27])} + {7'd0,(kernel[1][0] ~^ image[8][23])} + {7'd0,(kernel[1][1] ~^ image[8][24])} + {7'd0,(kernel[1][2] ~^ image[8][25])} + {7'd0,(kernel[1][3] ~^ image[8][26])} + {7'd0,(kernel[1][4] ~^ image[8][27])} + {7'd0,(kernel[2][0] ~^ image[9][23])} + {7'd0,(kernel[2][1] ~^ image[9][24])} + {7'd0,(kernel[2][2] ~^ image[9][25])} + {7'd0,(kernel[2][3] ~^ image[9][26])} + {7'd0,(kernel[2][4] ~^ image[9][27])} + {7'd0,(kernel[3][0] ~^ image[10][23])} + {7'd0,(kernel[3][1] ~^ image[10][24])} + {7'd0,(kernel[3][2] ~^ image[10][25])} + {7'd0,(kernel[3][3] ~^ image[10][26])} + {7'd0,(kernel[3][4] ~^ image[10][27])} + {7'd0,(kernel[4][0] ~^ image[11][23])} + {7'd0,(kernel[4][1] ~^ image[11][24])} + {7'd0,(kernel[4][2] ~^ image[11][25])} + {7'd0,(kernel[4][3] ~^ image[11][26])} + {7'd0,(kernel[4][4] ~^ image[11][27])};
assign out_fmap[8][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[8][0])} + {7'd0,(kernel[0][1] ~^ image[8][1])} + {7'd0,(kernel[0][2] ~^ image[8][2])} + {7'd0,(kernel[0][3] ~^ image[8][3])} + {7'd0,(kernel[0][4] ~^ image[8][4])} + {7'd0,(kernel[1][0] ~^ image[9][0])} + {7'd0,(kernel[1][1] ~^ image[9][1])} + {7'd0,(kernel[1][2] ~^ image[9][2])} + {7'd0,(kernel[1][3] ~^ image[9][3])} + {7'd0,(kernel[1][4] ~^ image[9][4])} + {7'd0,(kernel[2][0] ~^ image[10][0])} + {7'd0,(kernel[2][1] ~^ image[10][1])} + {7'd0,(kernel[2][2] ~^ image[10][2])} + {7'd0,(kernel[2][3] ~^ image[10][3])} + {7'd0,(kernel[2][4] ~^ image[10][4])} + {7'd0,(kernel[3][0] ~^ image[11][0])} + {7'd0,(kernel[3][1] ~^ image[11][1])} + {7'd0,(kernel[3][2] ~^ image[11][2])} + {7'd0,(kernel[3][3] ~^ image[11][3])} + {7'd0,(kernel[3][4] ~^ image[11][4])} + {7'd0,(kernel[4][0] ~^ image[12][0])} + {7'd0,(kernel[4][1] ~^ image[12][1])} + {7'd0,(kernel[4][2] ~^ image[12][2])} + {7'd0,(kernel[4][3] ~^ image[12][3])} + {7'd0,(kernel[4][4] ~^ image[12][4])};
assign out_fmap[8][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[8][1])} + {7'd0,(kernel[0][1] ~^ image[8][2])} + {7'd0,(kernel[0][2] ~^ image[8][3])} + {7'd0,(kernel[0][3] ~^ image[8][4])} + {7'd0,(kernel[0][4] ~^ image[8][5])} + {7'd0,(kernel[1][0] ~^ image[9][1])} + {7'd0,(kernel[1][1] ~^ image[9][2])} + {7'd0,(kernel[1][2] ~^ image[9][3])} + {7'd0,(kernel[1][3] ~^ image[9][4])} + {7'd0,(kernel[1][4] ~^ image[9][5])} + {7'd0,(kernel[2][0] ~^ image[10][1])} + {7'd0,(kernel[2][1] ~^ image[10][2])} + {7'd0,(kernel[2][2] ~^ image[10][3])} + {7'd0,(kernel[2][3] ~^ image[10][4])} + {7'd0,(kernel[2][4] ~^ image[10][5])} + {7'd0,(kernel[3][0] ~^ image[11][1])} + {7'd0,(kernel[3][1] ~^ image[11][2])} + {7'd0,(kernel[3][2] ~^ image[11][3])} + {7'd0,(kernel[3][3] ~^ image[11][4])} + {7'd0,(kernel[3][4] ~^ image[11][5])} + {7'd0,(kernel[4][0] ~^ image[12][1])} + {7'd0,(kernel[4][1] ~^ image[12][2])} + {7'd0,(kernel[4][2] ~^ image[12][3])} + {7'd0,(kernel[4][3] ~^ image[12][4])} + {7'd0,(kernel[4][4] ~^ image[12][5])};
assign out_fmap[8][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[8][2])} + {7'd0,(kernel[0][1] ~^ image[8][3])} + {7'd0,(kernel[0][2] ~^ image[8][4])} + {7'd0,(kernel[0][3] ~^ image[8][5])} + {7'd0,(kernel[0][4] ~^ image[8][6])} + {7'd0,(kernel[1][0] ~^ image[9][2])} + {7'd0,(kernel[1][1] ~^ image[9][3])} + {7'd0,(kernel[1][2] ~^ image[9][4])} + {7'd0,(kernel[1][3] ~^ image[9][5])} + {7'd0,(kernel[1][4] ~^ image[9][6])} + {7'd0,(kernel[2][0] ~^ image[10][2])} + {7'd0,(kernel[2][1] ~^ image[10][3])} + {7'd0,(kernel[2][2] ~^ image[10][4])} + {7'd0,(kernel[2][3] ~^ image[10][5])} + {7'd0,(kernel[2][4] ~^ image[10][6])} + {7'd0,(kernel[3][0] ~^ image[11][2])} + {7'd0,(kernel[3][1] ~^ image[11][3])} + {7'd0,(kernel[3][2] ~^ image[11][4])} + {7'd0,(kernel[3][3] ~^ image[11][5])} + {7'd0,(kernel[3][4] ~^ image[11][6])} + {7'd0,(kernel[4][0] ~^ image[12][2])} + {7'd0,(kernel[4][1] ~^ image[12][3])} + {7'd0,(kernel[4][2] ~^ image[12][4])} + {7'd0,(kernel[4][3] ~^ image[12][5])} + {7'd0,(kernel[4][4] ~^ image[12][6])};
assign out_fmap[8][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[8][3])} + {7'd0,(kernel[0][1] ~^ image[8][4])} + {7'd0,(kernel[0][2] ~^ image[8][5])} + {7'd0,(kernel[0][3] ~^ image[8][6])} + {7'd0,(kernel[0][4] ~^ image[8][7])} + {7'd0,(kernel[1][0] ~^ image[9][3])} + {7'd0,(kernel[1][1] ~^ image[9][4])} + {7'd0,(kernel[1][2] ~^ image[9][5])} + {7'd0,(kernel[1][3] ~^ image[9][6])} + {7'd0,(kernel[1][4] ~^ image[9][7])} + {7'd0,(kernel[2][0] ~^ image[10][3])} + {7'd0,(kernel[2][1] ~^ image[10][4])} + {7'd0,(kernel[2][2] ~^ image[10][5])} + {7'd0,(kernel[2][3] ~^ image[10][6])} + {7'd0,(kernel[2][4] ~^ image[10][7])} + {7'd0,(kernel[3][0] ~^ image[11][3])} + {7'd0,(kernel[3][1] ~^ image[11][4])} + {7'd0,(kernel[3][2] ~^ image[11][5])} + {7'd0,(kernel[3][3] ~^ image[11][6])} + {7'd0,(kernel[3][4] ~^ image[11][7])} + {7'd0,(kernel[4][0] ~^ image[12][3])} + {7'd0,(kernel[4][1] ~^ image[12][4])} + {7'd0,(kernel[4][2] ~^ image[12][5])} + {7'd0,(kernel[4][3] ~^ image[12][6])} + {7'd0,(kernel[4][4] ~^ image[12][7])};
assign out_fmap[8][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[8][4])} + {7'd0,(kernel[0][1] ~^ image[8][5])} + {7'd0,(kernel[0][2] ~^ image[8][6])} + {7'd0,(kernel[0][3] ~^ image[8][7])} + {7'd0,(kernel[0][4] ~^ image[8][8])} + {7'd0,(kernel[1][0] ~^ image[9][4])} + {7'd0,(kernel[1][1] ~^ image[9][5])} + {7'd0,(kernel[1][2] ~^ image[9][6])} + {7'd0,(kernel[1][3] ~^ image[9][7])} + {7'd0,(kernel[1][4] ~^ image[9][8])} + {7'd0,(kernel[2][0] ~^ image[10][4])} + {7'd0,(kernel[2][1] ~^ image[10][5])} + {7'd0,(kernel[2][2] ~^ image[10][6])} + {7'd0,(kernel[2][3] ~^ image[10][7])} + {7'd0,(kernel[2][4] ~^ image[10][8])} + {7'd0,(kernel[3][0] ~^ image[11][4])} + {7'd0,(kernel[3][1] ~^ image[11][5])} + {7'd0,(kernel[3][2] ~^ image[11][6])} + {7'd0,(kernel[3][3] ~^ image[11][7])} + {7'd0,(kernel[3][4] ~^ image[11][8])} + {7'd0,(kernel[4][0] ~^ image[12][4])} + {7'd0,(kernel[4][1] ~^ image[12][5])} + {7'd0,(kernel[4][2] ~^ image[12][6])} + {7'd0,(kernel[4][3] ~^ image[12][7])} + {7'd0,(kernel[4][4] ~^ image[12][8])};
assign out_fmap[8][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[8][5])} + {7'd0,(kernel[0][1] ~^ image[8][6])} + {7'd0,(kernel[0][2] ~^ image[8][7])} + {7'd0,(kernel[0][3] ~^ image[8][8])} + {7'd0,(kernel[0][4] ~^ image[8][9])} + {7'd0,(kernel[1][0] ~^ image[9][5])} + {7'd0,(kernel[1][1] ~^ image[9][6])} + {7'd0,(kernel[1][2] ~^ image[9][7])} + {7'd0,(kernel[1][3] ~^ image[9][8])} + {7'd0,(kernel[1][4] ~^ image[9][9])} + {7'd0,(kernel[2][0] ~^ image[10][5])} + {7'd0,(kernel[2][1] ~^ image[10][6])} + {7'd0,(kernel[2][2] ~^ image[10][7])} + {7'd0,(kernel[2][3] ~^ image[10][8])} + {7'd0,(kernel[2][4] ~^ image[10][9])} + {7'd0,(kernel[3][0] ~^ image[11][5])} + {7'd0,(kernel[3][1] ~^ image[11][6])} + {7'd0,(kernel[3][2] ~^ image[11][7])} + {7'd0,(kernel[3][3] ~^ image[11][8])} + {7'd0,(kernel[3][4] ~^ image[11][9])} + {7'd0,(kernel[4][0] ~^ image[12][5])} + {7'd0,(kernel[4][1] ~^ image[12][6])} + {7'd0,(kernel[4][2] ~^ image[12][7])} + {7'd0,(kernel[4][3] ~^ image[12][8])} + {7'd0,(kernel[4][4] ~^ image[12][9])};
assign out_fmap[8][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[8][6])} + {7'd0,(kernel[0][1] ~^ image[8][7])} + {7'd0,(kernel[0][2] ~^ image[8][8])} + {7'd0,(kernel[0][3] ~^ image[8][9])} + {7'd0,(kernel[0][4] ~^ image[8][10])} + {7'd0,(kernel[1][0] ~^ image[9][6])} + {7'd0,(kernel[1][1] ~^ image[9][7])} + {7'd0,(kernel[1][2] ~^ image[9][8])} + {7'd0,(kernel[1][3] ~^ image[9][9])} + {7'd0,(kernel[1][4] ~^ image[9][10])} + {7'd0,(kernel[2][0] ~^ image[10][6])} + {7'd0,(kernel[2][1] ~^ image[10][7])} + {7'd0,(kernel[2][2] ~^ image[10][8])} + {7'd0,(kernel[2][3] ~^ image[10][9])} + {7'd0,(kernel[2][4] ~^ image[10][10])} + {7'd0,(kernel[3][0] ~^ image[11][6])} + {7'd0,(kernel[3][1] ~^ image[11][7])} + {7'd0,(kernel[3][2] ~^ image[11][8])} + {7'd0,(kernel[3][3] ~^ image[11][9])} + {7'd0,(kernel[3][4] ~^ image[11][10])} + {7'd0,(kernel[4][0] ~^ image[12][6])} + {7'd0,(kernel[4][1] ~^ image[12][7])} + {7'd0,(kernel[4][2] ~^ image[12][8])} + {7'd0,(kernel[4][3] ~^ image[12][9])} + {7'd0,(kernel[4][4] ~^ image[12][10])};
assign out_fmap[8][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[8][7])} + {7'd0,(kernel[0][1] ~^ image[8][8])} + {7'd0,(kernel[0][2] ~^ image[8][9])} + {7'd0,(kernel[0][3] ~^ image[8][10])} + {7'd0,(kernel[0][4] ~^ image[8][11])} + {7'd0,(kernel[1][0] ~^ image[9][7])} + {7'd0,(kernel[1][1] ~^ image[9][8])} + {7'd0,(kernel[1][2] ~^ image[9][9])} + {7'd0,(kernel[1][3] ~^ image[9][10])} + {7'd0,(kernel[1][4] ~^ image[9][11])} + {7'd0,(kernel[2][0] ~^ image[10][7])} + {7'd0,(kernel[2][1] ~^ image[10][8])} + {7'd0,(kernel[2][2] ~^ image[10][9])} + {7'd0,(kernel[2][3] ~^ image[10][10])} + {7'd0,(kernel[2][4] ~^ image[10][11])} + {7'd0,(kernel[3][0] ~^ image[11][7])} + {7'd0,(kernel[3][1] ~^ image[11][8])} + {7'd0,(kernel[3][2] ~^ image[11][9])} + {7'd0,(kernel[3][3] ~^ image[11][10])} + {7'd0,(kernel[3][4] ~^ image[11][11])} + {7'd0,(kernel[4][0] ~^ image[12][7])} + {7'd0,(kernel[4][1] ~^ image[12][8])} + {7'd0,(kernel[4][2] ~^ image[12][9])} + {7'd0,(kernel[4][3] ~^ image[12][10])} + {7'd0,(kernel[4][4] ~^ image[12][11])};
assign out_fmap[8][8][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[8][8])} + {7'd0,(kernel[0][1] ~^ image[8][9])} + {7'd0,(kernel[0][2] ~^ image[8][10])} + {7'd0,(kernel[0][3] ~^ image[8][11])} + {7'd0,(kernel[0][4] ~^ image[8][12])} + {7'd0,(kernel[1][0] ~^ image[9][8])} + {7'd0,(kernel[1][1] ~^ image[9][9])} + {7'd0,(kernel[1][2] ~^ image[9][10])} + {7'd0,(kernel[1][3] ~^ image[9][11])} + {7'd0,(kernel[1][4] ~^ image[9][12])} + {7'd0,(kernel[2][0] ~^ image[10][8])} + {7'd0,(kernel[2][1] ~^ image[10][9])} + {7'd0,(kernel[2][2] ~^ image[10][10])} + {7'd0,(kernel[2][3] ~^ image[10][11])} + {7'd0,(kernel[2][4] ~^ image[10][12])} + {7'd0,(kernel[3][0] ~^ image[11][8])} + {7'd0,(kernel[3][1] ~^ image[11][9])} + {7'd0,(kernel[3][2] ~^ image[11][10])} + {7'd0,(kernel[3][3] ~^ image[11][11])} + {7'd0,(kernel[3][4] ~^ image[11][12])} + {7'd0,(kernel[4][0] ~^ image[12][8])} + {7'd0,(kernel[4][1] ~^ image[12][9])} + {7'd0,(kernel[4][2] ~^ image[12][10])} + {7'd0,(kernel[4][3] ~^ image[12][11])} + {7'd0,(kernel[4][4] ~^ image[12][12])};
assign out_fmap[8][9][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[8][9])} + {7'd0,(kernel[0][1] ~^ image[8][10])} + {7'd0,(kernel[0][2] ~^ image[8][11])} + {7'd0,(kernel[0][3] ~^ image[8][12])} + {7'd0,(kernel[0][4] ~^ image[8][13])} + {7'd0,(kernel[1][0] ~^ image[9][9])} + {7'd0,(kernel[1][1] ~^ image[9][10])} + {7'd0,(kernel[1][2] ~^ image[9][11])} + {7'd0,(kernel[1][3] ~^ image[9][12])} + {7'd0,(kernel[1][4] ~^ image[9][13])} + {7'd0,(kernel[2][0] ~^ image[10][9])} + {7'd0,(kernel[2][1] ~^ image[10][10])} + {7'd0,(kernel[2][2] ~^ image[10][11])} + {7'd0,(kernel[2][3] ~^ image[10][12])} + {7'd0,(kernel[2][4] ~^ image[10][13])} + {7'd0,(kernel[3][0] ~^ image[11][9])} + {7'd0,(kernel[3][1] ~^ image[11][10])} + {7'd0,(kernel[3][2] ~^ image[11][11])} + {7'd0,(kernel[3][3] ~^ image[11][12])} + {7'd0,(kernel[3][4] ~^ image[11][13])} + {7'd0,(kernel[4][0] ~^ image[12][9])} + {7'd0,(kernel[4][1] ~^ image[12][10])} + {7'd0,(kernel[4][2] ~^ image[12][11])} + {7'd0,(kernel[4][3] ~^ image[12][12])} + {7'd0,(kernel[4][4] ~^ image[12][13])};
assign out_fmap[8][10][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[8][10])} + {7'd0,(kernel[0][1] ~^ image[8][11])} + {7'd0,(kernel[0][2] ~^ image[8][12])} + {7'd0,(kernel[0][3] ~^ image[8][13])} + {7'd0,(kernel[0][4] ~^ image[8][14])} + {7'd0,(kernel[1][0] ~^ image[9][10])} + {7'd0,(kernel[1][1] ~^ image[9][11])} + {7'd0,(kernel[1][2] ~^ image[9][12])} + {7'd0,(kernel[1][3] ~^ image[9][13])} + {7'd0,(kernel[1][4] ~^ image[9][14])} + {7'd0,(kernel[2][0] ~^ image[10][10])} + {7'd0,(kernel[2][1] ~^ image[10][11])} + {7'd0,(kernel[2][2] ~^ image[10][12])} + {7'd0,(kernel[2][3] ~^ image[10][13])} + {7'd0,(kernel[2][4] ~^ image[10][14])} + {7'd0,(kernel[3][0] ~^ image[11][10])} + {7'd0,(kernel[3][1] ~^ image[11][11])} + {7'd0,(kernel[3][2] ~^ image[11][12])} + {7'd0,(kernel[3][3] ~^ image[11][13])} + {7'd0,(kernel[3][4] ~^ image[11][14])} + {7'd0,(kernel[4][0] ~^ image[12][10])} + {7'd0,(kernel[4][1] ~^ image[12][11])} + {7'd0,(kernel[4][2] ~^ image[12][12])} + {7'd0,(kernel[4][3] ~^ image[12][13])} + {7'd0,(kernel[4][4] ~^ image[12][14])};
assign out_fmap[8][11][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[8][11])} + {7'd0,(kernel[0][1] ~^ image[8][12])} + {7'd0,(kernel[0][2] ~^ image[8][13])} + {7'd0,(kernel[0][3] ~^ image[8][14])} + {7'd0,(kernel[0][4] ~^ image[8][15])} + {7'd0,(kernel[1][0] ~^ image[9][11])} + {7'd0,(kernel[1][1] ~^ image[9][12])} + {7'd0,(kernel[1][2] ~^ image[9][13])} + {7'd0,(kernel[1][3] ~^ image[9][14])} + {7'd0,(kernel[1][4] ~^ image[9][15])} + {7'd0,(kernel[2][0] ~^ image[10][11])} + {7'd0,(kernel[2][1] ~^ image[10][12])} + {7'd0,(kernel[2][2] ~^ image[10][13])} + {7'd0,(kernel[2][3] ~^ image[10][14])} + {7'd0,(kernel[2][4] ~^ image[10][15])} + {7'd0,(kernel[3][0] ~^ image[11][11])} + {7'd0,(kernel[3][1] ~^ image[11][12])} + {7'd0,(kernel[3][2] ~^ image[11][13])} + {7'd0,(kernel[3][3] ~^ image[11][14])} + {7'd0,(kernel[3][4] ~^ image[11][15])} + {7'd0,(kernel[4][0] ~^ image[12][11])} + {7'd0,(kernel[4][1] ~^ image[12][12])} + {7'd0,(kernel[4][2] ~^ image[12][13])} + {7'd0,(kernel[4][3] ~^ image[12][14])} + {7'd0,(kernel[4][4] ~^ image[12][15])};
assign out_fmap[8][12][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[8][12])} + {7'd0,(kernel[0][1] ~^ image[8][13])} + {7'd0,(kernel[0][2] ~^ image[8][14])} + {7'd0,(kernel[0][3] ~^ image[8][15])} + {7'd0,(kernel[0][4] ~^ image[8][16])} + {7'd0,(kernel[1][0] ~^ image[9][12])} + {7'd0,(kernel[1][1] ~^ image[9][13])} + {7'd0,(kernel[1][2] ~^ image[9][14])} + {7'd0,(kernel[1][3] ~^ image[9][15])} + {7'd0,(kernel[1][4] ~^ image[9][16])} + {7'd0,(kernel[2][0] ~^ image[10][12])} + {7'd0,(kernel[2][1] ~^ image[10][13])} + {7'd0,(kernel[2][2] ~^ image[10][14])} + {7'd0,(kernel[2][3] ~^ image[10][15])} + {7'd0,(kernel[2][4] ~^ image[10][16])} + {7'd0,(kernel[3][0] ~^ image[11][12])} + {7'd0,(kernel[3][1] ~^ image[11][13])} + {7'd0,(kernel[3][2] ~^ image[11][14])} + {7'd0,(kernel[3][3] ~^ image[11][15])} + {7'd0,(kernel[3][4] ~^ image[11][16])} + {7'd0,(kernel[4][0] ~^ image[12][12])} + {7'd0,(kernel[4][1] ~^ image[12][13])} + {7'd0,(kernel[4][2] ~^ image[12][14])} + {7'd0,(kernel[4][3] ~^ image[12][15])} + {7'd0,(kernel[4][4] ~^ image[12][16])};
assign out_fmap[8][13][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[8][13])} + {7'd0,(kernel[0][1] ~^ image[8][14])} + {7'd0,(kernel[0][2] ~^ image[8][15])} + {7'd0,(kernel[0][3] ~^ image[8][16])} + {7'd0,(kernel[0][4] ~^ image[8][17])} + {7'd0,(kernel[1][0] ~^ image[9][13])} + {7'd0,(kernel[1][1] ~^ image[9][14])} + {7'd0,(kernel[1][2] ~^ image[9][15])} + {7'd0,(kernel[1][3] ~^ image[9][16])} + {7'd0,(kernel[1][4] ~^ image[9][17])} + {7'd0,(kernel[2][0] ~^ image[10][13])} + {7'd0,(kernel[2][1] ~^ image[10][14])} + {7'd0,(kernel[2][2] ~^ image[10][15])} + {7'd0,(kernel[2][3] ~^ image[10][16])} + {7'd0,(kernel[2][4] ~^ image[10][17])} + {7'd0,(kernel[3][0] ~^ image[11][13])} + {7'd0,(kernel[3][1] ~^ image[11][14])} + {7'd0,(kernel[3][2] ~^ image[11][15])} + {7'd0,(kernel[3][3] ~^ image[11][16])} + {7'd0,(kernel[3][4] ~^ image[11][17])} + {7'd0,(kernel[4][0] ~^ image[12][13])} + {7'd0,(kernel[4][1] ~^ image[12][14])} + {7'd0,(kernel[4][2] ~^ image[12][15])} + {7'd0,(kernel[4][3] ~^ image[12][16])} + {7'd0,(kernel[4][4] ~^ image[12][17])};
assign out_fmap[8][14][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[8][14])} + {7'd0,(kernel[0][1] ~^ image[8][15])} + {7'd0,(kernel[0][2] ~^ image[8][16])} + {7'd0,(kernel[0][3] ~^ image[8][17])} + {7'd0,(kernel[0][4] ~^ image[8][18])} + {7'd0,(kernel[1][0] ~^ image[9][14])} + {7'd0,(kernel[1][1] ~^ image[9][15])} + {7'd0,(kernel[1][2] ~^ image[9][16])} + {7'd0,(kernel[1][3] ~^ image[9][17])} + {7'd0,(kernel[1][4] ~^ image[9][18])} + {7'd0,(kernel[2][0] ~^ image[10][14])} + {7'd0,(kernel[2][1] ~^ image[10][15])} + {7'd0,(kernel[2][2] ~^ image[10][16])} + {7'd0,(kernel[2][3] ~^ image[10][17])} + {7'd0,(kernel[2][4] ~^ image[10][18])} + {7'd0,(kernel[3][0] ~^ image[11][14])} + {7'd0,(kernel[3][1] ~^ image[11][15])} + {7'd0,(kernel[3][2] ~^ image[11][16])} + {7'd0,(kernel[3][3] ~^ image[11][17])} + {7'd0,(kernel[3][4] ~^ image[11][18])} + {7'd0,(kernel[4][0] ~^ image[12][14])} + {7'd0,(kernel[4][1] ~^ image[12][15])} + {7'd0,(kernel[4][2] ~^ image[12][16])} + {7'd0,(kernel[4][3] ~^ image[12][17])} + {7'd0,(kernel[4][4] ~^ image[12][18])};
assign out_fmap[8][15][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[8][15])} + {7'd0,(kernel[0][1] ~^ image[8][16])} + {7'd0,(kernel[0][2] ~^ image[8][17])} + {7'd0,(kernel[0][3] ~^ image[8][18])} + {7'd0,(kernel[0][4] ~^ image[8][19])} + {7'd0,(kernel[1][0] ~^ image[9][15])} + {7'd0,(kernel[1][1] ~^ image[9][16])} + {7'd0,(kernel[1][2] ~^ image[9][17])} + {7'd0,(kernel[1][3] ~^ image[9][18])} + {7'd0,(kernel[1][4] ~^ image[9][19])} + {7'd0,(kernel[2][0] ~^ image[10][15])} + {7'd0,(kernel[2][1] ~^ image[10][16])} + {7'd0,(kernel[2][2] ~^ image[10][17])} + {7'd0,(kernel[2][3] ~^ image[10][18])} + {7'd0,(kernel[2][4] ~^ image[10][19])} + {7'd0,(kernel[3][0] ~^ image[11][15])} + {7'd0,(kernel[3][1] ~^ image[11][16])} + {7'd0,(kernel[3][2] ~^ image[11][17])} + {7'd0,(kernel[3][3] ~^ image[11][18])} + {7'd0,(kernel[3][4] ~^ image[11][19])} + {7'd0,(kernel[4][0] ~^ image[12][15])} + {7'd0,(kernel[4][1] ~^ image[12][16])} + {7'd0,(kernel[4][2] ~^ image[12][17])} + {7'd0,(kernel[4][3] ~^ image[12][18])} + {7'd0,(kernel[4][4] ~^ image[12][19])};
assign out_fmap[8][16][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[8][16])} + {7'd0,(kernel[0][1] ~^ image[8][17])} + {7'd0,(kernel[0][2] ~^ image[8][18])} + {7'd0,(kernel[0][3] ~^ image[8][19])} + {7'd0,(kernel[0][4] ~^ image[8][20])} + {7'd0,(kernel[1][0] ~^ image[9][16])} + {7'd0,(kernel[1][1] ~^ image[9][17])} + {7'd0,(kernel[1][2] ~^ image[9][18])} + {7'd0,(kernel[1][3] ~^ image[9][19])} + {7'd0,(kernel[1][4] ~^ image[9][20])} + {7'd0,(kernel[2][0] ~^ image[10][16])} + {7'd0,(kernel[2][1] ~^ image[10][17])} + {7'd0,(kernel[2][2] ~^ image[10][18])} + {7'd0,(kernel[2][3] ~^ image[10][19])} + {7'd0,(kernel[2][4] ~^ image[10][20])} + {7'd0,(kernel[3][0] ~^ image[11][16])} + {7'd0,(kernel[3][1] ~^ image[11][17])} + {7'd0,(kernel[3][2] ~^ image[11][18])} + {7'd0,(kernel[3][3] ~^ image[11][19])} + {7'd0,(kernel[3][4] ~^ image[11][20])} + {7'd0,(kernel[4][0] ~^ image[12][16])} + {7'd0,(kernel[4][1] ~^ image[12][17])} + {7'd0,(kernel[4][2] ~^ image[12][18])} + {7'd0,(kernel[4][3] ~^ image[12][19])} + {7'd0,(kernel[4][4] ~^ image[12][20])};
assign out_fmap[8][17][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[8][17])} + {7'd0,(kernel[0][1] ~^ image[8][18])} + {7'd0,(kernel[0][2] ~^ image[8][19])} + {7'd0,(kernel[0][3] ~^ image[8][20])} + {7'd0,(kernel[0][4] ~^ image[8][21])} + {7'd0,(kernel[1][0] ~^ image[9][17])} + {7'd0,(kernel[1][1] ~^ image[9][18])} + {7'd0,(kernel[1][2] ~^ image[9][19])} + {7'd0,(kernel[1][3] ~^ image[9][20])} + {7'd0,(kernel[1][4] ~^ image[9][21])} + {7'd0,(kernel[2][0] ~^ image[10][17])} + {7'd0,(kernel[2][1] ~^ image[10][18])} + {7'd0,(kernel[2][2] ~^ image[10][19])} + {7'd0,(kernel[2][3] ~^ image[10][20])} + {7'd0,(kernel[2][4] ~^ image[10][21])} + {7'd0,(kernel[3][0] ~^ image[11][17])} + {7'd0,(kernel[3][1] ~^ image[11][18])} + {7'd0,(kernel[3][2] ~^ image[11][19])} + {7'd0,(kernel[3][3] ~^ image[11][20])} + {7'd0,(kernel[3][4] ~^ image[11][21])} + {7'd0,(kernel[4][0] ~^ image[12][17])} + {7'd0,(kernel[4][1] ~^ image[12][18])} + {7'd0,(kernel[4][2] ~^ image[12][19])} + {7'd0,(kernel[4][3] ~^ image[12][20])} + {7'd0,(kernel[4][4] ~^ image[12][21])};
assign out_fmap[8][18][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[8][18])} + {7'd0,(kernel[0][1] ~^ image[8][19])} + {7'd0,(kernel[0][2] ~^ image[8][20])} + {7'd0,(kernel[0][3] ~^ image[8][21])} + {7'd0,(kernel[0][4] ~^ image[8][22])} + {7'd0,(kernel[1][0] ~^ image[9][18])} + {7'd0,(kernel[1][1] ~^ image[9][19])} + {7'd0,(kernel[1][2] ~^ image[9][20])} + {7'd0,(kernel[1][3] ~^ image[9][21])} + {7'd0,(kernel[1][4] ~^ image[9][22])} + {7'd0,(kernel[2][0] ~^ image[10][18])} + {7'd0,(kernel[2][1] ~^ image[10][19])} + {7'd0,(kernel[2][2] ~^ image[10][20])} + {7'd0,(kernel[2][3] ~^ image[10][21])} + {7'd0,(kernel[2][4] ~^ image[10][22])} + {7'd0,(kernel[3][0] ~^ image[11][18])} + {7'd0,(kernel[3][1] ~^ image[11][19])} + {7'd0,(kernel[3][2] ~^ image[11][20])} + {7'd0,(kernel[3][3] ~^ image[11][21])} + {7'd0,(kernel[3][4] ~^ image[11][22])} + {7'd0,(kernel[4][0] ~^ image[12][18])} + {7'd0,(kernel[4][1] ~^ image[12][19])} + {7'd0,(kernel[4][2] ~^ image[12][20])} + {7'd0,(kernel[4][3] ~^ image[12][21])} + {7'd0,(kernel[4][4] ~^ image[12][22])};
assign out_fmap[8][19][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[8][19])} + {7'd0,(kernel[0][1] ~^ image[8][20])} + {7'd0,(kernel[0][2] ~^ image[8][21])} + {7'd0,(kernel[0][3] ~^ image[8][22])} + {7'd0,(kernel[0][4] ~^ image[8][23])} + {7'd0,(kernel[1][0] ~^ image[9][19])} + {7'd0,(kernel[1][1] ~^ image[9][20])} + {7'd0,(kernel[1][2] ~^ image[9][21])} + {7'd0,(kernel[1][3] ~^ image[9][22])} + {7'd0,(kernel[1][4] ~^ image[9][23])} + {7'd0,(kernel[2][0] ~^ image[10][19])} + {7'd0,(kernel[2][1] ~^ image[10][20])} + {7'd0,(kernel[2][2] ~^ image[10][21])} + {7'd0,(kernel[2][3] ~^ image[10][22])} + {7'd0,(kernel[2][4] ~^ image[10][23])} + {7'd0,(kernel[3][0] ~^ image[11][19])} + {7'd0,(kernel[3][1] ~^ image[11][20])} + {7'd0,(kernel[3][2] ~^ image[11][21])} + {7'd0,(kernel[3][3] ~^ image[11][22])} + {7'd0,(kernel[3][4] ~^ image[11][23])} + {7'd0,(kernel[4][0] ~^ image[12][19])} + {7'd0,(kernel[4][1] ~^ image[12][20])} + {7'd0,(kernel[4][2] ~^ image[12][21])} + {7'd0,(kernel[4][3] ~^ image[12][22])} + {7'd0,(kernel[4][4] ~^ image[12][23])};
assign out_fmap[8][20][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[8][20])} + {7'd0,(kernel[0][1] ~^ image[8][21])} + {7'd0,(kernel[0][2] ~^ image[8][22])} + {7'd0,(kernel[0][3] ~^ image[8][23])} + {7'd0,(kernel[0][4] ~^ image[8][24])} + {7'd0,(kernel[1][0] ~^ image[9][20])} + {7'd0,(kernel[1][1] ~^ image[9][21])} + {7'd0,(kernel[1][2] ~^ image[9][22])} + {7'd0,(kernel[1][3] ~^ image[9][23])} + {7'd0,(kernel[1][4] ~^ image[9][24])} + {7'd0,(kernel[2][0] ~^ image[10][20])} + {7'd0,(kernel[2][1] ~^ image[10][21])} + {7'd0,(kernel[2][2] ~^ image[10][22])} + {7'd0,(kernel[2][3] ~^ image[10][23])} + {7'd0,(kernel[2][4] ~^ image[10][24])} + {7'd0,(kernel[3][0] ~^ image[11][20])} + {7'd0,(kernel[3][1] ~^ image[11][21])} + {7'd0,(kernel[3][2] ~^ image[11][22])} + {7'd0,(kernel[3][3] ~^ image[11][23])} + {7'd0,(kernel[3][4] ~^ image[11][24])} + {7'd0,(kernel[4][0] ~^ image[12][20])} + {7'd0,(kernel[4][1] ~^ image[12][21])} + {7'd0,(kernel[4][2] ~^ image[12][22])} + {7'd0,(kernel[4][3] ~^ image[12][23])} + {7'd0,(kernel[4][4] ~^ image[12][24])};
assign out_fmap[8][21][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[8][21])} + {7'd0,(kernel[0][1] ~^ image[8][22])} + {7'd0,(kernel[0][2] ~^ image[8][23])} + {7'd0,(kernel[0][3] ~^ image[8][24])} + {7'd0,(kernel[0][4] ~^ image[8][25])} + {7'd0,(kernel[1][0] ~^ image[9][21])} + {7'd0,(kernel[1][1] ~^ image[9][22])} + {7'd0,(kernel[1][2] ~^ image[9][23])} + {7'd0,(kernel[1][3] ~^ image[9][24])} + {7'd0,(kernel[1][4] ~^ image[9][25])} + {7'd0,(kernel[2][0] ~^ image[10][21])} + {7'd0,(kernel[2][1] ~^ image[10][22])} + {7'd0,(kernel[2][2] ~^ image[10][23])} + {7'd0,(kernel[2][3] ~^ image[10][24])} + {7'd0,(kernel[2][4] ~^ image[10][25])} + {7'd0,(kernel[3][0] ~^ image[11][21])} + {7'd0,(kernel[3][1] ~^ image[11][22])} + {7'd0,(kernel[3][2] ~^ image[11][23])} + {7'd0,(kernel[3][3] ~^ image[11][24])} + {7'd0,(kernel[3][4] ~^ image[11][25])} + {7'd0,(kernel[4][0] ~^ image[12][21])} + {7'd0,(kernel[4][1] ~^ image[12][22])} + {7'd0,(kernel[4][2] ~^ image[12][23])} + {7'd0,(kernel[4][3] ~^ image[12][24])} + {7'd0,(kernel[4][4] ~^ image[12][25])};
assign out_fmap[8][22][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[8][22])} + {7'd0,(kernel[0][1] ~^ image[8][23])} + {7'd0,(kernel[0][2] ~^ image[8][24])} + {7'd0,(kernel[0][3] ~^ image[8][25])} + {7'd0,(kernel[0][4] ~^ image[8][26])} + {7'd0,(kernel[1][0] ~^ image[9][22])} + {7'd0,(kernel[1][1] ~^ image[9][23])} + {7'd0,(kernel[1][2] ~^ image[9][24])} + {7'd0,(kernel[1][3] ~^ image[9][25])} + {7'd0,(kernel[1][4] ~^ image[9][26])} + {7'd0,(kernel[2][0] ~^ image[10][22])} + {7'd0,(kernel[2][1] ~^ image[10][23])} + {7'd0,(kernel[2][2] ~^ image[10][24])} + {7'd0,(kernel[2][3] ~^ image[10][25])} + {7'd0,(kernel[2][4] ~^ image[10][26])} + {7'd0,(kernel[3][0] ~^ image[11][22])} + {7'd0,(kernel[3][1] ~^ image[11][23])} + {7'd0,(kernel[3][2] ~^ image[11][24])} + {7'd0,(kernel[3][3] ~^ image[11][25])} + {7'd0,(kernel[3][4] ~^ image[11][26])} + {7'd0,(kernel[4][0] ~^ image[12][22])} + {7'd0,(kernel[4][1] ~^ image[12][23])} + {7'd0,(kernel[4][2] ~^ image[12][24])} + {7'd0,(kernel[4][3] ~^ image[12][25])} + {7'd0,(kernel[4][4] ~^ image[12][26])};
assign out_fmap[8][23][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[8][23])} + {7'd0,(kernel[0][1] ~^ image[8][24])} + {7'd0,(kernel[0][2] ~^ image[8][25])} + {7'd0,(kernel[0][3] ~^ image[8][26])} + {7'd0,(kernel[0][4] ~^ image[8][27])} + {7'd0,(kernel[1][0] ~^ image[9][23])} + {7'd0,(kernel[1][1] ~^ image[9][24])} + {7'd0,(kernel[1][2] ~^ image[9][25])} + {7'd0,(kernel[1][3] ~^ image[9][26])} + {7'd0,(kernel[1][4] ~^ image[9][27])} + {7'd0,(kernel[2][0] ~^ image[10][23])} + {7'd0,(kernel[2][1] ~^ image[10][24])} + {7'd0,(kernel[2][2] ~^ image[10][25])} + {7'd0,(kernel[2][3] ~^ image[10][26])} + {7'd0,(kernel[2][4] ~^ image[10][27])} + {7'd0,(kernel[3][0] ~^ image[11][23])} + {7'd0,(kernel[3][1] ~^ image[11][24])} + {7'd0,(kernel[3][2] ~^ image[11][25])} + {7'd0,(kernel[3][3] ~^ image[11][26])} + {7'd0,(kernel[3][4] ~^ image[11][27])} + {7'd0,(kernel[4][0] ~^ image[12][23])} + {7'd0,(kernel[4][1] ~^ image[12][24])} + {7'd0,(kernel[4][2] ~^ image[12][25])} + {7'd0,(kernel[4][3] ~^ image[12][26])} + {7'd0,(kernel[4][4] ~^ image[12][27])};
assign out_fmap[9][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[9][0])} + {7'd0,(kernel[0][1] ~^ image[9][1])} + {7'd0,(kernel[0][2] ~^ image[9][2])} + {7'd0,(kernel[0][3] ~^ image[9][3])} + {7'd0,(kernel[0][4] ~^ image[9][4])} + {7'd0,(kernel[1][0] ~^ image[10][0])} + {7'd0,(kernel[1][1] ~^ image[10][1])} + {7'd0,(kernel[1][2] ~^ image[10][2])} + {7'd0,(kernel[1][3] ~^ image[10][3])} + {7'd0,(kernel[1][4] ~^ image[10][4])} + {7'd0,(kernel[2][0] ~^ image[11][0])} + {7'd0,(kernel[2][1] ~^ image[11][1])} + {7'd0,(kernel[2][2] ~^ image[11][2])} + {7'd0,(kernel[2][3] ~^ image[11][3])} + {7'd0,(kernel[2][4] ~^ image[11][4])} + {7'd0,(kernel[3][0] ~^ image[12][0])} + {7'd0,(kernel[3][1] ~^ image[12][1])} + {7'd0,(kernel[3][2] ~^ image[12][2])} + {7'd0,(kernel[3][3] ~^ image[12][3])} + {7'd0,(kernel[3][4] ~^ image[12][4])} + {7'd0,(kernel[4][0] ~^ image[13][0])} + {7'd0,(kernel[4][1] ~^ image[13][1])} + {7'd0,(kernel[4][2] ~^ image[13][2])} + {7'd0,(kernel[4][3] ~^ image[13][3])} + {7'd0,(kernel[4][4] ~^ image[13][4])};
assign out_fmap[9][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[9][1])} + {7'd0,(kernel[0][1] ~^ image[9][2])} + {7'd0,(kernel[0][2] ~^ image[9][3])} + {7'd0,(kernel[0][3] ~^ image[9][4])} + {7'd0,(kernel[0][4] ~^ image[9][5])} + {7'd0,(kernel[1][0] ~^ image[10][1])} + {7'd0,(kernel[1][1] ~^ image[10][2])} + {7'd0,(kernel[1][2] ~^ image[10][3])} + {7'd0,(kernel[1][3] ~^ image[10][4])} + {7'd0,(kernel[1][4] ~^ image[10][5])} + {7'd0,(kernel[2][0] ~^ image[11][1])} + {7'd0,(kernel[2][1] ~^ image[11][2])} + {7'd0,(kernel[2][2] ~^ image[11][3])} + {7'd0,(kernel[2][3] ~^ image[11][4])} + {7'd0,(kernel[2][4] ~^ image[11][5])} + {7'd0,(kernel[3][0] ~^ image[12][1])} + {7'd0,(kernel[3][1] ~^ image[12][2])} + {7'd0,(kernel[3][2] ~^ image[12][3])} + {7'd0,(kernel[3][3] ~^ image[12][4])} + {7'd0,(kernel[3][4] ~^ image[12][5])} + {7'd0,(kernel[4][0] ~^ image[13][1])} + {7'd0,(kernel[4][1] ~^ image[13][2])} + {7'd0,(kernel[4][2] ~^ image[13][3])} + {7'd0,(kernel[4][3] ~^ image[13][4])} + {7'd0,(kernel[4][4] ~^ image[13][5])};
assign out_fmap[9][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[9][2])} + {7'd0,(kernel[0][1] ~^ image[9][3])} + {7'd0,(kernel[0][2] ~^ image[9][4])} + {7'd0,(kernel[0][3] ~^ image[9][5])} + {7'd0,(kernel[0][4] ~^ image[9][6])} + {7'd0,(kernel[1][0] ~^ image[10][2])} + {7'd0,(kernel[1][1] ~^ image[10][3])} + {7'd0,(kernel[1][2] ~^ image[10][4])} + {7'd0,(kernel[1][3] ~^ image[10][5])} + {7'd0,(kernel[1][4] ~^ image[10][6])} + {7'd0,(kernel[2][0] ~^ image[11][2])} + {7'd0,(kernel[2][1] ~^ image[11][3])} + {7'd0,(kernel[2][2] ~^ image[11][4])} + {7'd0,(kernel[2][3] ~^ image[11][5])} + {7'd0,(kernel[2][4] ~^ image[11][6])} + {7'd0,(kernel[3][0] ~^ image[12][2])} + {7'd0,(kernel[3][1] ~^ image[12][3])} + {7'd0,(kernel[3][2] ~^ image[12][4])} + {7'd0,(kernel[3][3] ~^ image[12][5])} + {7'd0,(kernel[3][4] ~^ image[12][6])} + {7'd0,(kernel[4][0] ~^ image[13][2])} + {7'd0,(kernel[4][1] ~^ image[13][3])} + {7'd0,(kernel[4][2] ~^ image[13][4])} + {7'd0,(kernel[4][3] ~^ image[13][5])} + {7'd0,(kernel[4][4] ~^ image[13][6])};
assign out_fmap[9][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[9][3])} + {7'd0,(kernel[0][1] ~^ image[9][4])} + {7'd0,(kernel[0][2] ~^ image[9][5])} + {7'd0,(kernel[0][3] ~^ image[9][6])} + {7'd0,(kernel[0][4] ~^ image[9][7])} + {7'd0,(kernel[1][0] ~^ image[10][3])} + {7'd0,(kernel[1][1] ~^ image[10][4])} + {7'd0,(kernel[1][2] ~^ image[10][5])} + {7'd0,(kernel[1][3] ~^ image[10][6])} + {7'd0,(kernel[1][4] ~^ image[10][7])} + {7'd0,(kernel[2][0] ~^ image[11][3])} + {7'd0,(kernel[2][1] ~^ image[11][4])} + {7'd0,(kernel[2][2] ~^ image[11][5])} + {7'd0,(kernel[2][3] ~^ image[11][6])} + {7'd0,(kernel[2][4] ~^ image[11][7])} + {7'd0,(kernel[3][0] ~^ image[12][3])} + {7'd0,(kernel[3][1] ~^ image[12][4])} + {7'd0,(kernel[3][2] ~^ image[12][5])} + {7'd0,(kernel[3][3] ~^ image[12][6])} + {7'd0,(kernel[3][4] ~^ image[12][7])} + {7'd0,(kernel[4][0] ~^ image[13][3])} + {7'd0,(kernel[4][1] ~^ image[13][4])} + {7'd0,(kernel[4][2] ~^ image[13][5])} + {7'd0,(kernel[4][3] ~^ image[13][6])} + {7'd0,(kernel[4][4] ~^ image[13][7])};
assign out_fmap[9][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[9][4])} + {7'd0,(kernel[0][1] ~^ image[9][5])} + {7'd0,(kernel[0][2] ~^ image[9][6])} + {7'd0,(kernel[0][3] ~^ image[9][7])} + {7'd0,(kernel[0][4] ~^ image[9][8])} + {7'd0,(kernel[1][0] ~^ image[10][4])} + {7'd0,(kernel[1][1] ~^ image[10][5])} + {7'd0,(kernel[1][2] ~^ image[10][6])} + {7'd0,(kernel[1][3] ~^ image[10][7])} + {7'd0,(kernel[1][4] ~^ image[10][8])} + {7'd0,(kernel[2][0] ~^ image[11][4])} + {7'd0,(kernel[2][1] ~^ image[11][5])} + {7'd0,(kernel[2][2] ~^ image[11][6])} + {7'd0,(kernel[2][3] ~^ image[11][7])} + {7'd0,(kernel[2][4] ~^ image[11][8])} + {7'd0,(kernel[3][0] ~^ image[12][4])} + {7'd0,(kernel[3][1] ~^ image[12][5])} + {7'd0,(kernel[3][2] ~^ image[12][6])} + {7'd0,(kernel[3][3] ~^ image[12][7])} + {7'd0,(kernel[3][4] ~^ image[12][8])} + {7'd0,(kernel[4][0] ~^ image[13][4])} + {7'd0,(kernel[4][1] ~^ image[13][5])} + {7'd0,(kernel[4][2] ~^ image[13][6])} + {7'd0,(kernel[4][3] ~^ image[13][7])} + {7'd0,(kernel[4][4] ~^ image[13][8])};
assign out_fmap[9][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[9][5])} + {7'd0,(kernel[0][1] ~^ image[9][6])} + {7'd0,(kernel[0][2] ~^ image[9][7])} + {7'd0,(kernel[0][3] ~^ image[9][8])} + {7'd0,(kernel[0][4] ~^ image[9][9])} + {7'd0,(kernel[1][0] ~^ image[10][5])} + {7'd0,(kernel[1][1] ~^ image[10][6])} + {7'd0,(kernel[1][2] ~^ image[10][7])} + {7'd0,(kernel[1][3] ~^ image[10][8])} + {7'd0,(kernel[1][4] ~^ image[10][9])} + {7'd0,(kernel[2][0] ~^ image[11][5])} + {7'd0,(kernel[2][1] ~^ image[11][6])} + {7'd0,(kernel[2][2] ~^ image[11][7])} + {7'd0,(kernel[2][3] ~^ image[11][8])} + {7'd0,(kernel[2][4] ~^ image[11][9])} + {7'd0,(kernel[3][0] ~^ image[12][5])} + {7'd0,(kernel[3][1] ~^ image[12][6])} + {7'd0,(kernel[3][2] ~^ image[12][7])} + {7'd0,(kernel[3][3] ~^ image[12][8])} + {7'd0,(kernel[3][4] ~^ image[12][9])} + {7'd0,(kernel[4][0] ~^ image[13][5])} + {7'd0,(kernel[4][1] ~^ image[13][6])} + {7'd0,(kernel[4][2] ~^ image[13][7])} + {7'd0,(kernel[4][3] ~^ image[13][8])} + {7'd0,(kernel[4][4] ~^ image[13][9])};
assign out_fmap[9][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[9][6])} + {7'd0,(kernel[0][1] ~^ image[9][7])} + {7'd0,(kernel[0][2] ~^ image[9][8])} + {7'd0,(kernel[0][3] ~^ image[9][9])} + {7'd0,(kernel[0][4] ~^ image[9][10])} + {7'd0,(kernel[1][0] ~^ image[10][6])} + {7'd0,(kernel[1][1] ~^ image[10][7])} + {7'd0,(kernel[1][2] ~^ image[10][8])} + {7'd0,(kernel[1][3] ~^ image[10][9])} + {7'd0,(kernel[1][4] ~^ image[10][10])} + {7'd0,(kernel[2][0] ~^ image[11][6])} + {7'd0,(kernel[2][1] ~^ image[11][7])} + {7'd0,(kernel[2][2] ~^ image[11][8])} + {7'd0,(kernel[2][3] ~^ image[11][9])} + {7'd0,(kernel[2][4] ~^ image[11][10])} + {7'd0,(kernel[3][0] ~^ image[12][6])} + {7'd0,(kernel[3][1] ~^ image[12][7])} + {7'd0,(kernel[3][2] ~^ image[12][8])} + {7'd0,(kernel[3][3] ~^ image[12][9])} + {7'd0,(kernel[3][4] ~^ image[12][10])} + {7'd0,(kernel[4][0] ~^ image[13][6])} + {7'd0,(kernel[4][1] ~^ image[13][7])} + {7'd0,(kernel[4][2] ~^ image[13][8])} + {7'd0,(kernel[4][3] ~^ image[13][9])} + {7'd0,(kernel[4][4] ~^ image[13][10])};
assign out_fmap[9][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[9][7])} + {7'd0,(kernel[0][1] ~^ image[9][8])} + {7'd0,(kernel[0][2] ~^ image[9][9])} + {7'd0,(kernel[0][3] ~^ image[9][10])} + {7'd0,(kernel[0][4] ~^ image[9][11])} + {7'd0,(kernel[1][0] ~^ image[10][7])} + {7'd0,(kernel[1][1] ~^ image[10][8])} + {7'd0,(kernel[1][2] ~^ image[10][9])} + {7'd0,(kernel[1][3] ~^ image[10][10])} + {7'd0,(kernel[1][4] ~^ image[10][11])} + {7'd0,(kernel[2][0] ~^ image[11][7])} + {7'd0,(kernel[2][1] ~^ image[11][8])} + {7'd0,(kernel[2][2] ~^ image[11][9])} + {7'd0,(kernel[2][3] ~^ image[11][10])} + {7'd0,(kernel[2][4] ~^ image[11][11])} + {7'd0,(kernel[3][0] ~^ image[12][7])} + {7'd0,(kernel[3][1] ~^ image[12][8])} + {7'd0,(kernel[3][2] ~^ image[12][9])} + {7'd0,(kernel[3][3] ~^ image[12][10])} + {7'd0,(kernel[3][4] ~^ image[12][11])} + {7'd0,(kernel[4][0] ~^ image[13][7])} + {7'd0,(kernel[4][1] ~^ image[13][8])} + {7'd0,(kernel[4][2] ~^ image[13][9])} + {7'd0,(kernel[4][3] ~^ image[13][10])} + {7'd0,(kernel[4][4] ~^ image[13][11])};
assign out_fmap[9][8][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[9][8])} + {7'd0,(kernel[0][1] ~^ image[9][9])} + {7'd0,(kernel[0][2] ~^ image[9][10])} + {7'd0,(kernel[0][3] ~^ image[9][11])} + {7'd0,(kernel[0][4] ~^ image[9][12])} + {7'd0,(kernel[1][0] ~^ image[10][8])} + {7'd0,(kernel[1][1] ~^ image[10][9])} + {7'd0,(kernel[1][2] ~^ image[10][10])} + {7'd0,(kernel[1][3] ~^ image[10][11])} + {7'd0,(kernel[1][4] ~^ image[10][12])} + {7'd0,(kernel[2][0] ~^ image[11][8])} + {7'd0,(kernel[2][1] ~^ image[11][9])} + {7'd0,(kernel[2][2] ~^ image[11][10])} + {7'd0,(kernel[2][3] ~^ image[11][11])} + {7'd0,(kernel[2][4] ~^ image[11][12])} + {7'd0,(kernel[3][0] ~^ image[12][8])} + {7'd0,(kernel[3][1] ~^ image[12][9])} + {7'd0,(kernel[3][2] ~^ image[12][10])} + {7'd0,(kernel[3][3] ~^ image[12][11])} + {7'd0,(kernel[3][4] ~^ image[12][12])} + {7'd0,(kernel[4][0] ~^ image[13][8])} + {7'd0,(kernel[4][1] ~^ image[13][9])} + {7'd0,(kernel[4][2] ~^ image[13][10])} + {7'd0,(kernel[4][3] ~^ image[13][11])} + {7'd0,(kernel[4][4] ~^ image[13][12])};
assign out_fmap[9][9][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[9][9])} + {7'd0,(kernel[0][1] ~^ image[9][10])} + {7'd0,(kernel[0][2] ~^ image[9][11])} + {7'd0,(kernel[0][3] ~^ image[9][12])} + {7'd0,(kernel[0][4] ~^ image[9][13])} + {7'd0,(kernel[1][0] ~^ image[10][9])} + {7'd0,(kernel[1][1] ~^ image[10][10])} + {7'd0,(kernel[1][2] ~^ image[10][11])} + {7'd0,(kernel[1][3] ~^ image[10][12])} + {7'd0,(kernel[1][4] ~^ image[10][13])} + {7'd0,(kernel[2][0] ~^ image[11][9])} + {7'd0,(kernel[2][1] ~^ image[11][10])} + {7'd0,(kernel[2][2] ~^ image[11][11])} + {7'd0,(kernel[2][3] ~^ image[11][12])} + {7'd0,(kernel[2][4] ~^ image[11][13])} + {7'd0,(kernel[3][0] ~^ image[12][9])} + {7'd0,(kernel[3][1] ~^ image[12][10])} + {7'd0,(kernel[3][2] ~^ image[12][11])} + {7'd0,(kernel[3][3] ~^ image[12][12])} + {7'd0,(kernel[3][4] ~^ image[12][13])} + {7'd0,(kernel[4][0] ~^ image[13][9])} + {7'd0,(kernel[4][1] ~^ image[13][10])} + {7'd0,(kernel[4][2] ~^ image[13][11])} + {7'd0,(kernel[4][3] ~^ image[13][12])} + {7'd0,(kernel[4][4] ~^ image[13][13])};
assign out_fmap[9][10][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[9][10])} + {7'd0,(kernel[0][1] ~^ image[9][11])} + {7'd0,(kernel[0][2] ~^ image[9][12])} + {7'd0,(kernel[0][3] ~^ image[9][13])} + {7'd0,(kernel[0][4] ~^ image[9][14])} + {7'd0,(kernel[1][0] ~^ image[10][10])} + {7'd0,(kernel[1][1] ~^ image[10][11])} + {7'd0,(kernel[1][2] ~^ image[10][12])} + {7'd0,(kernel[1][3] ~^ image[10][13])} + {7'd0,(kernel[1][4] ~^ image[10][14])} + {7'd0,(kernel[2][0] ~^ image[11][10])} + {7'd0,(kernel[2][1] ~^ image[11][11])} + {7'd0,(kernel[2][2] ~^ image[11][12])} + {7'd0,(kernel[2][3] ~^ image[11][13])} + {7'd0,(kernel[2][4] ~^ image[11][14])} + {7'd0,(kernel[3][0] ~^ image[12][10])} + {7'd0,(kernel[3][1] ~^ image[12][11])} + {7'd0,(kernel[3][2] ~^ image[12][12])} + {7'd0,(kernel[3][3] ~^ image[12][13])} + {7'd0,(kernel[3][4] ~^ image[12][14])} + {7'd0,(kernel[4][0] ~^ image[13][10])} + {7'd0,(kernel[4][1] ~^ image[13][11])} + {7'd0,(kernel[4][2] ~^ image[13][12])} + {7'd0,(kernel[4][3] ~^ image[13][13])} + {7'd0,(kernel[4][4] ~^ image[13][14])};
assign out_fmap[9][11][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[9][11])} + {7'd0,(kernel[0][1] ~^ image[9][12])} + {7'd0,(kernel[0][2] ~^ image[9][13])} + {7'd0,(kernel[0][3] ~^ image[9][14])} + {7'd0,(kernel[0][4] ~^ image[9][15])} + {7'd0,(kernel[1][0] ~^ image[10][11])} + {7'd0,(kernel[1][1] ~^ image[10][12])} + {7'd0,(kernel[1][2] ~^ image[10][13])} + {7'd0,(kernel[1][3] ~^ image[10][14])} + {7'd0,(kernel[1][4] ~^ image[10][15])} + {7'd0,(kernel[2][0] ~^ image[11][11])} + {7'd0,(kernel[2][1] ~^ image[11][12])} + {7'd0,(kernel[2][2] ~^ image[11][13])} + {7'd0,(kernel[2][3] ~^ image[11][14])} + {7'd0,(kernel[2][4] ~^ image[11][15])} + {7'd0,(kernel[3][0] ~^ image[12][11])} + {7'd0,(kernel[3][1] ~^ image[12][12])} + {7'd0,(kernel[3][2] ~^ image[12][13])} + {7'd0,(kernel[3][3] ~^ image[12][14])} + {7'd0,(kernel[3][4] ~^ image[12][15])} + {7'd0,(kernel[4][0] ~^ image[13][11])} + {7'd0,(kernel[4][1] ~^ image[13][12])} + {7'd0,(kernel[4][2] ~^ image[13][13])} + {7'd0,(kernel[4][3] ~^ image[13][14])} + {7'd0,(kernel[4][4] ~^ image[13][15])};
assign out_fmap[9][12][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[9][12])} + {7'd0,(kernel[0][1] ~^ image[9][13])} + {7'd0,(kernel[0][2] ~^ image[9][14])} + {7'd0,(kernel[0][3] ~^ image[9][15])} + {7'd0,(kernel[0][4] ~^ image[9][16])} + {7'd0,(kernel[1][0] ~^ image[10][12])} + {7'd0,(kernel[1][1] ~^ image[10][13])} + {7'd0,(kernel[1][2] ~^ image[10][14])} + {7'd0,(kernel[1][3] ~^ image[10][15])} + {7'd0,(kernel[1][4] ~^ image[10][16])} + {7'd0,(kernel[2][0] ~^ image[11][12])} + {7'd0,(kernel[2][1] ~^ image[11][13])} + {7'd0,(kernel[2][2] ~^ image[11][14])} + {7'd0,(kernel[2][3] ~^ image[11][15])} + {7'd0,(kernel[2][4] ~^ image[11][16])} + {7'd0,(kernel[3][0] ~^ image[12][12])} + {7'd0,(kernel[3][1] ~^ image[12][13])} + {7'd0,(kernel[3][2] ~^ image[12][14])} + {7'd0,(kernel[3][3] ~^ image[12][15])} + {7'd0,(kernel[3][4] ~^ image[12][16])} + {7'd0,(kernel[4][0] ~^ image[13][12])} + {7'd0,(kernel[4][1] ~^ image[13][13])} + {7'd0,(kernel[4][2] ~^ image[13][14])} + {7'd0,(kernel[4][3] ~^ image[13][15])} + {7'd0,(kernel[4][4] ~^ image[13][16])};
assign out_fmap[9][13][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[9][13])} + {7'd0,(kernel[0][1] ~^ image[9][14])} + {7'd0,(kernel[0][2] ~^ image[9][15])} + {7'd0,(kernel[0][3] ~^ image[9][16])} + {7'd0,(kernel[0][4] ~^ image[9][17])} + {7'd0,(kernel[1][0] ~^ image[10][13])} + {7'd0,(kernel[1][1] ~^ image[10][14])} + {7'd0,(kernel[1][2] ~^ image[10][15])} + {7'd0,(kernel[1][3] ~^ image[10][16])} + {7'd0,(kernel[1][4] ~^ image[10][17])} + {7'd0,(kernel[2][0] ~^ image[11][13])} + {7'd0,(kernel[2][1] ~^ image[11][14])} + {7'd0,(kernel[2][2] ~^ image[11][15])} + {7'd0,(kernel[2][3] ~^ image[11][16])} + {7'd0,(kernel[2][4] ~^ image[11][17])} + {7'd0,(kernel[3][0] ~^ image[12][13])} + {7'd0,(kernel[3][1] ~^ image[12][14])} + {7'd0,(kernel[3][2] ~^ image[12][15])} + {7'd0,(kernel[3][3] ~^ image[12][16])} + {7'd0,(kernel[3][4] ~^ image[12][17])} + {7'd0,(kernel[4][0] ~^ image[13][13])} + {7'd0,(kernel[4][1] ~^ image[13][14])} + {7'd0,(kernel[4][2] ~^ image[13][15])} + {7'd0,(kernel[4][3] ~^ image[13][16])} + {7'd0,(kernel[4][4] ~^ image[13][17])};
assign out_fmap[9][14][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[9][14])} + {7'd0,(kernel[0][1] ~^ image[9][15])} + {7'd0,(kernel[0][2] ~^ image[9][16])} + {7'd0,(kernel[0][3] ~^ image[9][17])} + {7'd0,(kernel[0][4] ~^ image[9][18])} + {7'd0,(kernel[1][0] ~^ image[10][14])} + {7'd0,(kernel[1][1] ~^ image[10][15])} + {7'd0,(kernel[1][2] ~^ image[10][16])} + {7'd0,(kernel[1][3] ~^ image[10][17])} + {7'd0,(kernel[1][4] ~^ image[10][18])} + {7'd0,(kernel[2][0] ~^ image[11][14])} + {7'd0,(kernel[2][1] ~^ image[11][15])} + {7'd0,(kernel[2][2] ~^ image[11][16])} + {7'd0,(kernel[2][3] ~^ image[11][17])} + {7'd0,(kernel[2][4] ~^ image[11][18])} + {7'd0,(kernel[3][0] ~^ image[12][14])} + {7'd0,(kernel[3][1] ~^ image[12][15])} + {7'd0,(kernel[3][2] ~^ image[12][16])} + {7'd0,(kernel[3][3] ~^ image[12][17])} + {7'd0,(kernel[3][4] ~^ image[12][18])} + {7'd0,(kernel[4][0] ~^ image[13][14])} + {7'd0,(kernel[4][1] ~^ image[13][15])} + {7'd0,(kernel[4][2] ~^ image[13][16])} + {7'd0,(kernel[4][3] ~^ image[13][17])} + {7'd0,(kernel[4][4] ~^ image[13][18])};
assign out_fmap[9][15][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[9][15])} + {7'd0,(kernel[0][1] ~^ image[9][16])} + {7'd0,(kernel[0][2] ~^ image[9][17])} + {7'd0,(kernel[0][3] ~^ image[9][18])} + {7'd0,(kernel[0][4] ~^ image[9][19])} + {7'd0,(kernel[1][0] ~^ image[10][15])} + {7'd0,(kernel[1][1] ~^ image[10][16])} + {7'd0,(kernel[1][2] ~^ image[10][17])} + {7'd0,(kernel[1][3] ~^ image[10][18])} + {7'd0,(kernel[1][4] ~^ image[10][19])} + {7'd0,(kernel[2][0] ~^ image[11][15])} + {7'd0,(kernel[2][1] ~^ image[11][16])} + {7'd0,(kernel[2][2] ~^ image[11][17])} + {7'd0,(kernel[2][3] ~^ image[11][18])} + {7'd0,(kernel[2][4] ~^ image[11][19])} + {7'd0,(kernel[3][0] ~^ image[12][15])} + {7'd0,(kernel[3][1] ~^ image[12][16])} + {7'd0,(kernel[3][2] ~^ image[12][17])} + {7'd0,(kernel[3][3] ~^ image[12][18])} + {7'd0,(kernel[3][4] ~^ image[12][19])} + {7'd0,(kernel[4][0] ~^ image[13][15])} + {7'd0,(kernel[4][1] ~^ image[13][16])} + {7'd0,(kernel[4][2] ~^ image[13][17])} + {7'd0,(kernel[4][3] ~^ image[13][18])} + {7'd0,(kernel[4][4] ~^ image[13][19])};
assign out_fmap[9][16][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[9][16])} + {7'd0,(kernel[0][1] ~^ image[9][17])} + {7'd0,(kernel[0][2] ~^ image[9][18])} + {7'd0,(kernel[0][3] ~^ image[9][19])} + {7'd0,(kernel[0][4] ~^ image[9][20])} + {7'd0,(kernel[1][0] ~^ image[10][16])} + {7'd0,(kernel[1][1] ~^ image[10][17])} + {7'd0,(kernel[1][2] ~^ image[10][18])} + {7'd0,(kernel[1][3] ~^ image[10][19])} + {7'd0,(kernel[1][4] ~^ image[10][20])} + {7'd0,(kernel[2][0] ~^ image[11][16])} + {7'd0,(kernel[2][1] ~^ image[11][17])} + {7'd0,(kernel[2][2] ~^ image[11][18])} + {7'd0,(kernel[2][3] ~^ image[11][19])} + {7'd0,(kernel[2][4] ~^ image[11][20])} + {7'd0,(kernel[3][0] ~^ image[12][16])} + {7'd0,(kernel[3][1] ~^ image[12][17])} + {7'd0,(kernel[3][2] ~^ image[12][18])} + {7'd0,(kernel[3][3] ~^ image[12][19])} + {7'd0,(kernel[3][4] ~^ image[12][20])} + {7'd0,(kernel[4][0] ~^ image[13][16])} + {7'd0,(kernel[4][1] ~^ image[13][17])} + {7'd0,(kernel[4][2] ~^ image[13][18])} + {7'd0,(kernel[4][3] ~^ image[13][19])} + {7'd0,(kernel[4][4] ~^ image[13][20])};
assign out_fmap[9][17][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[9][17])} + {7'd0,(kernel[0][1] ~^ image[9][18])} + {7'd0,(kernel[0][2] ~^ image[9][19])} + {7'd0,(kernel[0][3] ~^ image[9][20])} + {7'd0,(kernel[0][4] ~^ image[9][21])} + {7'd0,(kernel[1][0] ~^ image[10][17])} + {7'd0,(kernel[1][1] ~^ image[10][18])} + {7'd0,(kernel[1][2] ~^ image[10][19])} + {7'd0,(kernel[1][3] ~^ image[10][20])} + {7'd0,(kernel[1][4] ~^ image[10][21])} + {7'd0,(kernel[2][0] ~^ image[11][17])} + {7'd0,(kernel[2][1] ~^ image[11][18])} + {7'd0,(kernel[2][2] ~^ image[11][19])} + {7'd0,(kernel[2][3] ~^ image[11][20])} + {7'd0,(kernel[2][4] ~^ image[11][21])} + {7'd0,(kernel[3][0] ~^ image[12][17])} + {7'd0,(kernel[3][1] ~^ image[12][18])} + {7'd0,(kernel[3][2] ~^ image[12][19])} + {7'd0,(kernel[3][3] ~^ image[12][20])} + {7'd0,(kernel[3][4] ~^ image[12][21])} + {7'd0,(kernel[4][0] ~^ image[13][17])} + {7'd0,(kernel[4][1] ~^ image[13][18])} + {7'd0,(kernel[4][2] ~^ image[13][19])} + {7'd0,(kernel[4][3] ~^ image[13][20])} + {7'd0,(kernel[4][4] ~^ image[13][21])};
assign out_fmap[9][18][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[9][18])} + {7'd0,(kernel[0][1] ~^ image[9][19])} + {7'd0,(kernel[0][2] ~^ image[9][20])} + {7'd0,(kernel[0][3] ~^ image[9][21])} + {7'd0,(kernel[0][4] ~^ image[9][22])} + {7'd0,(kernel[1][0] ~^ image[10][18])} + {7'd0,(kernel[1][1] ~^ image[10][19])} + {7'd0,(kernel[1][2] ~^ image[10][20])} + {7'd0,(kernel[1][3] ~^ image[10][21])} + {7'd0,(kernel[1][4] ~^ image[10][22])} + {7'd0,(kernel[2][0] ~^ image[11][18])} + {7'd0,(kernel[2][1] ~^ image[11][19])} + {7'd0,(kernel[2][2] ~^ image[11][20])} + {7'd0,(kernel[2][3] ~^ image[11][21])} + {7'd0,(kernel[2][4] ~^ image[11][22])} + {7'd0,(kernel[3][0] ~^ image[12][18])} + {7'd0,(kernel[3][1] ~^ image[12][19])} + {7'd0,(kernel[3][2] ~^ image[12][20])} + {7'd0,(kernel[3][3] ~^ image[12][21])} + {7'd0,(kernel[3][4] ~^ image[12][22])} + {7'd0,(kernel[4][0] ~^ image[13][18])} + {7'd0,(kernel[4][1] ~^ image[13][19])} + {7'd0,(kernel[4][2] ~^ image[13][20])} + {7'd0,(kernel[4][3] ~^ image[13][21])} + {7'd0,(kernel[4][4] ~^ image[13][22])};
assign out_fmap[9][19][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[9][19])} + {7'd0,(kernel[0][1] ~^ image[9][20])} + {7'd0,(kernel[0][2] ~^ image[9][21])} + {7'd0,(kernel[0][3] ~^ image[9][22])} + {7'd0,(kernel[0][4] ~^ image[9][23])} + {7'd0,(kernel[1][0] ~^ image[10][19])} + {7'd0,(kernel[1][1] ~^ image[10][20])} + {7'd0,(kernel[1][2] ~^ image[10][21])} + {7'd0,(kernel[1][3] ~^ image[10][22])} + {7'd0,(kernel[1][4] ~^ image[10][23])} + {7'd0,(kernel[2][0] ~^ image[11][19])} + {7'd0,(kernel[2][1] ~^ image[11][20])} + {7'd0,(kernel[2][2] ~^ image[11][21])} + {7'd0,(kernel[2][3] ~^ image[11][22])} + {7'd0,(kernel[2][4] ~^ image[11][23])} + {7'd0,(kernel[3][0] ~^ image[12][19])} + {7'd0,(kernel[3][1] ~^ image[12][20])} + {7'd0,(kernel[3][2] ~^ image[12][21])} + {7'd0,(kernel[3][3] ~^ image[12][22])} + {7'd0,(kernel[3][4] ~^ image[12][23])} + {7'd0,(kernel[4][0] ~^ image[13][19])} + {7'd0,(kernel[4][1] ~^ image[13][20])} + {7'd0,(kernel[4][2] ~^ image[13][21])} + {7'd0,(kernel[4][3] ~^ image[13][22])} + {7'd0,(kernel[4][4] ~^ image[13][23])};
assign out_fmap[9][20][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[9][20])} + {7'd0,(kernel[0][1] ~^ image[9][21])} + {7'd0,(kernel[0][2] ~^ image[9][22])} + {7'd0,(kernel[0][3] ~^ image[9][23])} + {7'd0,(kernel[0][4] ~^ image[9][24])} + {7'd0,(kernel[1][0] ~^ image[10][20])} + {7'd0,(kernel[1][1] ~^ image[10][21])} + {7'd0,(kernel[1][2] ~^ image[10][22])} + {7'd0,(kernel[1][3] ~^ image[10][23])} + {7'd0,(kernel[1][4] ~^ image[10][24])} + {7'd0,(kernel[2][0] ~^ image[11][20])} + {7'd0,(kernel[2][1] ~^ image[11][21])} + {7'd0,(kernel[2][2] ~^ image[11][22])} + {7'd0,(kernel[2][3] ~^ image[11][23])} + {7'd0,(kernel[2][4] ~^ image[11][24])} + {7'd0,(kernel[3][0] ~^ image[12][20])} + {7'd0,(kernel[3][1] ~^ image[12][21])} + {7'd0,(kernel[3][2] ~^ image[12][22])} + {7'd0,(kernel[3][3] ~^ image[12][23])} + {7'd0,(kernel[3][4] ~^ image[12][24])} + {7'd0,(kernel[4][0] ~^ image[13][20])} + {7'd0,(kernel[4][1] ~^ image[13][21])} + {7'd0,(kernel[4][2] ~^ image[13][22])} + {7'd0,(kernel[4][3] ~^ image[13][23])} + {7'd0,(kernel[4][4] ~^ image[13][24])};
assign out_fmap[9][21][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[9][21])} + {7'd0,(kernel[0][1] ~^ image[9][22])} + {7'd0,(kernel[0][2] ~^ image[9][23])} + {7'd0,(kernel[0][3] ~^ image[9][24])} + {7'd0,(kernel[0][4] ~^ image[9][25])} + {7'd0,(kernel[1][0] ~^ image[10][21])} + {7'd0,(kernel[1][1] ~^ image[10][22])} + {7'd0,(kernel[1][2] ~^ image[10][23])} + {7'd0,(kernel[1][3] ~^ image[10][24])} + {7'd0,(kernel[1][4] ~^ image[10][25])} + {7'd0,(kernel[2][0] ~^ image[11][21])} + {7'd0,(kernel[2][1] ~^ image[11][22])} + {7'd0,(kernel[2][2] ~^ image[11][23])} + {7'd0,(kernel[2][3] ~^ image[11][24])} + {7'd0,(kernel[2][4] ~^ image[11][25])} + {7'd0,(kernel[3][0] ~^ image[12][21])} + {7'd0,(kernel[3][1] ~^ image[12][22])} + {7'd0,(kernel[3][2] ~^ image[12][23])} + {7'd0,(kernel[3][3] ~^ image[12][24])} + {7'd0,(kernel[3][4] ~^ image[12][25])} + {7'd0,(kernel[4][0] ~^ image[13][21])} + {7'd0,(kernel[4][1] ~^ image[13][22])} + {7'd0,(kernel[4][2] ~^ image[13][23])} + {7'd0,(kernel[4][3] ~^ image[13][24])} + {7'd0,(kernel[4][4] ~^ image[13][25])};
assign out_fmap[9][22][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[9][22])} + {7'd0,(kernel[0][1] ~^ image[9][23])} + {7'd0,(kernel[0][2] ~^ image[9][24])} + {7'd0,(kernel[0][3] ~^ image[9][25])} + {7'd0,(kernel[0][4] ~^ image[9][26])} + {7'd0,(kernel[1][0] ~^ image[10][22])} + {7'd0,(kernel[1][1] ~^ image[10][23])} + {7'd0,(kernel[1][2] ~^ image[10][24])} + {7'd0,(kernel[1][3] ~^ image[10][25])} + {7'd0,(kernel[1][4] ~^ image[10][26])} + {7'd0,(kernel[2][0] ~^ image[11][22])} + {7'd0,(kernel[2][1] ~^ image[11][23])} + {7'd0,(kernel[2][2] ~^ image[11][24])} + {7'd0,(kernel[2][3] ~^ image[11][25])} + {7'd0,(kernel[2][4] ~^ image[11][26])} + {7'd0,(kernel[3][0] ~^ image[12][22])} + {7'd0,(kernel[3][1] ~^ image[12][23])} + {7'd0,(kernel[3][2] ~^ image[12][24])} + {7'd0,(kernel[3][3] ~^ image[12][25])} + {7'd0,(kernel[3][4] ~^ image[12][26])} + {7'd0,(kernel[4][0] ~^ image[13][22])} + {7'd0,(kernel[4][1] ~^ image[13][23])} + {7'd0,(kernel[4][2] ~^ image[13][24])} + {7'd0,(kernel[4][3] ~^ image[13][25])} + {7'd0,(kernel[4][4] ~^ image[13][26])};
assign out_fmap[9][23][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[9][23])} + {7'd0,(kernel[0][1] ~^ image[9][24])} + {7'd0,(kernel[0][2] ~^ image[9][25])} + {7'd0,(kernel[0][3] ~^ image[9][26])} + {7'd0,(kernel[0][4] ~^ image[9][27])} + {7'd0,(kernel[1][0] ~^ image[10][23])} + {7'd0,(kernel[1][1] ~^ image[10][24])} + {7'd0,(kernel[1][2] ~^ image[10][25])} + {7'd0,(kernel[1][3] ~^ image[10][26])} + {7'd0,(kernel[1][4] ~^ image[10][27])} + {7'd0,(kernel[2][0] ~^ image[11][23])} + {7'd0,(kernel[2][1] ~^ image[11][24])} + {7'd0,(kernel[2][2] ~^ image[11][25])} + {7'd0,(kernel[2][3] ~^ image[11][26])} + {7'd0,(kernel[2][4] ~^ image[11][27])} + {7'd0,(kernel[3][0] ~^ image[12][23])} + {7'd0,(kernel[3][1] ~^ image[12][24])} + {7'd0,(kernel[3][2] ~^ image[12][25])} + {7'd0,(kernel[3][3] ~^ image[12][26])} + {7'd0,(kernel[3][4] ~^ image[12][27])} + {7'd0,(kernel[4][0] ~^ image[13][23])} + {7'd0,(kernel[4][1] ~^ image[13][24])} + {7'd0,(kernel[4][2] ~^ image[13][25])} + {7'd0,(kernel[4][3] ~^ image[13][26])} + {7'd0,(kernel[4][4] ~^ image[13][27])};
assign out_fmap[10][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[10][0])} + {7'd0,(kernel[0][1] ~^ image[10][1])} + {7'd0,(kernel[0][2] ~^ image[10][2])} + {7'd0,(kernel[0][3] ~^ image[10][3])} + {7'd0,(kernel[0][4] ~^ image[10][4])} + {7'd0,(kernel[1][0] ~^ image[11][0])} + {7'd0,(kernel[1][1] ~^ image[11][1])} + {7'd0,(kernel[1][2] ~^ image[11][2])} + {7'd0,(kernel[1][3] ~^ image[11][3])} + {7'd0,(kernel[1][4] ~^ image[11][4])} + {7'd0,(kernel[2][0] ~^ image[12][0])} + {7'd0,(kernel[2][1] ~^ image[12][1])} + {7'd0,(kernel[2][2] ~^ image[12][2])} + {7'd0,(kernel[2][3] ~^ image[12][3])} + {7'd0,(kernel[2][4] ~^ image[12][4])} + {7'd0,(kernel[3][0] ~^ image[13][0])} + {7'd0,(kernel[3][1] ~^ image[13][1])} + {7'd0,(kernel[3][2] ~^ image[13][2])} + {7'd0,(kernel[3][3] ~^ image[13][3])} + {7'd0,(kernel[3][4] ~^ image[13][4])} + {7'd0,(kernel[4][0] ~^ image[14][0])} + {7'd0,(kernel[4][1] ~^ image[14][1])} + {7'd0,(kernel[4][2] ~^ image[14][2])} + {7'd0,(kernel[4][3] ~^ image[14][3])} + {7'd0,(kernel[4][4] ~^ image[14][4])};
assign out_fmap[10][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[10][1])} + {7'd0,(kernel[0][1] ~^ image[10][2])} + {7'd0,(kernel[0][2] ~^ image[10][3])} + {7'd0,(kernel[0][3] ~^ image[10][4])} + {7'd0,(kernel[0][4] ~^ image[10][5])} + {7'd0,(kernel[1][0] ~^ image[11][1])} + {7'd0,(kernel[1][1] ~^ image[11][2])} + {7'd0,(kernel[1][2] ~^ image[11][3])} + {7'd0,(kernel[1][3] ~^ image[11][4])} + {7'd0,(kernel[1][4] ~^ image[11][5])} + {7'd0,(kernel[2][0] ~^ image[12][1])} + {7'd0,(kernel[2][1] ~^ image[12][2])} + {7'd0,(kernel[2][2] ~^ image[12][3])} + {7'd0,(kernel[2][3] ~^ image[12][4])} + {7'd0,(kernel[2][4] ~^ image[12][5])} + {7'd0,(kernel[3][0] ~^ image[13][1])} + {7'd0,(kernel[3][1] ~^ image[13][2])} + {7'd0,(kernel[3][2] ~^ image[13][3])} + {7'd0,(kernel[3][3] ~^ image[13][4])} + {7'd0,(kernel[3][4] ~^ image[13][5])} + {7'd0,(kernel[4][0] ~^ image[14][1])} + {7'd0,(kernel[4][1] ~^ image[14][2])} + {7'd0,(kernel[4][2] ~^ image[14][3])} + {7'd0,(kernel[4][3] ~^ image[14][4])} + {7'd0,(kernel[4][4] ~^ image[14][5])};
assign out_fmap[10][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[10][2])} + {7'd0,(kernel[0][1] ~^ image[10][3])} + {7'd0,(kernel[0][2] ~^ image[10][4])} + {7'd0,(kernel[0][3] ~^ image[10][5])} + {7'd0,(kernel[0][4] ~^ image[10][6])} + {7'd0,(kernel[1][0] ~^ image[11][2])} + {7'd0,(kernel[1][1] ~^ image[11][3])} + {7'd0,(kernel[1][2] ~^ image[11][4])} + {7'd0,(kernel[1][3] ~^ image[11][5])} + {7'd0,(kernel[1][4] ~^ image[11][6])} + {7'd0,(kernel[2][0] ~^ image[12][2])} + {7'd0,(kernel[2][1] ~^ image[12][3])} + {7'd0,(kernel[2][2] ~^ image[12][4])} + {7'd0,(kernel[2][3] ~^ image[12][5])} + {7'd0,(kernel[2][4] ~^ image[12][6])} + {7'd0,(kernel[3][0] ~^ image[13][2])} + {7'd0,(kernel[3][1] ~^ image[13][3])} + {7'd0,(kernel[3][2] ~^ image[13][4])} + {7'd0,(kernel[3][3] ~^ image[13][5])} + {7'd0,(kernel[3][4] ~^ image[13][6])} + {7'd0,(kernel[4][0] ~^ image[14][2])} + {7'd0,(kernel[4][1] ~^ image[14][3])} + {7'd0,(kernel[4][2] ~^ image[14][4])} + {7'd0,(kernel[4][3] ~^ image[14][5])} + {7'd0,(kernel[4][4] ~^ image[14][6])};
assign out_fmap[10][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[10][3])} + {7'd0,(kernel[0][1] ~^ image[10][4])} + {7'd0,(kernel[0][2] ~^ image[10][5])} + {7'd0,(kernel[0][3] ~^ image[10][6])} + {7'd0,(kernel[0][4] ~^ image[10][7])} + {7'd0,(kernel[1][0] ~^ image[11][3])} + {7'd0,(kernel[1][1] ~^ image[11][4])} + {7'd0,(kernel[1][2] ~^ image[11][5])} + {7'd0,(kernel[1][3] ~^ image[11][6])} + {7'd0,(kernel[1][4] ~^ image[11][7])} + {7'd0,(kernel[2][0] ~^ image[12][3])} + {7'd0,(kernel[2][1] ~^ image[12][4])} + {7'd0,(kernel[2][2] ~^ image[12][5])} + {7'd0,(kernel[2][3] ~^ image[12][6])} + {7'd0,(kernel[2][4] ~^ image[12][7])} + {7'd0,(kernel[3][0] ~^ image[13][3])} + {7'd0,(kernel[3][1] ~^ image[13][4])} + {7'd0,(kernel[3][2] ~^ image[13][5])} + {7'd0,(kernel[3][3] ~^ image[13][6])} + {7'd0,(kernel[3][4] ~^ image[13][7])} + {7'd0,(kernel[4][0] ~^ image[14][3])} + {7'd0,(kernel[4][1] ~^ image[14][4])} + {7'd0,(kernel[4][2] ~^ image[14][5])} + {7'd0,(kernel[4][3] ~^ image[14][6])} + {7'd0,(kernel[4][4] ~^ image[14][7])};
assign out_fmap[10][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[10][4])} + {7'd0,(kernel[0][1] ~^ image[10][5])} + {7'd0,(kernel[0][2] ~^ image[10][6])} + {7'd0,(kernel[0][3] ~^ image[10][7])} + {7'd0,(kernel[0][4] ~^ image[10][8])} + {7'd0,(kernel[1][0] ~^ image[11][4])} + {7'd0,(kernel[1][1] ~^ image[11][5])} + {7'd0,(kernel[1][2] ~^ image[11][6])} + {7'd0,(kernel[1][3] ~^ image[11][7])} + {7'd0,(kernel[1][4] ~^ image[11][8])} + {7'd0,(kernel[2][0] ~^ image[12][4])} + {7'd0,(kernel[2][1] ~^ image[12][5])} + {7'd0,(kernel[2][2] ~^ image[12][6])} + {7'd0,(kernel[2][3] ~^ image[12][7])} + {7'd0,(kernel[2][4] ~^ image[12][8])} + {7'd0,(kernel[3][0] ~^ image[13][4])} + {7'd0,(kernel[3][1] ~^ image[13][5])} + {7'd0,(kernel[3][2] ~^ image[13][6])} + {7'd0,(kernel[3][3] ~^ image[13][7])} + {7'd0,(kernel[3][4] ~^ image[13][8])} + {7'd0,(kernel[4][0] ~^ image[14][4])} + {7'd0,(kernel[4][1] ~^ image[14][5])} + {7'd0,(kernel[4][2] ~^ image[14][6])} + {7'd0,(kernel[4][3] ~^ image[14][7])} + {7'd0,(kernel[4][4] ~^ image[14][8])};
assign out_fmap[10][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[10][5])} + {7'd0,(kernel[0][1] ~^ image[10][6])} + {7'd0,(kernel[0][2] ~^ image[10][7])} + {7'd0,(kernel[0][3] ~^ image[10][8])} + {7'd0,(kernel[0][4] ~^ image[10][9])} + {7'd0,(kernel[1][0] ~^ image[11][5])} + {7'd0,(kernel[1][1] ~^ image[11][6])} + {7'd0,(kernel[1][2] ~^ image[11][7])} + {7'd0,(kernel[1][3] ~^ image[11][8])} + {7'd0,(kernel[1][4] ~^ image[11][9])} + {7'd0,(kernel[2][0] ~^ image[12][5])} + {7'd0,(kernel[2][1] ~^ image[12][6])} + {7'd0,(kernel[2][2] ~^ image[12][7])} + {7'd0,(kernel[2][3] ~^ image[12][8])} + {7'd0,(kernel[2][4] ~^ image[12][9])} + {7'd0,(kernel[3][0] ~^ image[13][5])} + {7'd0,(kernel[3][1] ~^ image[13][6])} + {7'd0,(kernel[3][2] ~^ image[13][7])} + {7'd0,(kernel[3][3] ~^ image[13][8])} + {7'd0,(kernel[3][4] ~^ image[13][9])} + {7'd0,(kernel[4][0] ~^ image[14][5])} + {7'd0,(kernel[4][1] ~^ image[14][6])} + {7'd0,(kernel[4][2] ~^ image[14][7])} + {7'd0,(kernel[4][3] ~^ image[14][8])} + {7'd0,(kernel[4][4] ~^ image[14][9])};
assign out_fmap[10][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[10][6])} + {7'd0,(kernel[0][1] ~^ image[10][7])} + {7'd0,(kernel[0][2] ~^ image[10][8])} + {7'd0,(kernel[0][3] ~^ image[10][9])} + {7'd0,(kernel[0][4] ~^ image[10][10])} + {7'd0,(kernel[1][0] ~^ image[11][6])} + {7'd0,(kernel[1][1] ~^ image[11][7])} + {7'd0,(kernel[1][2] ~^ image[11][8])} + {7'd0,(kernel[1][3] ~^ image[11][9])} + {7'd0,(kernel[1][4] ~^ image[11][10])} + {7'd0,(kernel[2][0] ~^ image[12][6])} + {7'd0,(kernel[2][1] ~^ image[12][7])} + {7'd0,(kernel[2][2] ~^ image[12][8])} + {7'd0,(kernel[2][3] ~^ image[12][9])} + {7'd0,(kernel[2][4] ~^ image[12][10])} + {7'd0,(kernel[3][0] ~^ image[13][6])} + {7'd0,(kernel[3][1] ~^ image[13][7])} + {7'd0,(kernel[3][2] ~^ image[13][8])} + {7'd0,(kernel[3][3] ~^ image[13][9])} + {7'd0,(kernel[3][4] ~^ image[13][10])} + {7'd0,(kernel[4][0] ~^ image[14][6])} + {7'd0,(kernel[4][1] ~^ image[14][7])} + {7'd0,(kernel[4][2] ~^ image[14][8])} + {7'd0,(kernel[4][3] ~^ image[14][9])} + {7'd0,(kernel[4][4] ~^ image[14][10])};
assign out_fmap[10][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[10][7])} + {7'd0,(kernel[0][1] ~^ image[10][8])} + {7'd0,(kernel[0][2] ~^ image[10][9])} + {7'd0,(kernel[0][3] ~^ image[10][10])} + {7'd0,(kernel[0][4] ~^ image[10][11])} + {7'd0,(kernel[1][0] ~^ image[11][7])} + {7'd0,(kernel[1][1] ~^ image[11][8])} + {7'd0,(kernel[1][2] ~^ image[11][9])} + {7'd0,(kernel[1][3] ~^ image[11][10])} + {7'd0,(kernel[1][4] ~^ image[11][11])} + {7'd0,(kernel[2][0] ~^ image[12][7])} + {7'd0,(kernel[2][1] ~^ image[12][8])} + {7'd0,(kernel[2][2] ~^ image[12][9])} + {7'd0,(kernel[2][3] ~^ image[12][10])} + {7'd0,(kernel[2][4] ~^ image[12][11])} + {7'd0,(kernel[3][0] ~^ image[13][7])} + {7'd0,(kernel[3][1] ~^ image[13][8])} + {7'd0,(kernel[3][2] ~^ image[13][9])} + {7'd0,(kernel[3][3] ~^ image[13][10])} + {7'd0,(kernel[3][4] ~^ image[13][11])} + {7'd0,(kernel[4][0] ~^ image[14][7])} + {7'd0,(kernel[4][1] ~^ image[14][8])} + {7'd0,(kernel[4][2] ~^ image[14][9])} + {7'd0,(kernel[4][3] ~^ image[14][10])} + {7'd0,(kernel[4][4] ~^ image[14][11])};
assign out_fmap[10][8][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[10][8])} + {7'd0,(kernel[0][1] ~^ image[10][9])} + {7'd0,(kernel[0][2] ~^ image[10][10])} + {7'd0,(kernel[0][3] ~^ image[10][11])} + {7'd0,(kernel[0][4] ~^ image[10][12])} + {7'd0,(kernel[1][0] ~^ image[11][8])} + {7'd0,(kernel[1][1] ~^ image[11][9])} + {7'd0,(kernel[1][2] ~^ image[11][10])} + {7'd0,(kernel[1][3] ~^ image[11][11])} + {7'd0,(kernel[1][4] ~^ image[11][12])} + {7'd0,(kernel[2][0] ~^ image[12][8])} + {7'd0,(kernel[2][1] ~^ image[12][9])} + {7'd0,(kernel[2][2] ~^ image[12][10])} + {7'd0,(kernel[2][3] ~^ image[12][11])} + {7'd0,(kernel[2][4] ~^ image[12][12])} + {7'd0,(kernel[3][0] ~^ image[13][8])} + {7'd0,(kernel[3][1] ~^ image[13][9])} + {7'd0,(kernel[3][2] ~^ image[13][10])} + {7'd0,(kernel[3][3] ~^ image[13][11])} + {7'd0,(kernel[3][4] ~^ image[13][12])} + {7'd0,(kernel[4][0] ~^ image[14][8])} + {7'd0,(kernel[4][1] ~^ image[14][9])} + {7'd0,(kernel[4][2] ~^ image[14][10])} + {7'd0,(kernel[4][3] ~^ image[14][11])} + {7'd0,(kernel[4][4] ~^ image[14][12])};
assign out_fmap[10][9][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[10][9])} + {7'd0,(kernel[0][1] ~^ image[10][10])} + {7'd0,(kernel[0][2] ~^ image[10][11])} + {7'd0,(kernel[0][3] ~^ image[10][12])} + {7'd0,(kernel[0][4] ~^ image[10][13])} + {7'd0,(kernel[1][0] ~^ image[11][9])} + {7'd0,(kernel[1][1] ~^ image[11][10])} + {7'd0,(kernel[1][2] ~^ image[11][11])} + {7'd0,(kernel[1][3] ~^ image[11][12])} + {7'd0,(kernel[1][4] ~^ image[11][13])} + {7'd0,(kernel[2][0] ~^ image[12][9])} + {7'd0,(kernel[2][1] ~^ image[12][10])} + {7'd0,(kernel[2][2] ~^ image[12][11])} + {7'd0,(kernel[2][3] ~^ image[12][12])} + {7'd0,(kernel[2][4] ~^ image[12][13])} + {7'd0,(kernel[3][0] ~^ image[13][9])} + {7'd0,(kernel[3][1] ~^ image[13][10])} + {7'd0,(kernel[3][2] ~^ image[13][11])} + {7'd0,(kernel[3][3] ~^ image[13][12])} + {7'd0,(kernel[3][4] ~^ image[13][13])} + {7'd0,(kernel[4][0] ~^ image[14][9])} + {7'd0,(kernel[4][1] ~^ image[14][10])} + {7'd0,(kernel[4][2] ~^ image[14][11])} + {7'd0,(kernel[4][3] ~^ image[14][12])} + {7'd0,(kernel[4][4] ~^ image[14][13])};
assign out_fmap[10][10][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[10][10])} + {7'd0,(kernel[0][1] ~^ image[10][11])} + {7'd0,(kernel[0][2] ~^ image[10][12])} + {7'd0,(kernel[0][3] ~^ image[10][13])} + {7'd0,(kernel[0][4] ~^ image[10][14])} + {7'd0,(kernel[1][0] ~^ image[11][10])} + {7'd0,(kernel[1][1] ~^ image[11][11])} + {7'd0,(kernel[1][2] ~^ image[11][12])} + {7'd0,(kernel[1][3] ~^ image[11][13])} + {7'd0,(kernel[1][4] ~^ image[11][14])} + {7'd0,(kernel[2][0] ~^ image[12][10])} + {7'd0,(kernel[2][1] ~^ image[12][11])} + {7'd0,(kernel[2][2] ~^ image[12][12])} + {7'd0,(kernel[2][3] ~^ image[12][13])} + {7'd0,(kernel[2][4] ~^ image[12][14])} + {7'd0,(kernel[3][0] ~^ image[13][10])} + {7'd0,(kernel[3][1] ~^ image[13][11])} + {7'd0,(kernel[3][2] ~^ image[13][12])} + {7'd0,(kernel[3][3] ~^ image[13][13])} + {7'd0,(kernel[3][4] ~^ image[13][14])} + {7'd0,(kernel[4][0] ~^ image[14][10])} + {7'd0,(kernel[4][1] ~^ image[14][11])} + {7'd0,(kernel[4][2] ~^ image[14][12])} + {7'd0,(kernel[4][3] ~^ image[14][13])} + {7'd0,(kernel[4][4] ~^ image[14][14])};
assign out_fmap[10][11][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[10][11])} + {7'd0,(kernel[0][1] ~^ image[10][12])} + {7'd0,(kernel[0][2] ~^ image[10][13])} + {7'd0,(kernel[0][3] ~^ image[10][14])} + {7'd0,(kernel[0][4] ~^ image[10][15])} + {7'd0,(kernel[1][0] ~^ image[11][11])} + {7'd0,(kernel[1][1] ~^ image[11][12])} + {7'd0,(kernel[1][2] ~^ image[11][13])} + {7'd0,(kernel[1][3] ~^ image[11][14])} + {7'd0,(kernel[1][4] ~^ image[11][15])} + {7'd0,(kernel[2][0] ~^ image[12][11])} + {7'd0,(kernel[2][1] ~^ image[12][12])} + {7'd0,(kernel[2][2] ~^ image[12][13])} + {7'd0,(kernel[2][3] ~^ image[12][14])} + {7'd0,(kernel[2][4] ~^ image[12][15])} + {7'd0,(kernel[3][0] ~^ image[13][11])} + {7'd0,(kernel[3][1] ~^ image[13][12])} + {7'd0,(kernel[3][2] ~^ image[13][13])} + {7'd0,(kernel[3][3] ~^ image[13][14])} + {7'd0,(kernel[3][4] ~^ image[13][15])} + {7'd0,(kernel[4][0] ~^ image[14][11])} + {7'd0,(kernel[4][1] ~^ image[14][12])} + {7'd0,(kernel[4][2] ~^ image[14][13])} + {7'd0,(kernel[4][3] ~^ image[14][14])} + {7'd0,(kernel[4][4] ~^ image[14][15])};
assign out_fmap[10][12][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[10][12])} + {7'd0,(kernel[0][1] ~^ image[10][13])} + {7'd0,(kernel[0][2] ~^ image[10][14])} + {7'd0,(kernel[0][3] ~^ image[10][15])} + {7'd0,(kernel[0][4] ~^ image[10][16])} + {7'd0,(kernel[1][0] ~^ image[11][12])} + {7'd0,(kernel[1][1] ~^ image[11][13])} + {7'd0,(kernel[1][2] ~^ image[11][14])} + {7'd0,(kernel[1][3] ~^ image[11][15])} + {7'd0,(kernel[1][4] ~^ image[11][16])} + {7'd0,(kernel[2][0] ~^ image[12][12])} + {7'd0,(kernel[2][1] ~^ image[12][13])} + {7'd0,(kernel[2][2] ~^ image[12][14])} + {7'd0,(kernel[2][3] ~^ image[12][15])} + {7'd0,(kernel[2][4] ~^ image[12][16])} + {7'd0,(kernel[3][0] ~^ image[13][12])} + {7'd0,(kernel[3][1] ~^ image[13][13])} + {7'd0,(kernel[3][2] ~^ image[13][14])} + {7'd0,(kernel[3][3] ~^ image[13][15])} + {7'd0,(kernel[3][4] ~^ image[13][16])} + {7'd0,(kernel[4][0] ~^ image[14][12])} + {7'd0,(kernel[4][1] ~^ image[14][13])} + {7'd0,(kernel[4][2] ~^ image[14][14])} + {7'd0,(kernel[4][3] ~^ image[14][15])} + {7'd0,(kernel[4][4] ~^ image[14][16])};
assign out_fmap[10][13][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[10][13])} + {7'd0,(kernel[0][1] ~^ image[10][14])} + {7'd0,(kernel[0][2] ~^ image[10][15])} + {7'd0,(kernel[0][3] ~^ image[10][16])} + {7'd0,(kernel[0][4] ~^ image[10][17])} + {7'd0,(kernel[1][0] ~^ image[11][13])} + {7'd0,(kernel[1][1] ~^ image[11][14])} + {7'd0,(kernel[1][2] ~^ image[11][15])} + {7'd0,(kernel[1][3] ~^ image[11][16])} + {7'd0,(kernel[1][4] ~^ image[11][17])} + {7'd0,(kernel[2][0] ~^ image[12][13])} + {7'd0,(kernel[2][1] ~^ image[12][14])} + {7'd0,(kernel[2][2] ~^ image[12][15])} + {7'd0,(kernel[2][3] ~^ image[12][16])} + {7'd0,(kernel[2][4] ~^ image[12][17])} + {7'd0,(kernel[3][0] ~^ image[13][13])} + {7'd0,(kernel[3][1] ~^ image[13][14])} + {7'd0,(kernel[3][2] ~^ image[13][15])} + {7'd0,(kernel[3][3] ~^ image[13][16])} + {7'd0,(kernel[3][4] ~^ image[13][17])} + {7'd0,(kernel[4][0] ~^ image[14][13])} + {7'd0,(kernel[4][1] ~^ image[14][14])} + {7'd0,(kernel[4][2] ~^ image[14][15])} + {7'd0,(kernel[4][3] ~^ image[14][16])} + {7'd0,(kernel[4][4] ~^ image[14][17])};
assign out_fmap[10][14][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[10][14])} + {7'd0,(kernel[0][1] ~^ image[10][15])} + {7'd0,(kernel[0][2] ~^ image[10][16])} + {7'd0,(kernel[0][3] ~^ image[10][17])} + {7'd0,(kernel[0][4] ~^ image[10][18])} + {7'd0,(kernel[1][0] ~^ image[11][14])} + {7'd0,(kernel[1][1] ~^ image[11][15])} + {7'd0,(kernel[1][2] ~^ image[11][16])} + {7'd0,(kernel[1][3] ~^ image[11][17])} + {7'd0,(kernel[1][4] ~^ image[11][18])} + {7'd0,(kernel[2][0] ~^ image[12][14])} + {7'd0,(kernel[2][1] ~^ image[12][15])} + {7'd0,(kernel[2][2] ~^ image[12][16])} + {7'd0,(kernel[2][3] ~^ image[12][17])} + {7'd0,(kernel[2][4] ~^ image[12][18])} + {7'd0,(kernel[3][0] ~^ image[13][14])} + {7'd0,(kernel[3][1] ~^ image[13][15])} + {7'd0,(kernel[3][2] ~^ image[13][16])} + {7'd0,(kernel[3][3] ~^ image[13][17])} + {7'd0,(kernel[3][4] ~^ image[13][18])} + {7'd0,(kernel[4][0] ~^ image[14][14])} + {7'd0,(kernel[4][1] ~^ image[14][15])} + {7'd0,(kernel[4][2] ~^ image[14][16])} + {7'd0,(kernel[4][3] ~^ image[14][17])} + {7'd0,(kernel[4][4] ~^ image[14][18])};
assign out_fmap[10][15][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[10][15])} + {7'd0,(kernel[0][1] ~^ image[10][16])} + {7'd0,(kernel[0][2] ~^ image[10][17])} + {7'd0,(kernel[0][3] ~^ image[10][18])} + {7'd0,(kernel[0][4] ~^ image[10][19])} + {7'd0,(kernel[1][0] ~^ image[11][15])} + {7'd0,(kernel[1][1] ~^ image[11][16])} + {7'd0,(kernel[1][2] ~^ image[11][17])} + {7'd0,(kernel[1][3] ~^ image[11][18])} + {7'd0,(kernel[1][4] ~^ image[11][19])} + {7'd0,(kernel[2][0] ~^ image[12][15])} + {7'd0,(kernel[2][1] ~^ image[12][16])} + {7'd0,(kernel[2][2] ~^ image[12][17])} + {7'd0,(kernel[2][3] ~^ image[12][18])} + {7'd0,(kernel[2][4] ~^ image[12][19])} + {7'd0,(kernel[3][0] ~^ image[13][15])} + {7'd0,(kernel[3][1] ~^ image[13][16])} + {7'd0,(kernel[3][2] ~^ image[13][17])} + {7'd0,(kernel[3][3] ~^ image[13][18])} + {7'd0,(kernel[3][4] ~^ image[13][19])} + {7'd0,(kernel[4][0] ~^ image[14][15])} + {7'd0,(kernel[4][1] ~^ image[14][16])} + {7'd0,(kernel[4][2] ~^ image[14][17])} + {7'd0,(kernel[4][3] ~^ image[14][18])} + {7'd0,(kernel[4][4] ~^ image[14][19])};
assign out_fmap[10][16][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[10][16])} + {7'd0,(kernel[0][1] ~^ image[10][17])} + {7'd0,(kernel[0][2] ~^ image[10][18])} + {7'd0,(kernel[0][3] ~^ image[10][19])} + {7'd0,(kernel[0][4] ~^ image[10][20])} + {7'd0,(kernel[1][0] ~^ image[11][16])} + {7'd0,(kernel[1][1] ~^ image[11][17])} + {7'd0,(kernel[1][2] ~^ image[11][18])} + {7'd0,(kernel[1][3] ~^ image[11][19])} + {7'd0,(kernel[1][4] ~^ image[11][20])} + {7'd0,(kernel[2][0] ~^ image[12][16])} + {7'd0,(kernel[2][1] ~^ image[12][17])} + {7'd0,(kernel[2][2] ~^ image[12][18])} + {7'd0,(kernel[2][3] ~^ image[12][19])} + {7'd0,(kernel[2][4] ~^ image[12][20])} + {7'd0,(kernel[3][0] ~^ image[13][16])} + {7'd0,(kernel[3][1] ~^ image[13][17])} + {7'd0,(kernel[3][2] ~^ image[13][18])} + {7'd0,(kernel[3][3] ~^ image[13][19])} + {7'd0,(kernel[3][4] ~^ image[13][20])} + {7'd0,(kernel[4][0] ~^ image[14][16])} + {7'd0,(kernel[4][1] ~^ image[14][17])} + {7'd0,(kernel[4][2] ~^ image[14][18])} + {7'd0,(kernel[4][3] ~^ image[14][19])} + {7'd0,(kernel[4][4] ~^ image[14][20])};
assign out_fmap[10][17][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[10][17])} + {7'd0,(kernel[0][1] ~^ image[10][18])} + {7'd0,(kernel[0][2] ~^ image[10][19])} + {7'd0,(kernel[0][3] ~^ image[10][20])} + {7'd0,(kernel[0][4] ~^ image[10][21])} + {7'd0,(kernel[1][0] ~^ image[11][17])} + {7'd0,(kernel[1][1] ~^ image[11][18])} + {7'd0,(kernel[1][2] ~^ image[11][19])} + {7'd0,(kernel[1][3] ~^ image[11][20])} + {7'd0,(kernel[1][4] ~^ image[11][21])} + {7'd0,(kernel[2][0] ~^ image[12][17])} + {7'd0,(kernel[2][1] ~^ image[12][18])} + {7'd0,(kernel[2][2] ~^ image[12][19])} + {7'd0,(kernel[2][3] ~^ image[12][20])} + {7'd0,(kernel[2][4] ~^ image[12][21])} + {7'd0,(kernel[3][0] ~^ image[13][17])} + {7'd0,(kernel[3][1] ~^ image[13][18])} + {7'd0,(kernel[3][2] ~^ image[13][19])} + {7'd0,(kernel[3][3] ~^ image[13][20])} + {7'd0,(kernel[3][4] ~^ image[13][21])} + {7'd0,(kernel[4][0] ~^ image[14][17])} + {7'd0,(kernel[4][1] ~^ image[14][18])} + {7'd0,(kernel[4][2] ~^ image[14][19])} + {7'd0,(kernel[4][3] ~^ image[14][20])} + {7'd0,(kernel[4][4] ~^ image[14][21])};
assign out_fmap[10][18][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[10][18])} + {7'd0,(kernel[0][1] ~^ image[10][19])} + {7'd0,(kernel[0][2] ~^ image[10][20])} + {7'd0,(kernel[0][3] ~^ image[10][21])} + {7'd0,(kernel[0][4] ~^ image[10][22])} + {7'd0,(kernel[1][0] ~^ image[11][18])} + {7'd0,(kernel[1][1] ~^ image[11][19])} + {7'd0,(kernel[1][2] ~^ image[11][20])} + {7'd0,(kernel[1][3] ~^ image[11][21])} + {7'd0,(kernel[1][4] ~^ image[11][22])} + {7'd0,(kernel[2][0] ~^ image[12][18])} + {7'd0,(kernel[2][1] ~^ image[12][19])} + {7'd0,(kernel[2][2] ~^ image[12][20])} + {7'd0,(kernel[2][3] ~^ image[12][21])} + {7'd0,(kernel[2][4] ~^ image[12][22])} + {7'd0,(kernel[3][0] ~^ image[13][18])} + {7'd0,(kernel[3][1] ~^ image[13][19])} + {7'd0,(kernel[3][2] ~^ image[13][20])} + {7'd0,(kernel[3][3] ~^ image[13][21])} + {7'd0,(kernel[3][4] ~^ image[13][22])} + {7'd0,(kernel[4][0] ~^ image[14][18])} + {7'd0,(kernel[4][1] ~^ image[14][19])} + {7'd0,(kernel[4][2] ~^ image[14][20])} + {7'd0,(kernel[4][3] ~^ image[14][21])} + {7'd0,(kernel[4][4] ~^ image[14][22])};
assign out_fmap[10][19][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[10][19])} + {7'd0,(kernel[0][1] ~^ image[10][20])} + {7'd0,(kernel[0][2] ~^ image[10][21])} + {7'd0,(kernel[0][3] ~^ image[10][22])} + {7'd0,(kernel[0][4] ~^ image[10][23])} + {7'd0,(kernel[1][0] ~^ image[11][19])} + {7'd0,(kernel[1][1] ~^ image[11][20])} + {7'd0,(kernel[1][2] ~^ image[11][21])} + {7'd0,(kernel[1][3] ~^ image[11][22])} + {7'd0,(kernel[1][4] ~^ image[11][23])} + {7'd0,(kernel[2][0] ~^ image[12][19])} + {7'd0,(kernel[2][1] ~^ image[12][20])} + {7'd0,(kernel[2][2] ~^ image[12][21])} + {7'd0,(kernel[2][3] ~^ image[12][22])} + {7'd0,(kernel[2][4] ~^ image[12][23])} + {7'd0,(kernel[3][0] ~^ image[13][19])} + {7'd0,(kernel[3][1] ~^ image[13][20])} + {7'd0,(kernel[3][2] ~^ image[13][21])} + {7'd0,(kernel[3][3] ~^ image[13][22])} + {7'd0,(kernel[3][4] ~^ image[13][23])} + {7'd0,(kernel[4][0] ~^ image[14][19])} + {7'd0,(kernel[4][1] ~^ image[14][20])} + {7'd0,(kernel[4][2] ~^ image[14][21])} + {7'd0,(kernel[4][3] ~^ image[14][22])} + {7'd0,(kernel[4][4] ~^ image[14][23])};
assign out_fmap[10][20][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[10][20])} + {7'd0,(kernel[0][1] ~^ image[10][21])} + {7'd0,(kernel[0][2] ~^ image[10][22])} + {7'd0,(kernel[0][3] ~^ image[10][23])} + {7'd0,(kernel[0][4] ~^ image[10][24])} + {7'd0,(kernel[1][0] ~^ image[11][20])} + {7'd0,(kernel[1][1] ~^ image[11][21])} + {7'd0,(kernel[1][2] ~^ image[11][22])} + {7'd0,(kernel[1][3] ~^ image[11][23])} + {7'd0,(kernel[1][4] ~^ image[11][24])} + {7'd0,(kernel[2][0] ~^ image[12][20])} + {7'd0,(kernel[2][1] ~^ image[12][21])} + {7'd0,(kernel[2][2] ~^ image[12][22])} + {7'd0,(kernel[2][3] ~^ image[12][23])} + {7'd0,(kernel[2][4] ~^ image[12][24])} + {7'd0,(kernel[3][0] ~^ image[13][20])} + {7'd0,(kernel[3][1] ~^ image[13][21])} + {7'd0,(kernel[3][2] ~^ image[13][22])} + {7'd0,(kernel[3][3] ~^ image[13][23])} + {7'd0,(kernel[3][4] ~^ image[13][24])} + {7'd0,(kernel[4][0] ~^ image[14][20])} + {7'd0,(kernel[4][1] ~^ image[14][21])} + {7'd0,(kernel[4][2] ~^ image[14][22])} + {7'd0,(kernel[4][3] ~^ image[14][23])} + {7'd0,(kernel[4][4] ~^ image[14][24])};
assign out_fmap[10][21][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[10][21])} + {7'd0,(kernel[0][1] ~^ image[10][22])} + {7'd0,(kernel[0][2] ~^ image[10][23])} + {7'd0,(kernel[0][3] ~^ image[10][24])} + {7'd0,(kernel[0][4] ~^ image[10][25])} + {7'd0,(kernel[1][0] ~^ image[11][21])} + {7'd0,(kernel[1][1] ~^ image[11][22])} + {7'd0,(kernel[1][2] ~^ image[11][23])} + {7'd0,(kernel[1][3] ~^ image[11][24])} + {7'd0,(kernel[1][4] ~^ image[11][25])} + {7'd0,(kernel[2][0] ~^ image[12][21])} + {7'd0,(kernel[2][1] ~^ image[12][22])} + {7'd0,(kernel[2][2] ~^ image[12][23])} + {7'd0,(kernel[2][3] ~^ image[12][24])} + {7'd0,(kernel[2][4] ~^ image[12][25])} + {7'd0,(kernel[3][0] ~^ image[13][21])} + {7'd0,(kernel[3][1] ~^ image[13][22])} + {7'd0,(kernel[3][2] ~^ image[13][23])} + {7'd0,(kernel[3][3] ~^ image[13][24])} + {7'd0,(kernel[3][4] ~^ image[13][25])} + {7'd0,(kernel[4][0] ~^ image[14][21])} + {7'd0,(kernel[4][1] ~^ image[14][22])} + {7'd0,(kernel[4][2] ~^ image[14][23])} + {7'd0,(kernel[4][3] ~^ image[14][24])} + {7'd0,(kernel[4][4] ~^ image[14][25])};
assign out_fmap[10][22][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[10][22])} + {7'd0,(kernel[0][1] ~^ image[10][23])} + {7'd0,(kernel[0][2] ~^ image[10][24])} + {7'd0,(kernel[0][3] ~^ image[10][25])} + {7'd0,(kernel[0][4] ~^ image[10][26])} + {7'd0,(kernel[1][0] ~^ image[11][22])} + {7'd0,(kernel[1][1] ~^ image[11][23])} + {7'd0,(kernel[1][2] ~^ image[11][24])} + {7'd0,(kernel[1][3] ~^ image[11][25])} + {7'd0,(kernel[1][4] ~^ image[11][26])} + {7'd0,(kernel[2][0] ~^ image[12][22])} + {7'd0,(kernel[2][1] ~^ image[12][23])} + {7'd0,(kernel[2][2] ~^ image[12][24])} + {7'd0,(kernel[2][3] ~^ image[12][25])} + {7'd0,(kernel[2][4] ~^ image[12][26])} + {7'd0,(kernel[3][0] ~^ image[13][22])} + {7'd0,(kernel[3][1] ~^ image[13][23])} + {7'd0,(kernel[3][2] ~^ image[13][24])} + {7'd0,(kernel[3][3] ~^ image[13][25])} + {7'd0,(kernel[3][4] ~^ image[13][26])} + {7'd0,(kernel[4][0] ~^ image[14][22])} + {7'd0,(kernel[4][1] ~^ image[14][23])} + {7'd0,(kernel[4][2] ~^ image[14][24])} + {7'd0,(kernel[4][3] ~^ image[14][25])} + {7'd0,(kernel[4][4] ~^ image[14][26])};
assign out_fmap[10][23][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[10][23])} + {7'd0,(kernel[0][1] ~^ image[10][24])} + {7'd0,(kernel[0][2] ~^ image[10][25])} + {7'd0,(kernel[0][3] ~^ image[10][26])} + {7'd0,(kernel[0][4] ~^ image[10][27])} + {7'd0,(kernel[1][0] ~^ image[11][23])} + {7'd0,(kernel[1][1] ~^ image[11][24])} + {7'd0,(kernel[1][2] ~^ image[11][25])} + {7'd0,(kernel[1][3] ~^ image[11][26])} + {7'd0,(kernel[1][4] ~^ image[11][27])} + {7'd0,(kernel[2][0] ~^ image[12][23])} + {7'd0,(kernel[2][1] ~^ image[12][24])} + {7'd0,(kernel[2][2] ~^ image[12][25])} + {7'd0,(kernel[2][3] ~^ image[12][26])} + {7'd0,(kernel[2][4] ~^ image[12][27])} + {7'd0,(kernel[3][0] ~^ image[13][23])} + {7'd0,(kernel[3][1] ~^ image[13][24])} + {7'd0,(kernel[3][2] ~^ image[13][25])} + {7'd0,(kernel[3][3] ~^ image[13][26])} + {7'd0,(kernel[3][4] ~^ image[13][27])} + {7'd0,(kernel[4][0] ~^ image[14][23])} + {7'd0,(kernel[4][1] ~^ image[14][24])} + {7'd0,(kernel[4][2] ~^ image[14][25])} + {7'd0,(kernel[4][3] ~^ image[14][26])} + {7'd0,(kernel[4][4] ~^ image[14][27])};
assign out_fmap[11][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[11][0])} + {7'd0,(kernel[0][1] ~^ image[11][1])} + {7'd0,(kernel[0][2] ~^ image[11][2])} + {7'd0,(kernel[0][3] ~^ image[11][3])} + {7'd0,(kernel[0][4] ~^ image[11][4])} + {7'd0,(kernel[1][0] ~^ image[12][0])} + {7'd0,(kernel[1][1] ~^ image[12][1])} + {7'd0,(kernel[1][2] ~^ image[12][2])} + {7'd0,(kernel[1][3] ~^ image[12][3])} + {7'd0,(kernel[1][4] ~^ image[12][4])} + {7'd0,(kernel[2][0] ~^ image[13][0])} + {7'd0,(kernel[2][1] ~^ image[13][1])} + {7'd0,(kernel[2][2] ~^ image[13][2])} + {7'd0,(kernel[2][3] ~^ image[13][3])} + {7'd0,(kernel[2][4] ~^ image[13][4])} + {7'd0,(kernel[3][0] ~^ image[14][0])} + {7'd0,(kernel[3][1] ~^ image[14][1])} + {7'd0,(kernel[3][2] ~^ image[14][2])} + {7'd0,(kernel[3][3] ~^ image[14][3])} + {7'd0,(kernel[3][4] ~^ image[14][4])} + {7'd0,(kernel[4][0] ~^ image[15][0])} + {7'd0,(kernel[4][1] ~^ image[15][1])} + {7'd0,(kernel[4][2] ~^ image[15][2])} + {7'd0,(kernel[4][3] ~^ image[15][3])} + {7'd0,(kernel[4][4] ~^ image[15][4])};
assign out_fmap[11][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[11][1])} + {7'd0,(kernel[0][1] ~^ image[11][2])} + {7'd0,(kernel[0][2] ~^ image[11][3])} + {7'd0,(kernel[0][3] ~^ image[11][4])} + {7'd0,(kernel[0][4] ~^ image[11][5])} + {7'd0,(kernel[1][0] ~^ image[12][1])} + {7'd0,(kernel[1][1] ~^ image[12][2])} + {7'd0,(kernel[1][2] ~^ image[12][3])} + {7'd0,(kernel[1][3] ~^ image[12][4])} + {7'd0,(kernel[1][4] ~^ image[12][5])} + {7'd0,(kernel[2][0] ~^ image[13][1])} + {7'd0,(kernel[2][1] ~^ image[13][2])} + {7'd0,(kernel[2][2] ~^ image[13][3])} + {7'd0,(kernel[2][3] ~^ image[13][4])} + {7'd0,(kernel[2][4] ~^ image[13][5])} + {7'd0,(kernel[3][0] ~^ image[14][1])} + {7'd0,(kernel[3][1] ~^ image[14][2])} + {7'd0,(kernel[3][2] ~^ image[14][3])} + {7'd0,(kernel[3][3] ~^ image[14][4])} + {7'd0,(kernel[3][4] ~^ image[14][5])} + {7'd0,(kernel[4][0] ~^ image[15][1])} + {7'd0,(kernel[4][1] ~^ image[15][2])} + {7'd0,(kernel[4][2] ~^ image[15][3])} + {7'd0,(kernel[4][3] ~^ image[15][4])} + {7'd0,(kernel[4][4] ~^ image[15][5])};
assign out_fmap[11][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[11][2])} + {7'd0,(kernel[0][1] ~^ image[11][3])} + {7'd0,(kernel[0][2] ~^ image[11][4])} + {7'd0,(kernel[0][3] ~^ image[11][5])} + {7'd0,(kernel[0][4] ~^ image[11][6])} + {7'd0,(kernel[1][0] ~^ image[12][2])} + {7'd0,(kernel[1][1] ~^ image[12][3])} + {7'd0,(kernel[1][2] ~^ image[12][4])} + {7'd0,(kernel[1][3] ~^ image[12][5])} + {7'd0,(kernel[1][4] ~^ image[12][6])} + {7'd0,(kernel[2][0] ~^ image[13][2])} + {7'd0,(kernel[2][1] ~^ image[13][3])} + {7'd0,(kernel[2][2] ~^ image[13][4])} + {7'd0,(kernel[2][3] ~^ image[13][5])} + {7'd0,(kernel[2][4] ~^ image[13][6])} + {7'd0,(kernel[3][0] ~^ image[14][2])} + {7'd0,(kernel[3][1] ~^ image[14][3])} + {7'd0,(kernel[3][2] ~^ image[14][4])} + {7'd0,(kernel[3][3] ~^ image[14][5])} + {7'd0,(kernel[3][4] ~^ image[14][6])} + {7'd0,(kernel[4][0] ~^ image[15][2])} + {7'd0,(kernel[4][1] ~^ image[15][3])} + {7'd0,(kernel[4][2] ~^ image[15][4])} + {7'd0,(kernel[4][3] ~^ image[15][5])} + {7'd0,(kernel[4][4] ~^ image[15][6])};
assign out_fmap[11][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[11][3])} + {7'd0,(kernel[0][1] ~^ image[11][4])} + {7'd0,(kernel[0][2] ~^ image[11][5])} + {7'd0,(kernel[0][3] ~^ image[11][6])} + {7'd0,(kernel[0][4] ~^ image[11][7])} + {7'd0,(kernel[1][0] ~^ image[12][3])} + {7'd0,(kernel[1][1] ~^ image[12][4])} + {7'd0,(kernel[1][2] ~^ image[12][5])} + {7'd0,(kernel[1][3] ~^ image[12][6])} + {7'd0,(kernel[1][4] ~^ image[12][7])} + {7'd0,(kernel[2][0] ~^ image[13][3])} + {7'd0,(kernel[2][1] ~^ image[13][4])} + {7'd0,(kernel[2][2] ~^ image[13][5])} + {7'd0,(kernel[2][3] ~^ image[13][6])} + {7'd0,(kernel[2][4] ~^ image[13][7])} + {7'd0,(kernel[3][0] ~^ image[14][3])} + {7'd0,(kernel[3][1] ~^ image[14][4])} + {7'd0,(kernel[3][2] ~^ image[14][5])} + {7'd0,(kernel[3][3] ~^ image[14][6])} + {7'd0,(kernel[3][4] ~^ image[14][7])} + {7'd0,(kernel[4][0] ~^ image[15][3])} + {7'd0,(kernel[4][1] ~^ image[15][4])} + {7'd0,(kernel[4][2] ~^ image[15][5])} + {7'd0,(kernel[4][3] ~^ image[15][6])} + {7'd0,(kernel[4][4] ~^ image[15][7])};
assign out_fmap[11][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[11][4])} + {7'd0,(kernel[0][1] ~^ image[11][5])} + {7'd0,(kernel[0][2] ~^ image[11][6])} + {7'd0,(kernel[0][3] ~^ image[11][7])} + {7'd0,(kernel[0][4] ~^ image[11][8])} + {7'd0,(kernel[1][0] ~^ image[12][4])} + {7'd0,(kernel[1][1] ~^ image[12][5])} + {7'd0,(kernel[1][2] ~^ image[12][6])} + {7'd0,(kernel[1][3] ~^ image[12][7])} + {7'd0,(kernel[1][4] ~^ image[12][8])} + {7'd0,(kernel[2][0] ~^ image[13][4])} + {7'd0,(kernel[2][1] ~^ image[13][5])} + {7'd0,(kernel[2][2] ~^ image[13][6])} + {7'd0,(kernel[2][3] ~^ image[13][7])} + {7'd0,(kernel[2][4] ~^ image[13][8])} + {7'd0,(kernel[3][0] ~^ image[14][4])} + {7'd0,(kernel[3][1] ~^ image[14][5])} + {7'd0,(kernel[3][2] ~^ image[14][6])} + {7'd0,(kernel[3][3] ~^ image[14][7])} + {7'd0,(kernel[3][4] ~^ image[14][8])} + {7'd0,(kernel[4][0] ~^ image[15][4])} + {7'd0,(kernel[4][1] ~^ image[15][5])} + {7'd0,(kernel[4][2] ~^ image[15][6])} + {7'd0,(kernel[4][3] ~^ image[15][7])} + {7'd0,(kernel[4][4] ~^ image[15][8])};
assign out_fmap[11][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[11][5])} + {7'd0,(kernel[0][1] ~^ image[11][6])} + {7'd0,(kernel[0][2] ~^ image[11][7])} + {7'd0,(kernel[0][3] ~^ image[11][8])} + {7'd0,(kernel[0][4] ~^ image[11][9])} + {7'd0,(kernel[1][0] ~^ image[12][5])} + {7'd0,(kernel[1][1] ~^ image[12][6])} + {7'd0,(kernel[1][2] ~^ image[12][7])} + {7'd0,(kernel[1][3] ~^ image[12][8])} + {7'd0,(kernel[1][4] ~^ image[12][9])} + {7'd0,(kernel[2][0] ~^ image[13][5])} + {7'd0,(kernel[2][1] ~^ image[13][6])} + {7'd0,(kernel[2][2] ~^ image[13][7])} + {7'd0,(kernel[2][3] ~^ image[13][8])} + {7'd0,(kernel[2][4] ~^ image[13][9])} + {7'd0,(kernel[3][0] ~^ image[14][5])} + {7'd0,(kernel[3][1] ~^ image[14][6])} + {7'd0,(kernel[3][2] ~^ image[14][7])} + {7'd0,(kernel[3][3] ~^ image[14][8])} + {7'd0,(kernel[3][4] ~^ image[14][9])} + {7'd0,(kernel[4][0] ~^ image[15][5])} + {7'd0,(kernel[4][1] ~^ image[15][6])} + {7'd0,(kernel[4][2] ~^ image[15][7])} + {7'd0,(kernel[4][3] ~^ image[15][8])} + {7'd0,(kernel[4][4] ~^ image[15][9])};
assign out_fmap[11][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[11][6])} + {7'd0,(kernel[0][1] ~^ image[11][7])} + {7'd0,(kernel[0][2] ~^ image[11][8])} + {7'd0,(kernel[0][3] ~^ image[11][9])} + {7'd0,(kernel[0][4] ~^ image[11][10])} + {7'd0,(kernel[1][0] ~^ image[12][6])} + {7'd0,(kernel[1][1] ~^ image[12][7])} + {7'd0,(kernel[1][2] ~^ image[12][8])} + {7'd0,(kernel[1][3] ~^ image[12][9])} + {7'd0,(kernel[1][4] ~^ image[12][10])} + {7'd0,(kernel[2][0] ~^ image[13][6])} + {7'd0,(kernel[2][1] ~^ image[13][7])} + {7'd0,(kernel[2][2] ~^ image[13][8])} + {7'd0,(kernel[2][3] ~^ image[13][9])} + {7'd0,(kernel[2][4] ~^ image[13][10])} + {7'd0,(kernel[3][0] ~^ image[14][6])} + {7'd0,(kernel[3][1] ~^ image[14][7])} + {7'd0,(kernel[3][2] ~^ image[14][8])} + {7'd0,(kernel[3][3] ~^ image[14][9])} + {7'd0,(kernel[3][4] ~^ image[14][10])} + {7'd0,(kernel[4][0] ~^ image[15][6])} + {7'd0,(kernel[4][1] ~^ image[15][7])} + {7'd0,(kernel[4][2] ~^ image[15][8])} + {7'd0,(kernel[4][3] ~^ image[15][9])} + {7'd0,(kernel[4][4] ~^ image[15][10])};
assign out_fmap[11][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[11][7])} + {7'd0,(kernel[0][1] ~^ image[11][8])} + {7'd0,(kernel[0][2] ~^ image[11][9])} + {7'd0,(kernel[0][3] ~^ image[11][10])} + {7'd0,(kernel[0][4] ~^ image[11][11])} + {7'd0,(kernel[1][0] ~^ image[12][7])} + {7'd0,(kernel[1][1] ~^ image[12][8])} + {7'd0,(kernel[1][2] ~^ image[12][9])} + {7'd0,(kernel[1][3] ~^ image[12][10])} + {7'd0,(kernel[1][4] ~^ image[12][11])} + {7'd0,(kernel[2][0] ~^ image[13][7])} + {7'd0,(kernel[2][1] ~^ image[13][8])} + {7'd0,(kernel[2][2] ~^ image[13][9])} + {7'd0,(kernel[2][3] ~^ image[13][10])} + {7'd0,(kernel[2][4] ~^ image[13][11])} + {7'd0,(kernel[3][0] ~^ image[14][7])} + {7'd0,(kernel[3][1] ~^ image[14][8])} + {7'd0,(kernel[3][2] ~^ image[14][9])} + {7'd0,(kernel[3][3] ~^ image[14][10])} + {7'd0,(kernel[3][4] ~^ image[14][11])} + {7'd0,(kernel[4][0] ~^ image[15][7])} + {7'd0,(kernel[4][1] ~^ image[15][8])} + {7'd0,(kernel[4][2] ~^ image[15][9])} + {7'd0,(kernel[4][3] ~^ image[15][10])} + {7'd0,(kernel[4][4] ~^ image[15][11])};
assign out_fmap[11][8][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[11][8])} + {7'd0,(kernel[0][1] ~^ image[11][9])} + {7'd0,(kernel[0][2] ~^ image[11][10])} + {7'd0,(kernel[0][3] ~^ image[11][11])} + {7'd0,(kernel[0][4] ~^ image[11][12])} + {7'd0,(kernel[1][0] ~^ image[12][8])} + {7'd0,(kernel[1][1] ~^ image[12][9])} + {7'd0,(kernel[1][2] ~^ image[12][10])} + {7'd0,(kernel[1][3] ~^ image[12][11])} + {7'd0,(kernel[1][4] ~^ image[12][12])} + {7'd0,(kernel[2][0] ~^ image[13][8])} + {7'd0,(kernel[2][1] ~^ image[13][9])} + {7'd0,(kernel[2][2] ~^ image[13][10])} + {7'd0,(kernel[2][3] ~^ image[13][11])} + {7'd0,(kernel[2][4] ~^ image[13][12])} + {7'd0,(kernel[3][0] ~^ image[14][8])} + {7'd0,(kernel[3][1] ~^ image[14][9])} + {7'd0,(kernel[3][2] ~^ image[14][10])} + {7'd0,(kernel[3][3] ~^ image[14][11])} + {7'd0,(kernel[3][4] ~^ image[14][12])} + {7'd0,(kernel[4][0] ~^ image[15][8])} + {7'd0,(kernel[4][1] ~^ image[15][9])} + {7'd0,(kernel[4][2] ~^ image[15][10])} + {7'd0,(kernel[4][3] ~^ image[15][11])} + {7'd0,(kernel[4][4] ~^ image[15][12])};
assign out_fmap[11][9][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[11][9])} + {7'd0,(kernel[0][1] ~^ image[11][10])} + {7'd0,(kernel[0][2] ~^ image[11][11])} + {7'd0,(kernel[0][3] ~^ image[11][12])} + {7'd0,(kernel[0][4] ~^ image[11][13])} + {7'd0,(kernel[1][0] ~^ image[12][9])} + {7'd0,(kernel[1][1] ~^ image[12][10])} + {7'd0,(kernel[1][2] ~^ image[12][11])} + {7'd0,(kernel[1][3] ~^ image[12][12])} + {7'd0,(kernel[1][4] ~^ image[12][13])} + {7'd0,(kernel[2][0] ~^ image[13][9])} + {7'd0,(kernel[2][1] ~^ image[13][10])} + {7'd0,(kernel[2][2] ~^ image[13][11])} + {7'd0,(kernel[2][3] ~^ image[13][12])} + {7'd0,(kernel[2][4] ~^ image[13][13])} + {7'd0,(kernel[3][0] ~^ image[14][9])} + {7'd0,(kernel[3][1] ~^ image[14][10])} + {7'd0,(kernel[3][2] ~^ image[14][11])} + {7'd0,(kernel[3][3] ~^ image[14][12])} + {7'd0,(kernel[3][4] ~^ image[14][13])} + {7'd0,(kernel[4][0] ~^ image[15][9])} + {7'd0,(kernel[4][1] ~^ image[15][10])} + {7'd0,(kernel[4][2] ~^ image[15][11])} + {7'd0,(kernel[4][3] ~^ image[15][12])} + {7'd0,(kernel[4][4] ~^ image[15][13])};
assign out_fmap[11][10][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[11][10])} + {7'd0,(kernel[0][1] ~^ image[11][11])} + {7'd0,(kernel[0][2] ~^ image[11][12])} + {7'd0,(kernel[0][3] ~^ image[11][13])} + {7'd0,(kernel[0][4] ~^ image[11][14])} + {7'd0,(kernel[1][0] ~^ image[12][10])} + {7'd0,(kernel[1][1] ~^ image[12][11])} + {7'd0,(kernel[1][2] ~^ image[12][12])} + {7'd0,(kernel[1][3] ~^ image[12][13])} + {7'd0,(kernel[1][4] ~^ image[12][14])} + {7'd0,(kernel[2][0] ~^ image[13][10])} + {7'd0,(kernel[2][1] ~^ image[13][11])} + {7'd0,(kernel[2][2] ~^ image[13][12])} + {7'd0,(kernel[2][3] ~^ image[13][13])} + {7'd0,(kernel[2][4] ~^ image[13][14])} + {7'd0,(kernel[3][0] ~^ image[14][10])} + {7'd0,(kernel[3][1] ~^ image[14][11])} + {7'd0,(kernel[3][2] ~^ image[14][12])} + {7'd0,(kernel[3][3] ~^ image[14][13])} + {7'd0,(kernel[3][4] ~^ image[14][14])} + {7'd0,(kernel[4][0] ~^ image[15][10])} + {7'd0,(kernel[4][1] ~^ image[15][11])} + {7'd0,(kernel[4][2] ~^ image[15][12])} + {7'd0,(kernel[4][3] ~^ image[15][13])} + {7'd0,(kernel[4][4] ~^ image[15][14])};
assign out_fmap[11][11][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[11][11])} + {7'd0,(kernel[0][1] ~^ image[11][12])} + {7'd0,(kernel[0][2] ~^ image[11][13])} + {7'd0,(kernel[0][3] ~^ image[11][14])} + {7'd0,(kernel[0][4] ~^ image[11][15])} + {7'd0,(kernel[1][0] ~^ image[12][11])} + {7'd0,(kernel[1][1] ~^ image[12][12])} + {7'd0,(kernel[1][2] ~^ image[12][13])} + {7'd0,(kernel[1][3] ~^ image[12][14])} + {7'd0,(kernel[1][4] ~^ image[12][15])} + {7'd0,(kernel[2][0] ~^ image[13][11])} + {7'd0,(kernel[2][1] ~^ image[13][12])} + {7'd0,(kernel[2][2] ~^ image[13][13])} + {7'd0,(kernel[2][3] ~^ image[13][14])} + {7'd0,(kernel[2][4] ~^ image[13][15])} + {7'd0,(kernel[3][0] ~^ image[14][11])} + {7'd0,(kernel[3][1] ~^ image[14][12])} + {7'd0,(kernel[3][2] ~^ image[14][13])} + {7'd0,(kernel[3][3] ~^ image[14][14])} + {7'd0,(kernel[3][4] ~^ image[14][15])} + {7'd0,(kernel[4][0] ~^ image[15][11])} + {7'd0,(kernel[4][1] ~^ image[15][12])} + {7'd0,(kernel[4][2] ~^ image[15][13])} + {7'd0,(kernel[4][3] ~^ image[15][14])} + {7'd0,(kernel[4][4] ~^ image[15][15])};
assign out_fmap[11][12][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[11][12])} + {7'd0,(kernel[0][1] ~^ image[11][13])} + {7'd0,(kernel[0][2] ~^ image[11][14])} + {7'd0,(kernel[0][3] ~^ image[11][15])} + {7'd0,(kernel[0][4] ~^ image[11][16])} + {7'd0,(kernel[1][0] ~^ image[12][12])} + {7'd0,(kernel[1][1] ~^ image[12][13])} + {7'd0,(kernel[1][2] ~^ image[12][14])} + {7'd0,(kernel[1][3] ~^ image[12][15])} + {7'd0,(kernel[1][4] ~^ image[12][16])} + {7'd0,(kernel[2][0] ~^ image[13][12])} + {7'd0,(kernel[2][1] ~^ image[13][13])} + {7'd0,(kernel[2][2] ~^ image[13][14])} + {7'd0,(kernel[2][3] ~^ image[13][15])} + {7'd0,(kernel[2][4] ~^ image[13][16])} + {7'd0,(kernel[3][0] ~^ image[14][12])} + {7'd0,(kernel[3][1] ~^ image[14][13])} + {7'd0,(kernel[3][2] ~^ image[14][14])} + {7'd0,(kernel[3][3] ~^ image[14][15])} + {7'd0,(kernel[3][4] ~^ image[14][16])} + {7'd0,(kernel[4][0] ~^ image[15][12])} + {7'd0,(kernel[4][1] ~^ image[15][13])} + {7'd0,(kernel[4][2] ~^ image[15][14])} + {7'd0,(kernel[4][3] ~^ image[15][15])} + {7'd0,(kernel[4][4] ~^ image[15][16])};
assign out_fmap[11][13][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[11][13])} + {7'd0,(kernel[0][1] ~^ image[11][14])} + {7'd0,(kernel[0][2] ~^ image[11][15])} + {7'd0,(kernel[0][3] ~^ image[11][16])} + {7'd0,(kernel[0][4] ~^ image[11][17])} + {7'd0,(kernel[1][0] ~^ image[12][13])} + {7'd0,(kernel[1][1] ~^ image[12][14])} + {7'd0,(kernel[1][2] ~^ image[12][15])} + {7'd0,(kernel[1][3] ~^ image[12][16])} + {7'd0,(kernel[1][4] ~^ image[12][17])} + {7'd0,(kernel[2][0] ~^ image[13][13])} + {7'd0,(kernel[2][1] ~^ image[13][14])} + {7'd0,(kernel[2][2] ~^ image[13][15])} + {7'd0,(kernel[2][3] ~^ image[13][16])} + {7'd0,(kernel[2][4] ~^ image[13][17])} + {7'd0,(kernel[3][0] ~^ image[14][13])} + {7'd0,(kernel[3][1] ~^ image[14][14])} + {7'd0,(kernel[3][2] ~^ image[14][15])} + {7'd0,(kernel[3][3] ~^ image[14][16])} + {7'd0,(kernel[3][4] ~^ image[14][17])} + {7'd0,(kernel[4][0] ~^ image[15][13])} + {7'd0,(kernel[4][1] ~^ image[15][14])} + {7'd0,(kernel[4][2] ~^ image[15][15])} + {7'd0,(kernel[4][3] ~^ image[15][16])} + {7'd0,(kernel[4][4] ~^ image[15][17])};
assign out_fmap[11][14][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[11][14])} + {7'd0,(kernel[0][1] ~^ image[11][15])} + {7'd0,(kernel[0][2] ~^ image[11][16])} + {7'd0,(kernel[0][3] ~^ image[11][17])} + {7'd0,(kernel[0][4] ~^ image[11][18])} + {7'd0,(kernel[1][0] ~^ image[12][14])} + {7'd0,(kernel[1][1] ~^ image[12][15])} + {7'd0,(kernel[1][2] ~^ image[12][16])} + {7'd0,(kernel[1][3] ~^ image[12][17])} + {7'd0,(kernel[1][4] ~^ image[12][18])} + {7'd0,(kernel[2][0] ~^ image[13][14])} + {7'd0,(kernel[2][1] ~^ image[13][15])} + {7'd0,(kernel[2][2] ~^ image[13][16])} + {7'd0,(kernel[2][3] ~^ image[13][17])} + {7'd0,(kernel[2][4] ~^ image[13][18])} + {7'd0,(kernel[3][0] ~^ image[14][14])} + {7'd0,(kernel[3][1] ~^ image[14][15])} + {7'd0,(kernel[3][2] ~^ image[14][16])} + {7'd0,(kernel[3][3] ~^ image[14][17])} + {7'd0,(kernel[3][4] ~^ image[14][18])} + {7'd0,(kernel[4][0] ~^ image[15][14])} + {7'd0,(kernel[4][1] ~^ image[15][15])} + {7'd0,(kernel[4][2] ~^ image[15][16])} + {7'd0,(kernel[4][3] ~^ image[15][17])} + {7'd0,(kernel[4][4] ~^ image[15][18])};
assign out_fmap[11][15][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[11][15])} + {7'd0,(kernel[0][1] ~^ image[11][16])} + {7'd0,(kernel[0][2] ~^ image[11][17])} + {7'd0,(kernel[0][3] ~^ image[11][18])} + {7'd0,(kernel[0][4] ~^ image[11][19])} + {7'd0,(kernel[1][0] ~^ image[12][15])} + {7'd0,(kernel[1][1] ~^ image[12][16])} + {7'd0,(kernel[1][2] ~^ image[12][17])} + {7'd0,(kernel[1][3] ~^ image[12][18])} + {7'd0,(kernel[1][4] ~^ image[12][19])} + {7'd0,(kernel[2][0] ~^ image[13][15])} + {7'd0,(kernel[2][1] ~^ image[13][16])} + {7'd0,(kernel[2][2] ~^ image[13][17])} + {7'd0,(kernel[2][3] ~^ image[13][18])} + {7'd0,(kernel[2][4] ~^ image[13][19])} + {7'd0,(kernel[3][0] ~^ image[14][15])} + {7'd0,(kernel[3][1] ~^ image[14][16])} + {7'd0,(kernel[3][2] ~^ image[14][17])} + {7'd0,(kernel[3][3] ~^ image[14][18])} + {7'd0,(kernel[3][4] ~^ image[14][19])} + {7'd0,(kernel[4][0] ~^ image[15][15])} + {7'd0,(kernel[4][1] ~^ image[15][16])} + {7'd0,(kernel[4][2] ~^ image[15][17])} + {7'd0,(kernel[4][3] ~^ image[15][18])} + {7'd0,(kernel[4][4] ~^ image[15][19])};
assign out_fmap[11][16][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[11][16])} + {7'd0,(kernel[0][1] ~^ image[11][17])} + {7'd0,(kernel[0][2] ~^ image[11][18])} + {7'd0,(kernel[0][3] ~^ image[11][19])} + {7'd0,(kernel[0][4] ~^ image[11][20])} + {7'd0,(kernel[1][0] ~^ image[12][16])} + {7'd0,(kernel[1][1] ~^ image[12][17])} + {7'd0,(kernel[1][2] ~^ image[12][18])} + {7'd0,(kernel[1][3] ~^ image[12][19])} + {7'd0,(kernel[1][4] ~^ image[12][20])} + {7'd0,(kernel[2][0] ~^ image[13][16])} + {7'd0,(kernel[2][1] ~^ image[13][17])} + {7'd0,(kernel[2][2] ~^ image[13][18])} + {7'd0,(kernel[2][3] ~^ image[13][19])} + {7'd0,(kernel[2][4] ~^ image[13][20])} + {7'd0,(kernel[3][0] ~^ image[14][16])} + {7'd0,(kernel[3][1] ~^ image[14][17])} + {7'd0,(kernel[3][2] ~^ image[14][18])} + {7'd0,(kernel[3][3] ~^ image[14][19])} + {7'd0,(kernel[3][4] ~^ image[14][20])} + {7'd0,(kernel[4][0] ~^ image[15][16])} + {7'd0,(kernel[4][1] ~^ image[15][17])} + {7'd0,(kernel[4][2] ~^ image[15][18])} + {7'd0,(kernel[4][3] ~^ image[15][19])} + {7'd0,(kernel[4][4] ~^ image[15][20])};
assign out_fmap[11][17][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[11][17])} + {7'd0,(kernel[0][1] ~^ image[11][18])} + {7'd0,(kernel[0][2] ~^ image[11][19])} + {7'd0,(kernel[0][3] ~^ image[11][20])} + {7'd0,(kernel[0][4] ~^ image[11][21])} + {7'd0,(kernel[1][0] ~^ image[12][17])} + {7'd0,(kernel[1][1] ~^ image[12][18])} + {7'd0,(kernel[1][2] ~^ image[12][19])} + {7'd0,(kernel[1][3] ~^ image[12][20])} + {7'd0,(kernel[1][4] ~^ image[12][21])} + {7'd0,(kernel[2][0] ~^ image[13][17])} + {7'd0,(kernel[2][1] ~^ image[13][18])} + {7'd0,(kernel[2][2] ~^ image[13][19])} + {7'd0,(kernel[2][3] ~^ image[13][20])} + {7'd0,(kernel[2][4] ~^ image[13][21])} + {7'd0,(kernel[3][0] ~^ image[14][17])} + {7'd0,(kernel[3][1] ~^ image[14][18])} + {7'd0,(kernel[3][2] ~^ image[14][19])} + {7'd0,(kernel[3][3] ~^ image[14][20])} + {7'd0,(kernel[3][4] ~^ image[14][21])} + {7'd0,(kernel[4][0] ~^ image[15][17])} + {7'd0,(kernel[4][1] ~^ image[15][18])} + {7'd0,(kernel[4][2] ~^ image[15][19])} + {7'd0,(kernel[4][3] ~^ image[15][20])} + {7'd0,(kernel[4][4] ~^ image[15][21])};
assign out_fmap[11][18][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[11][18])} + {7'd0,(kernel[0][1] ~^ image[11][19])} + {7'd0,(kernel[0][2] ~^ image[11][20])} + {7'd0,(kernel[0][3] ~^ image[11][21])} + {7'd0,(kernel[0][4] ~^ image[11][22])} + {7'd0,(kernel[1][0] ~^ image[12][18])} + {7'd0,(kernel[1][1] ~^ image[12][19])} + {7'd0,(kernel[1][2] ~^ image[12][20])} + {7'd0,(kernel[1][3] ~^ image[12][21])} + {7'd0,(kernel[1][4] ~^ image[12][22])} + {7'd0,(kernel[2][0] ~^ image[13][18])} + {7'd0,(kernel[2][1] ~^ image[13][19])} + {7'd0,(kernel[2][2] ~^ image[13][20])} + {7'd0,(kernel[2][3] ~^ image[13][21])} + {7'd0,(kernel[2][4] ~^ image[13][22])} + {7'd0,(kernel[3][0] ~^ image[14][18])} + {7'd0,(kernel[3][1] ~^ image[14][19])} + {7'd0,(kernel[3][2] ~^ image[14][20])} + {7'd0,(kernel[3][3] ~^ image[14][21])} + {7'd0,(kernel[3][4] ~^ image[14][22])} + {7'd0,(kernel[4][0] ~^ image[15][18])} + {7'd0,(kernel[4][1] ~^ image[15][19])} + {7'd0,(kernel[4][2] ~^ image[15][20])} + {7'd0,(kernel[4][3] ~^ image[15][21])} + {7'd0,(kernel[4][4] ~^ image[15][22])};
assign out_fmap[11][19][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[11][19])} + {7'd0,(kernel[0][1] ~^ image[11][20])} + {7'd0,(kernel[0][2] ~^ image[11][21])} + {7'd0,(kernel[0][3] ~^ image[11][22])} + {7'd0,(kernel[0][4] ~^ image[11][23])} + {7'd0,(kernel[1][0] ~^ image[12][19])} + {7'd0,(kernel[1][1] ~^ image[12][20])} + {7'd0,(kernel[1][2] ~^ image[12][21])} + {7'd0,(kernel[1][3] ~^ image[12][22])} + {7'd0,(kernel[1][4] ~^ image[12][23])} + {7'd0,(kernel[2][0] ~^ image[13][19])} + {7'd0,(kernel[2][1] ~^ image[13][20])} + {7'd0,(kernel[2][2] ~^ image[13][21])} + {7'd0,(kernel[2][3] ~^ image[13][22])} + {7'd0,(kernel[2][4] ~^ image[13][23])} + {7'd0,(kernel[3][0] ~^ image[14][19])} + {7'd0,(kernel[3][1] ~^ image[14][20])} + {7'd0,(kernel[3][2] ~^ image[14][21])} + {7'd0,(kernel[3][3] ~^ image[14][22])} + {7'd0,(kernel[3][4] ~^ image[14][23])} + {7'd0,(kernel[4][0] ~^ image[15][19])} + {7'd0,(kernel[4][1] ~^ image[15][20])} + {7'd0,(kernel[4][2] ~^ image[15][21])} + {7'd0,(kernel[4][3] ~^ image[15][22])} + {7'd0,(kernel[4][4] ~^ image[15][23])};
assign out_fmap[11][20][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[11][20])} + {7'd0,(kernel[0][1] ~^ image[11][21])} + {7'd0,(kernel[0][2] ~^ image[11][22])} + {7'd0,(kernel[0][3] ~^ image[11][23])} + {7'd0,(kernel[0][4] ~^ image[11][24])} + {7'd0,(kernel[1][0] ~^ image[12][20])} + {7'd0,(kernel[1][1] ~^ image[12][21])} + {7'd0,(kernel[1][2] ~^ image[12][22])} + {7'd0,(kernel[1][3] ~^ image[12][23])} + {7'd0,(kernel[1][4] ~^ image[12][24])} + {7'd0,(kernel[2][0] ~^ image[13][20])} + {7'd0,(kernel[2][1] ~^ image[13][21])} + {7'd0,(kernel[2][2] ~^ image[13][22])} + {7'd0,(kernel[2][3] ~^ image[13][23])} + {7'd0,(kernel[2][4] ~^ image[13][24])} + {7'd0,(kernel[3][0] ~^ image[14][20])} + {7'd0,(kernel[3][1] ~^ image[14][21])} + {7'd0,(kernel[3][2] ~^ image[14][22])} + {7'd0,(kernel[3][3] ~^ image[14][23])} + {7'd0,(kernel[3][4] ~^ image[14][24])} + {7'd0,(kernel[4][0] ~^ image[15][20])} + {7'd0,(kernel[4][1] ~^ image[15][21])} + {7'd0,(kernel[4][2] ~^ image[15][22])} + {7'd0,(kernel[4][3] ~^ image[15][23])} + {7'd0,(kernel[4][4] ~^ image[15][24])};
assign out_fmap[11][21][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[11][21])} + {7'd0,(kernel[0][1] ~^ image[11][22])} + {7'd0,(kernel[0][2] ~^ image[11][23])} + {7'd0,(kernel[0][3] ~^ image[11][24])} + {7'd0,(kernel[0][4] ~^ image[11][25])} + {7'd0,(kernel[1][0] ~^ image[12][21])} + {7'd0,(kernel[1][1] ~^ image[12][22])} + {7'd0,(kernel[1][2] ~^ image[12][23])} + {7'd0,(kernel[1][3] ~^ image[12][24])} + {7'd0,(kernel[1][4] ~^ image[12][25])} + {7'd0,(kernel[2][0] ~^ image[13][21])} + {7'd0,(kernel[2][1] ~^ image[13][22])} + {7'd0,(kernel[2][2] ~^ image[13][23])} + {7'd0,(kernel[2][3] ~^ image[13][24])} + {7'd0,(kernel[2][4] ~^ image[13][25])} + {7'd0,(kernel[3][0] ~^ image[14][21])} + {7'd0,(kernel[3][1] ~^ image[14][22])} + {7'd0,(kernel[3][2] ~^ image[14][23])} + {7'd0,(kernel[3][3] ~^ image[14][24])} + {7'd0,(kernel[3][4] ~^ image[14][25])} + {7'd0,(kernel[4][0] ~^ image[15][21])} + {7'd0,(kernel[4][1] ~^ image[15][22])} + {7'd0,(kernel[4][2] ~^ image[15][23])} + {7'd0,(kernel[4][3] ~^ image[15][24])} + {7'd0,(kernel[4][4] ~^ image[15][25])};
assign out_fmap[11][22][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[11][22])} + {7'd0,(kernel[0][1] ~^ image[11][23])} + {7'd0,(kernel[0][2] ~^ image[11][24])} + {7'd0,(kernel[0][3] ~^ image[11][25])} + {7'd0,(kernel[0][4] ~^ image[11][26])} + {7'd0,(kernel[1][0] ~^ image[12][22])} + {7'd0,(kernel[1][1] ~^ image[12][23])} + {7'd0,(kernel[1][2] ~^ image[12][24])} + {7'd0,(kernel[1][3] ~^ image[12][25])} + {7'd0,(kernel[1][4] ~^ image[12][26])} + {7'd0,(kernel[2][0] ~^ image[13][22])} + {7'd0,(kernel[2][1] ~^ image[13][23])} + {7'd0,(kernel[2][2] ~^ image[13][24])} + {7'd0,(kernel[2][3] ~^ image[13][25])} + {7'd0,(kernel[2][4] ~^ image[13][26])} + {7'd0,(kernel[3][0] ~^ image[14][22])} + {7'd0,(kernel[3][1] ~^ image[14][23])} + {7'd0,(kernel[3][2] ~^ image[14][24])} + {7'd0,(kernel[3][3] ~^ image[14][25])} + {7'd0,(kernel[3][4] ~^ image[14][26])} + {7'd0,(kernel[4][0] ~^ image[15][22])} + {7'd0,(kernel[4][1] ~^ image[15][23])} + {7'd0,(kernel[4][2] ~^ image[15][24])} + {7'd0,(kernel[4][3] ~^ image[15][25])} + {7'd0,(kernel[4][4] ~^ image[15][26])};
assign out_fmap[11][23][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[11][23])} + {7'd0,(kernel[0][1] ~^ image[11][24])} + {7'd0,(kernel[0][2] ~^ image[11][25])} + {7'd0,(kernel[0][3] ~^ image[11][26])} + {7'd0,(kernel[0][4] ~^ image[11][27])} + {7'd0,(kernel[1][0] ~^ image[12][23])} + {7'd0,(kernel[1][1] ~^ image[12][24])} + {7'd0,(kernel[1][2] ~^ image[12][25])} + {7'd0,(kernel[1][3] ~^ image[12][26])} + {7'd0,(kernel[1][4] ~^ image[12][27])} + {7'd0,(kernel[2][0] ~^ image[13][23])} + {7'd0,(kernel[2][1] ~^ image[13][24])} + {7'd0,(kernel[2][2] ~^ image[13][25])} + {7'd0,(kernel[2][3] ~^ image[13][26])} + {7'd0,(kernel[2][4] ~^ image[13][27])} + {7'd0,(kernel[3][0] ~^ image[14][23])} + {7'd0,(kernel[3][1] ~^ image[14][24])} + {7'd0,(kernel[3][2] ~^ image[14][25])} + {7'd0,(kernel[3][3] ~^ image[14][26])} + {7'd0,(kernel[3][4] ~^ image[14][27])} + {7'd0,(kernel[4][0] ~^ image[15][23])} + {7'd0,(kernel[4][1] ~^ image[15][24])} + {7'd0,(kernel[4][2] ~^ image[15][25])} + {7'd0,(kernel[4][3] ~^ image[15][26])} + {7'd0,(kernel[4][4] ~^ image[15][27])};
assign out_fmap[12][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[12][0])} + {7'd0,(kernel[0][1] ~^ image[12][1])} + {7'd0,(kernel[0][2] ~^ image[12][2])} + {7'd0,(kernel[0][3] ~^ image[12][3])} + {7'd0,(kernel[0][4] ~^ image[12][4])} + {7'd0,(kernel[1][0] ~^ image[13][0])} + {7'd0,(kernel[1][1] ~^ image[13][1])} + {7'd0,(kernel[1][2] ~^ image[13][2])} + {7'd0,(kernel[1][3] ~^ image[13][3])} + {7'd0,(kernel[1][4] ~^ image[13][4])} + {7'd0,(kernel[2][0] ~^ image[14][0])} + {7'd0,(kernel[2][1] ~^ image[14][1])} + {7'd0,(kernel[2][2] ~^ image[14][2])} + {7'd0,(kernel[2][3] ~^ image[14][3])} + {7'd0,(kernel[2][4] ~^ image[14][4])} + {7'd0,(kernel[3][0] ~^ image[15][0])} + {7'd0,(kernel[3][1] ~^ image[15][1])} + {7'd0,(kernel[3][2] ~^ image[15][2])} + {7'd0,(kernel[3][3] ~^ image[15][3])} + {7'd0,(kernel[3][4] ~^ image[15][4])} + {7'd0,(kernel[4][0] ~^ image[16][0])} + {7'd0,(kernel[4][1] ~^ image[16][1])} + {7'd0,(kernel[4][2] ~^ image[16][2])} + {7'd0,(kernel[4][3] ~^ image[16][3])} + {7'd0,(kernel[4][4] ~^ image[16][4])};
assign out_fmap[12][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[12][1])} + {7'd0,(kernel[0][1] ~^ image[12][2])} + {7'd0,(kernel[0][2] ~^ image[12][3])} + {7'd0,(kernel[0][3] ~^ image[12][4])} + {7'd0,(kernel[0][4] ~^ image[12][5])} + {7'd0,(kernel[1][0] ~^ image[13][1])} + {7'd0,(kernel[1][1] ~^ image[13][2])} + {7'd0,(kernel[1][2] ~^ image[13][3])} + {7'd0,(kernel[1][3] ~^ image[13][4])} + {7'd0,(kernel[1][4] ~^ image[13][5])} + {7'd0,(kernel[2][0] ~^ image[14][1])} + {7'd0,(kernel[2][1] ~^ image[14][2])} + {7'd0,(kernel[2][2] ~^ image[14][3])} + {7'd0,(kernel[2][3] ~^ image[14][4])} + {7'd0,(kernel[2][4] ~^ image[14][5])} + {7'd0,(kernel[3][0] ~^ image[15][1])} + {7'd0,(kernel[3][1] ~^ image[15][2])} + {7'd0,(kernel[3][2] ~^ image[15][3])} + {7'd0,(kernel[3][3] ~^ image[15][4])} + {7'd0,(kernel[3][4] ~^ image[15][5])} + {7'd0,(kernel[4][0] ~^ image[16][1])} + {7'd0,(kernel[4][1] ~^ image[16][2])} + {7'd0,(kernel[4][2] ~^ image[16][3])} + {7'd0,(kernel[4][3] ~^ image[16][4])} + {7'd0,(kernel[4][4] ~^ image[16][5])};
assign out_fmap[12][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[12][2])} + {7'd0,(kernel[0][1] ~^ image[12][3])} + {7'd0,(kernel[0][2] ~^ image[12][4])} + {7'd0,(kernel[0][3] ~^ image[12][5])} + {7'd0,(kernel[0][4] ~^ image[12][6])} + {7'd0,(kernel[1][0] ~^ image[13][2])} + {7'd0,(kernel[1][1] ~^ image[13][3])} + {7'd0,(kernel[1][2] ~^ image[13][4])} + {7'd0,(kernel[1][3] ~^ image[13][5])} + {7'd0,(kernel[1][4] ~^ image[13][6])} + {7'd0,(kernel[2][0] ~^ image[14][2])} + {7'd0,(kernel[2][1] ~^ image[14][3])} + {7'd0,(kernel[2][2] ~^ image[14][4])} + {7'd0,(kernel[2][3] ~^ image[14][5])} + {7'd0,(kernel[2][4] ~^ image[14][6])} + {7'd0,(kernel[3][0] ~^ image[15][2])} + {7'd0,(kernel[3][1] ~^ image[15][3])} + {7'd0,(kernel[3][2] ~^ image[15][4])} + {7'd0,(kernel[3][3] ~^ image[15][5])} + {7'd0,(kernel[3][4] ~^ image[15][6])} + {7'd0,(kernel[4][0] ~^ image[16][2])} + {7'd0,(kernel[4][1] ~^ image[16][3])} + {7'd0,(kernel[4][2] ~^ image[16][4])} + {7'd0,(kernel[4][3] ~^ image[16][5])} + {7'd0,(kernel[4][4] ~^ image[16][6])};
assign out_fmap[12][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[12][3])} + {7'd0,(kernel[0][1] ~^ image[12][4])} + {7'd0,(kernel[0][2] ~^ image[12][5])} + {7'd0,(kernel[0][3] ~^ image[12][6])} + {7'd0,(kernel[0][4] ~^ image[12][7])} + {7'd0,(kernel[1][0] ~^ image[13][3])} + {7'd0,(kernel[1][1] ~^ image[13][4])} + {7'd0,(kernel[1][2] ~^ image[13][5])} + {7'd0,(kernel[1][3] ~^ image[13][6])} + {7'd0,(kernel[1][4] ~^ image[13][7])} + {7'd0,(kernel[2][0] ~^ image[14][3])} + {7'd0,(kernel[2][1] ~^ image[14][4])} + {7'd0,(kernel[2][2] ~^ image[14][5])} + {7'd0,(kernel[2][3] ~^ image[14][6])} + {7'd0,(kernel[2][4] ~^ image[14][7])} + {7'd0,(kernel[3][0] ~^ image[15][3])} + {7'd0,(kernel[3][1] ~^ image[15][4])} + {7'd0,(kernel[3][2] ~^ image[15][5])} + {7'd0,(kernel[3][3] ~^ image[15][6])} + {7'd0,(kernel[3][4] ~^ image[15][7])} + {7'd0,(kernel[4][0] ~^ image[16][3])} + {7'd0,(kernel[4][1] ~^ image[16][4])} + {7'd0,(kernel[4][2] ~^ image[16][5])} + {7'd0,(kernel[4][3] ~^ image[16][6])} + {7'd0,(kernel[4][4] ~^ image[16][7])};
assign out_fmap[12][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[12][4])} + {7'd0,(kernel[0][1] ~^ image[12][5])} + {7'd0,(kernel[0][2] ~^ image[12][6])} + {7'd0,(kernel[0][3] ~^ image[12][7])} + {7'd0,(kernel[0][4] ~^ image[12][8])} + {7'd0,(kernel[1][0] ~^ image[13][4])} + {7'd0,(kernel[1][1] ~^ image[13][5])} + {7'd0,(kernel[1][2] ~^ image[13][6])} + {7'd0,(kernel[1][3] ~^ image[13][7])} + {7'd0,(kernel[1][4] ~^ image[13][8])} + {7'd0,(kernel[2][0] ~^ image[14][4])} + {7'd0,(kernel[2][1] ~^ image[14][5])} + {7'd0,(kernel[2][2] ~^ image[14][6])} + {7'd0,(kernel[2][3] ~^ image[14][7])} + {7'd0,(kernel[2][4] ~^ image[14][8])} + {7'd0,(kernel[3][0] ~^ image[15][4])} + {7'd0,(kernel[3][1] ~^ image[15][5])} + {7'd0,(kernel[3][2] ~^ image[15][6])} + {7'd0,(kernel[3][3] ~^ image[15][7])} + {7'd0,(kernel[3][4] ~^ image[15][8])} + {7'd0,(kernel[4][0] ~^ image[16][4])} + {7'd0,(kernel[4][1] ~^ image[16][5])} + {7'd0,(kernel[4][2] ~^ image[16][6])} + {7'd0,(kernel[4][3] ~^ image[16][7])} + {7'd0,(kernel[4][4] ~^ image[16][8])};
assign out_fmap[12][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[12][5])} + {7'd0,(kernel[0][1] ~^ image[12][6])} + {7'd0,(kernel[0][2] ~^ image[12][7])} + {7'd0,(kernel[0][3] ~^ image[12][8])} + {7'd0,(kernel[0][4] ~^ image[12][9])} + {7'd0,(kernel[1][0] ~^ image[13][5])} + {7'd0,(kernel[1][1] ~^ image[13][6])} + {7'd0,(kernel[1][2] ~^ image[13][7])} + {7'd0,(kernel[1][3] ~^ image[13][8])} + {7'd0,(kernel[1][4] ~^ image[13][9])} + {7'd0,(kernel[2][0] ~^ image[14][5])} + {7'd0,(kernel[2][1] ~^ image[14][6])} + {7'd0,(kernel[2][2] ~^ image[14][7])} + {7'd0,(kernel[2][3] ~^ image[14][8])} + {7'd0,(kernel[2][4] ~^ image[14][9])} + {7'd0,(kernel[3][0] ~^ image[15][5])} + {7'd0,(kernel[3][1] ~^ image[15][6])} + {7'd0,(kernel[3][2] ~^ image[15][7])} + {7'd0,(kernel[3][3] ~^ image[15][8])} + {7'd0,(kernel[3][4] ~^ image[15][9])} + {7'd0,(kernel[4][0] ~^ image[16][5])} + {7'd0,(kernel[4][1] ~^ image[16][6])} + {7'd0,(kernel[4][2] ~^ image[16][7])} + {7'd0,(kernel[4][3] ~^ image[16][8])} + {7'd0,(kernel[4][4] ~^ image[16][9])};
assign out_fmap[12][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[12][6])} + {7'd0,(kernel[0][1] ~^ image[12][7])} + {7'd0,(kernel[0][2] ~^ image[12][8])} + {7'd0,(kernel[0][3] ~^ image[12][9])} + {7'd0,(kernel[0][4] ~^ image[12][10])} + {7'd0,(kernel[1][0] ~^ image[13][6])} + {7'd0,(kernel[1][1] ~^ image[13][7])} + {7'd0,(kernel[1][2] ~^ image[13][8])} + {7'd0,(kernel[1][3] ~^ image[13][9])} + {7'd0,(kernel[1][4] ~^ image[13][10])} + {7'd0,(kernel[2][0] ~^ image[14][6])} + {7'd0,(kernel[2][1] ~^ image[14][7])} + {7'd0,(kernel[2][2] ~^ image[14][8])} + {7'd0,(kernel[2][3] ~^ image[14][9])} + {7'd0,(kernel[2][4] ~^ image[14][10])} + {7'd0,(kernel[3][0] ~^ image[15][6])} + {7'd0,(kernel[3][1] ~^ image[15][7])} + {7'd0,(kernel[3][2] ~^ image[15][8])} + {7'd0,(kernel[3][3] ~^ image[15][9])} + {7'd0,(kernel[3][4] ~^ image[15][10])} + {7'd0,(kernel[4][0] ~^ image[16][6])} + {7'd0,(kernel[4][1] ~^ image[16][7])} + {7'd0,(kernel[4][2] ~^ image[16][8])} + {7'd0,(kernel[4][3] ~^ image[16][9])} + {7'd0,(kernel[4][4] ~^ image[16][10])};
assign out_fmap[12][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[12][7])} + {7'd0,(kernel[0][1] ~^ image[12][8])} + {7'd0,(kernel[0][2] ~^ image[12][9])} + {7'd0,(kernel[0][3] ~^ image[12][10])} + {7'd0,(kernel[0][4] ~^ image[12][11])} + {7'd0,(kernel[1][0] ~^ image[13][7])} + {7'd0,(kernel[1][1] ~^ image[13][8])} + {7'd0,(kernel[1][2] ~^ image[13][9])} + {7'd0,(kernel[1][3] ~^ image[13][10])} + {7'd0,(kernel[1][4] ~^ image[13][11])} + {7'd0,(kernel[2][0] ~^ image[14][7])} + {7'd0,(kernel[2][1] ~^ image[14][8])} + {7'd0,(kernel[2][2] ~^ image[14][9])} + {7'd0,(kernel[2][3] ~^ image[14][10])} + {7'd0,(kernel[2][4] ~^ image[14][11])} + {7'd0,(kernel[3][0] ~^ image[15][7])} + {7'd0,(kernel[3][1] ~^ image[15][8])} + {7'd0,(kernel[3][2] ~^ image[15][9])} + {7'd0,(kernel[3][3] ~^ image[15][10])} + {7'd0,(kernel[3][4] ~^ image[15][11])} + {7'd0,(kernel[4][0] ~^ image[16][7])} + {7'd0,(kernel[4][1] ~^ image[16][8])} + {7'd0,(kernel[4][2] ~^ image[16][9])} + {7'd0,(kernel[4][3] ~^ image[16][10])} + {7'd0,(kernel[4][4] ~^ image[16][11])};
assign out_fmap[12][8][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[12][8])} + {7'd0,(kernel[0][1] ~^ image[12][9])} + {7'd0,(kernel[0][2] ~^ image[12][10])} + {7'd0,(kernel[0][3] ~^ image[12][11])} + {7'd0,(kernel[0][4] ~^ image[12][12])} + {7'd0,(kernel[1][0] ~^ image[13][8])} + {7'd0,(kernel[1][1] ~^ image[13][9])} + {7'd0,(kernel[1][2] ~^ image[13][10])} + {7'd0,(kernel[1][3] ~^ image[13][11])} + {7'd0,(kernel[1][4] ~^ image[13][12])} + {7'd0,(kernel[2][0] ~^ image[14][8])} + {7'd0,(kernel[2][1] ~^ image[14][9])} + {7'd0,(kernel[2][2] ~^ image[14][10])} + {7'd0,(kernel[2][3] ~^ image[14][11])} + {7'd0,(kernel[2][4] ~^ image[14][12])} + {7'd0,(kernel[3][0] ~^ image[15][8])} + {7'd0,(kernel[3][1] ~^ image[15][9])} + {7'd0,(kernel[3][2] ~^ image[15][10])} + {7'd0,(kernel[3][3] ~^ image[15][11])} + {7'd0,(kernel[3][4] ~^ image[15][12])} + {7'd0,(kernel[4][0] ~^ image[16][8])} + {7'd0,(kernel[4][1] ~^ image[16][9])} + {7'd0,(kernel[4][2] ~^ image[16][10])} + {7'd0,(kernel[4][3] ~^ image[16][11])} + {7'd0,(kernel[4][4] ~^ image[16][12])};
assign out_fmap[12][9][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[12][9])} + {7'd0,(kernel[0][1] ~^ image[12][10])} + {7'd0,(kernel[0][2] ~^ image[12][11])} + {7'd0,(kernel[0][3] ~^ image[12][12])} + {7'd0,(kernel[0][4] ~^ image[12][13])} + {7'd0,(kernel[1][0] ~^ image[13][9])} + {7'd0,(kernel[1][1] ~^ image[13][10])} + {7'd0,(kernel[1][2] ~^ image[13][11])} + {7'd0,(kernel[1][3] ~^ image[13][12])} + {7'd0,(kernel[1][4] ~^ image[13][13])} + {7'd0,(kernel[2][0] ~^ image[14][9])} + {7'd0,(kernel[2][1] ~^ image[14][10])} + {7'd0,(kernel[2][2] ~^ image[14][11])} + {7'd0,(kernel[2][3] ~^ image[14][12])} + {7'd0,(kernel[2][4] ~^ image[14][13])} + {7'd0,(kernel[3][0] ~^ image[15][9])} + {7'd0,(kernel[3][1] ~^ image[15][10])} + {7'd0,(kernel[3][2] ~^ image[15][11])} + {7'd0,(kernel[3][3] ~^ image[15][12])} + {7'd0,(kernel[3][4] ~^ image[15][13])} + {7'd0,(kernel[4][0] ~^ image[16][9])} + {7'd0,(kernel[4][1] ~^ image[16][10])} + {7'd0,(kernel[4][2] ~^ image[16][11])} + {7'd0,(kernel[4][3] ~^ image[16][12])} + {7'd0,(kernel[4][4] ~^ image[16][13])};
assign out_fmap[12][10][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[12][10])} + {7'd0,(kernel[0][1] ~^ image[12][11])} + {7'd0,(kernel[0][2] ~^ image[12][12])} + {7'd0,(kernel[0][3] ~^ image[12][13])} + {7'd0,(kernel[0][4] ~^ image[12][14])} + {7'd0,(kernel[1][0] ~^ image[13][10])} + {7'd0,(kernel[1][1] ~^ image[13][11])} + {7'd0,(kernel[1][2] ~^ image[13][12])} + {7'd0,(kernel[1][3] ~^ image[13][13])} + {7'd0,(kernel[1][4] ~^ image[13][14])} + {7'd0,(kernel[2][0] ~^ image[14][10])} + {7'd0,(kernel[2][1] ~^ image[14][11])} + {7'd0,(kernel[2][2] ~^ image[14][12])} + {7'd0,(kernel[2][3] ~^ image[14][13])} + {7'd0,(kernel[2][4] ~^ image[14][14])} + {7'd0,(kernel[3][0] ~^ image[15][10])} + {7'd0,(kernel[3][1] ~^ image[15][11])} + {7'd0,(kernel[3][2] ~^ image[15][12])} + {7'd0,(kernel[3][3] ~^ image[15][13])} + {7'd0,(kernel[3][4] ~^ image[15][14])} + {7'd0,(kernel[4][0] ~^ image[16][10])} + {7'd0,(kernel[4][1] ~^ image[16][11])} + {7'd0,(kernel[4][2] ~^ image[16][12])} + {7'd0,(kernel[4][3] ~^ image[16][13])} + {7'd0,(kernel[4][4] ~^ image[16][14])};
assign out_fmap[12][11][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[12][11])} + {7'd0,(kernel[0][1] ~^ image[12][12])} + {7'd0,(kernel[0][2] ~^ image[12][13])} + {7'd0,(kernel[0][3] ~^ image[12][14])} + {7'd0,(kernel[0][4] ~^ image[12][15])} + {7'd0,(kernel[1][0] ~^ image[13][11])} + {7'd0,(kernel[1][1] ~^ image[13][12])} + {7'd0,(kernel[1][2] ~^ image[13][13])} + {7'd0,(kernel[1][3] ~^ image[13][14])} + {7'd0,(kernel[1][4] ~^ image[13][15])} + {7'd0,(kernel[2][0] ~^ image[14][11])} + {7'd0,(kernel[2][1] ~^ image[14][12])} + {7'd0,(kernel[2][2] ~^ image[14][13])} + {7'd0,(kernel[2][3] ~^ image[14][14])} + {7'd0,(kernel[2][4] ~^ image[14][15])} + {7'd0,(kernel[3][0] ~^ image[15][11])} + {7'd0,(kernel[3][1] ~^ image[15][12])} + {7'd0,(kernel[3][2] ~^ image[15][13])} + {7'd0,(kernel[3][3] ~^ image[15][14])} + {7'd0,(kernel[3][4] ~^ image[15][15])} + {7'd0,(kernel[4][0] ~^ image[16][11])} + {7'd0,(kernel[4][1] ~^ image[16][12])} + {7'd0,(kernel[4][2] ~^ image[16][13])} + {7'd0,(kernel[4][3] ~^ image[16][14])} + {7'd0,(kernel[4][4] ~^ image[16][15])};
assign out_fmap[12][12][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[12][12])} + {7'd0,(kernel[0][1] ~^ image[12][13])} + {7'd0,(kernel[0][2] ~^ image[12][14])} + {7'd0,(kernel[0][3] ~^ image[12][15])} + {7'd0,(kernel[0][4] ~^ image[12][16])} + {7'd0,(kernel[1][0] ~^ image[13][12])} + {7'd0,(kernel[1][1] ~^ image[13][13])} + {7'd0,(kernel[1][2] ~^ image[13][14])} + {7'd0,(kernel[1][3] ~^ image[13][15])} + {7'd0,(kernel[1][4] ~^ image[13][16])} + {7'd0,(kernel[2][0] ~^ image[14][12])} + {7'd0,(kernel[2][1] ~^ image[14][13])} + {7'd0,(kernel[2][2] ~^ image[14][14])} + {7'd0,(kernel[2][3] ~^ image[14][15])} + {7'd0,(kernel[2][4] ~^ image[14][16])} + {7'd0,(kernel[3][0] ~^ image[15][12])} + {7'd0,(kernel[3][1] ~^ image[15][13])} + {7'd0,(kernel[3][2] ~^ image[15][14])} + {7'd0,(kernel[3][3] ~^ image[15][15])} + {7'd0,(kernel[3][4] ~^ image[15][16])} + {7'd0,(kernel[4][0] ~^ image[16][12])} + {7'd0,(kernel[4][1] ~^ image[16][13])} + {7'd0,(kernel[4][2] ~^ image[16][14])} + {7'd0,(kernel[4][3] ~^ image[16][15])} + {7'd0,(kernel[4][4] ~^ image[16][16])};
assign out_fmap[12][13][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[12][13])} + {7'd0,(kernel[0][1] ~^ image[12][14])} + {7'd0,(kernel[0][2] ~^ image[12][15])} + {7'd0,(kernel[0][3] ~^ image[12][16])} + {7'd0,(kernel[0][4] ~^ image[12][17])} + {7'd0,(kernel[1][0] ~^ image[13][13])} + {7'd0,(kernel[1][1] ~^ image[13][14])} + {7'd0,(kernel[1][2] ~^ image[13][15])} + {7'd0,(kernel[1][3] ~^ image[13][16])} + {7'd0,(kernel[1][4] ~^ image[13][17])} + {7'd0,(kernel[2][0] ~^ image[14][13])} + {7'd0,(kernel[2][1] ~^ image[14][14])} + {7'd0,(kernel[2][2] ~^ image[14][15])} + {7'd0,(kernel[2][3] ~^ image[14][16])} + {7'd0,(kernel[2][4] ~^ image[14][17])} + {7'd0,(kernel[3][0] ~^ image[15][13])} + {7'd0,(kernel[3][1] ~^ image[15][14])} + {7'd0,(kernel[3][2] ~^ image[15][15])} + {7'd0,(kernel[3][3] ~^ image[15][16])} + {7'd0,(kernel[3][4] ~^ image[15][17])} + {7'd0,(kernel[4][0] ~^ image[16][13])} + {7'd0,(kernel[4][1] ~^ image[16][14])} + {7'd0,(kernel[4][2] ~^ image[16][15])} + {7'd0,(kernel[4][3] ~^ image[16][16])} + {7'd0,(kernel[4][4] ~^ image[16][17])};
assign out_fmap[12][14][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[12][14])} + {7'd0,(kernel[0][1] ~^ image[12][15])} + {7'd0,(kernel[0][2] ~^ image[12][16])} + {7'd0,(kernel[0][3] ~^ image[12][17])} + {7'd0,(kernel[0][4] ~^ image[12][18])} + {7'd0,(kernel[1][0] ~^ image[13][14])} + {7'd0,(kernel[1][1] ~^ image[13][15])} + {7'd0,(kernel[1][2] ~^ image[13][16])} + {7'd0,(kernel[1][3] ~^ image[13][17])} + {7'd0,(kernel[1][4] ~^ image[13][18])} + {7'd0,(kernel[2][0] ~^ image[14][14])} + {7'd0,(kernel[2][1] ~^ image[14][15])} + {7'd0,(kernel[2][2] ~^ image[14][16])} + {7'd0,(kernel[2][3] ~^ image[14][17])} + {7'd0,(kernel[2][4] ~^ image[14][18])} + {7'd0,(kernel[3][0] ~^ image[15][14])} + {7'd0,(kernel[3][1] ~^ image[15][15])} + {7'd0,(kernel[3][2] ~^ image[15][16])} + {7'd0,(kernel[3][3] ~^ image[15][17])} + {7'd0,(kernel[3][4] ~^ image[15][18])} + {7'd0,(kernel[4][0] ~^ image[16][14])} + {7'd0,(kernel[4][1] ~^ image[16][15])} + {7'd0,(kernel[4][2] ~^ image[16][16])} + {7'd0,(kernel[4][3] ~^ image[16][17])} + {7'd0,(kernel[4][4] ~^ image[16][18])};
assign out_fmap[12][15][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[12][15])} + {7'd0,(kernel[0][1] ~^ image[12][16])} + {7'd0,(kernel[0][2] ~^ image[12][17])} + {7'd0,(kernel[0][3] ~^ image[12][18])} + {7'd0,(kernel[0][4] ~^ image[12][19])} + {7'd0,(kernel[1][0] ~^ image[13][15])} + {7'd0,(kernel[1][1] ~^ image[13][16])} + {7'd0,(kernel[1][2] ~^ image[13][17])} + {7'd0,(kernel[1][3] ~^ image[13][18])} + {7'd0,(kernel[1][4] ~^ image[13][19])} + {7'd0,(kernel[2][0] ~^ image[14][15])} + {7'd0,(kernel[2][1] ~^ image[14][16])} + {7'd0,(kernel[2][2] ~^ image[14][17])} + {7'd0,(kernel[2][3] ~^ image[14][18])} + {7'd0,(kernel[2][4] ~^ image[14][19])} + {7'd0,(kernel[3][0] ~^ image[15][15])} + {7'd0,(kernel[3][1] ~^ image[15][16])} + {7'd0,(kernel[3][2] ~^ image[15][17])} + {7'd0,(kernel[3][3] ~^ image[15][18])} + {7'd0,(kernel[3][4] ~^ image[15][19])} + {7'd0,(kernel[4][0] ~^ image[16][15])} + {7'd0,(kernel[4][1] ~^ image[16][16])} + {7'd0,(kernel[4][2] ~^ image[16][17])} + {7'd0,(kernel[4][3] ~^ image[16][18])} + {7'd0,(kernel[4][4] ~^ image[16][19])};
assign out_fmap[12][16][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[12][16])} + {7'd0,(kernel[0][1] ~^ image[12][17])} + {7'd0,(kernel[0][2] ~^ image[12][18])} + {7'd0,(kernel[0][3] ~^ image[12][19])} + {7'd0,(kernel[0][4] ~^ image[12][20])} + {7'd0,(kernel[1][0] ~^ image[13][16])} + {7'd0,(kernel[1][1] ~^ image[13][17])} + {7'd0,(kernel[1][2] ~^ image[13][18])} + {7'd0,(kernel[1][3] ~^ image[13][19])} + {7'd0,(kernel[1][4] ~^ image[13][20])} + {7'd0,(kernel[2][0] ~^ image[14][16])} + {7'd0,(kernel[2][1] ~^ image[14][17])} + {7'd0,(kernel[2][2] ~^ image[14][18])} + {7'd0,(kernel[2][3] ~^ image[14][19])} + {7'd0,(kernel[2][4] ~^ image[14][20])} + {7'd0,(kernel[3][0] ~^ image[15][16])} + {7'd0,(kernel[3][1] ~^ image[15][17])} + {7'd0,(kernel[3][2] ~^ image[15][18])} + {7'd0,(kernel[3][3] ~^ image[15][19])} + {7'd0,(kernel[3][4] ~^ image[15][20])} + {7'd0,(kernel[4][0] ~^ image[16][16])} + {7'd0,(kernel[4][1] ~^ image[16][17])} + {7'd0,(kernel[4][2] ~^ image[16][18])} + {7'd0,(kernel[4][3] ~^ image[16][19])} + {7'd0,(kernel[4][4] ~^ image[16][20])};
assign out_fmap[12][17][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[12][17])} + {7'd0,(kernel[0][1] ~^ image[12][18])} + {7'd0,(kernel[0][2] ~^ image[12][19])} + {7'd0,(kernel[0][3] ~^ image[12][20])} + {7'd0,(kernel[0][4] ~^ image[12][21])} + {7'd0,(kernel[1][0] ~^ image[13][17])} + {7'd0,(kernel[1][1] ~^ image[13][18])} + {7'd0,(kernel[1][2] ~^ image[13][19])} + {7'd0,(kernel[1][3] ~^ image[13][20])} + {7'd0,(kernel[1][4] ~^ image[13][21])} + {7'd0,(kernel[2][0] ~^ image[14][17])} + {7'd0,(kernel[2][1] ~^ image[14][18])} + {7'd0,(kernel[2][2] ~^ image[14][19])} + {7'd0,(kernel[2][3] ~^ image[14][20])} + {7'd0,(kernel[2][4] ~^ image[14][21])} + {7'd0,(kernel[3][0] ~^ image[15][17])} + {7'd0,(kernel[3][1] ~^ image[15][18])} + {7'd0,(kernel[3][2] ~^ image[15][19])} + {7'd0,(kernel[3][3] ~^ image[15][20])} + {7'd0,(kernel[3][4] ~^ image[15][21])} + {7'd0,(kernel[4][0] ~^ image[16][17])} + {7'd0,(kernel[4][1] ~^ image[16][18])} + {7'd0,(kernel[4][2] ~^ image[16][19])} + {7'd0,(kernel[4][3] ~^ image[16][20])} + {7'd0,(kernel[4][4] ~^ image[16][21])};
assign out_fmap[12][18][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[12][18])} + {7'd0,(kernel[0][1] ~^ image[12][19])} + {7'd0,(kernel[0][2] ~^ image[12][20])} + {7'd0,(kernel[0][3] ~^ image[12][21])} + {7'd0,(kernel[0][4] ~^ image[12][22])} + {7'd0,(kernel[1][0] ~^ image[13][18])} + {7'd0,(kernel[1][1] ~^ image[13][19])} + {7'd0,(kernel[1][2] ~^ image[13][20])} + {7'd0,(kernel[1][3] ~^ image[13][21])} + {7'd0,(kernel[1][4] ~^ image[13][22])} + {7'd0,(kernel[2][0] ~^ image[14][18])} + {7'd0,(kernel[2][1] ~^ image[14][19])} + {7'd0,(kernel[2][2] ~^ image[14][20])} + {7'd0,(kernel[2][3] ~^ image[14][21])} + {7'd0,(kernel[2][4] ~^ image[14][22])} + {7'd0,(kernel[3][0] ~^ image[15][18])} + {7'd0,(kernel[3][1] ~^ image[15][19])} + {7'd0,(kernel[3][2] ~^ image[15][20])} + {7'd0,(kernel[3][3] ~^ image[15][21])} + {7'd0,(kernel[3][4] ~^ image[15][22])} + {7'd0,(kernel[4][0] ~^ image[16][18])} + {7'd0,(kernel[4][1] ~^ image[16][19])} + {7'd0,(kernel[4][2] ~^ image[16][20])} + {7'd0,(kernel[4][3] ~^ image[16][21])} + {7'd0,(kernel[4][4] ~^ image[16][22])};
assign out_fmap[12][19][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[12][19])} + {7'd0,(kernel[0][1] ~^ image[12][20])} + {7'd0,(kernel[0][2] ~^ image[12][21])} + {7'd0,(kernel[0][3] ~^ image[12][22])} + {7'd0,(kernel[0][4] ~^ image[12][23])} + {7'd0,(kernel[1][0] ~^ image[13][19])} + {7'd0,(kernel[1][1] ~^ image[13][20])} + {7'd0,(kernel[1][2] ~^ image[13][21])} + {7'd0,(kernel[1][3] ~^ image[13][22])} + {7'd0,(kernel[1][4] ~^ image[13][23])} + {7'd0,(kernel[2][0] ~^ image[14][19])} + {7'd0,(kernel[2][1] ~^ image[14][20])} + {7'd0,(kernel[2][2] ~^ image[14][21])} + {7'd0,(kernel[2][3] ~^ image[14][22])} + {7'd0,(kernel[2][4] ~^ image[14][23])} + {7'd0,(kernel[3][0] ~^ image[15][19])} + {7'd0,(kernel[3][1] ~^ image[15][20])} + {7'd0,(kernel[3][2] ~^ image[15][21])} + {7'd0,(kernel[3][3] ~^ image[15][22])} + {7'd0,(kernel[3][4] ~^ image[15][23])} + {7'd0,(kernel[4][0] ~^ image[16][19])} + {7'd0,(kernel[4][1] ~^ image[16][20])} + {7'd0,(kernel[4][2] ~^ image[16][21])} + {7'd0,(kernel[4][3] ~^ image[16][22])} + {7'd0,(kernel[4][4] ~^ image[16][23])};
assign out_fmap[12][20][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[12][20])} + {7'd0,(kernel[0][1] ~^ image[12][21])} + {7'd0,(kernel[0][2] ~^ image[12][22])} + {7'd0,(kernel[0][3] ~^ image[12][23])} + {7'd0,(kernel[0][4] ~^ image[12][24])} + {7'd0,(kernel[1][0] ~^ image[13][20])} + {7'd0,(kernel[1][1] ~^ image[13][21])} + {7'd0,(kernel[1][2] ~^ image[13][22])} + {7'd0,(kernel[1][3] ~^ image[13][23])} + {7'd0,(kernel[1][4] ~^ image[13][24])} + {7'd0,(kernel[2][0] ~^ image[14][20])} + {7'd0,(kernel[2][1] ~^ image[14][21])} + {7'd0,(kernel[2][2] ~^ image[14][22])} + {7'd0,(kernel[2][3] ~^ image[14][23])} + {7'd0,(kernel[2][4] ~^ image[14][24])} + {7'd0,(kernel[3][0] ~^ image[15][20])} + {7'd0,(kernel[3][1] ~^ image[15][21])} + {7'd0,(kernel[3][2] ~^ image[15][22])} + {7'd0,(kernel[3][3] ~^ image[15][23])} + {7'd0,(kernel[3][4] ~^ image[15][24])} + {7'd0,(kernel[4][0] ~^ image[16][20])} + {7'd0,(kernel[4][1] ~^ image[16][21])} + {7'd0,(kernel[4][2] ~^ image[16][22])} + {7'd0,(kernel[4][3] ~^ image[16][23])} + {7'd0,(kernel[4][4] ~^ image[16][24])};
assign out_fmap[12][21][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[12][21])} + {7'd0,(kernel[0][1] ~^ image[12][22])} + {7'd0,(kernel[0][2] ~^ image[12][23])} + {7'd0,(kernel[0][3] ~^ image[12][24])} + {7'd0,(kernel[0][4] ~^ image[12][25])} + {7'd0,(kernel[1][0] ~^ image[13][21])} + {7'd0,(kernel[1][1] ~^ image[13][22])} + {7'd0,(kernel[1][2] ~^ image[13][23])} + {7'd0,(kernel[1][3] ~^ image[13][24])} + {7'd0,(kernel[1][4] ~^ image[13][25])} + {7'd0,(kernel[2][0] ~^ image[14][21])} + {7'd0,(kernel[2][1] ~^ image[14][22])} + {7'd0,(kernel[2][2] ~^ image[14][23])} + {7'd0,(kernel[2][3] ~^ image[14][24])} + {7'd0,(kernel[2][4] ~^ image[14][25])} + {7'd0,(kernel[3][0] ~^ image[15][21])} + {7'd0,(kernel[3][1] ~^ image[15][22])} + {7'd0,(kernel[3][2] ~^ image[15][23])} + {7'd0,(kernel[3][3] ~^ image[15][24])} + {7'd0,(kernel[3][4] ~^ image[15][25])} + {7'd0,(kernel[4][0] ~^ image[16][21])} + {7'd0,(kernel[4][1] ~^ image[16][22])} + {7'd0,(kernel[4][2] ~^ image[16][23])} + {7'd0,(kernel[4][3] ~^ image[16][24])} + {7'd0,(kernel[4][4] ~^ image[16][25])};
assign out_fmap[12][22][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[12][22])} + {7'd0,(kernel[0][1] ~^ image[12][23])} + {7'd0,(kernel[0][2] ~^ image[12][24])} + {7'd0,(kernel[0][3] ~^ image[12][25])} + {7'd0,(kernel[0][4] ~^ image[12][26])} + {7'd0,(kernel[1][0] ~^ image[13][22])} + {7'd0,(kernel[1][1] ~^ image[13][23])} + {7'd0,(kernel[1][2] ~^ image[13][24])} + {7'd0,(kernel[1][3] ~^ image[13][25])} + {7'd0,(kernel[1][4] ~^ image[13][26])} + {7'd0,(kernel[2][0] ~^ image[14][22])} + {7'd0,(kernel[2][1] ~^ image[14][23])} + {7'd0,(kernel[2][2] ~^ image[14][24])} + {7'd0,(kernel[2][3] ~^ image[14][25])} + {7'd0,(kernel[2][4] ~^ image[14][26])} + {7'd0,(kernel[3][0] ~^ image[15][22])} + {7'd0,(kernel[3][1] ~^ image[15][23])} + {7'd0,(kernel[3][2] ~^ image[15][24])} + {7'd0,(kernel[3][3] ~^ image[15][25])} + {7'd0,(kernel[3][4] ~^ image[15][26])} + {7'd0,(kernel[4][0] ~^ image[16][22])} + {7'd0,(kernel[4][1] ~^ image[16][23])} + {7'd0,(kernel[4][2] ~^ image[16][24])} + {7'd0,(kernel[4][3] ~^ image[16][25])} + {7'd0,(kernel[4][4] ~^ image[16][26])};
assign out_fmap[12][23][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[12][23])} + {7'd0,(kernel[0][1] ~^ image[12][24])} + {7'd0,(kernel[0][2] ~^ image[12][25])} + {7'd0,(kernel[0][3] ~^ image[12][26])} + {7'd0,(kernel[0][4] ~^ image[12][27])} + {7'd0,(kernel[1][0] ~^ image[13][23])} + {7'd0,(kernel[1][1] ~^ image[13][24])} + {7'd0,(kernel[1][2] ~^ image[13][25])} + {7'd0,(kernel[1][3] ~^ image[13][26])} + {7'd0,(kernel[1][4] ~^ image[13][27])} + {7'd0,(kernel[2][0] ~^ image[14][23])} + {7'd0,(kernel[2][1] ~^ image[14][24])} + {7'd0,(kernel[2][2] ~^ image[14][25])} + {7'd0,(kernel[2][3] ~^ image[14][26])} + {7'd0,(kernel[2][4] ~^ image[14][27])} + {7'd0,(kernel[3][0] ~^ image[15][23])} + {7'd0,(kernel[3][1] ~^ image[15][24])} + {7'd0,(kernel[3][2] ~^ image[15][25])} + {7'd0,(kernel[3][3] ~^ image[15][26])} + {7'd0,(kernel[3][4] ~^ image[15][27])} + {7'd0,(kernel[4][0] ~^ image[16][23])} + {7'd0,(kernel[4][1] ~^ image[16][24])} + {7'd0,(kernel[4][2] ~^ image[16][25])} + {7'd0,(kernel[4][3] ~^ image[16][26])} + {7'd0,(kernel[4][4] ~^ image[16][27])};
assign out_fmap[13][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[13][0])} + {7'd0,(kernel[0][1] ~^ image[13][1])} + {7'd0,(kernel[0][2] ~^ image[13][2])} + {7'd0,(kernel[0][3] ~^ image[13][3])} + {7'd0,(kernel[0][4] ~^ image[13][4])} + {7'd0,(kernel[1][0] ~^ image[14][0])} + {7'd0,(kernel[1][1] ~^ image[14][1])} + {7'd0,(kernel[1][2] ~^ image[14][2])} + {7'd0,(kernel[1][3] ~^ image[14][3])} + {7'd0,(kernel[1][4] ~^ image[14][4])} + {7'd0,(kernel[2][0] ~^ image[15][0])} + {7'd0,(kernel[2][1] ~^ image[15][1])} + {7'd0,(kernel[2][2] ~^ image[15][2])} + {7'd0,(kernel[2][3] ~^ image[15][3])} + {7'd0,(kernel[2][4] ~^ image[15][4])} + {7'd0,(kernel[3][0] ~^ image[16][0])} + {7'd0,(kernel[3][1] ~^ image[16][1])} + {7'd0,(kernel[3][2] ~^ image[16][2])} + {7'd0,(kernel[3][3] ~^ image[16][3])} + {7'd0,(kernel[3][4] ~^ image[16][4])} + {7'd0,(kernel[4][0] ~^ image[17][0])} + {7'd0,(kernel[4][1] ~^ image[17][1])} + {7'd0,(kernel[4][2] ~^ image[17][2])} + {7'd0,(kernel[4][3] ~^ image[17][3])} + {7'd0,(kernel[4][4] ~^ image[17][4])};
assign out_fmap[13][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[13][1])} + {7'd0,(kernel[0][1] ~^ image[13][2])} + {7'd0,(kernel[0][2] ~^ image[13][3])} + {7'd0,(kernel[0][3] ~^ image[13][4])} + {7'd0,(kernel[0][4] ~^ image[13][5])} + {7'd0,(kernel[1][0] ~^ image[14][1])} + {7'd0,(kernel[1][1] ~^ image[14][2])} + {7'd0,(kernel[1][2] ~^ image[14][3])} + {7'd0,(kernel[1][3] ~^ image[14][4])} + {7'd0,(kernel[1][4] ~^ image[14][5])} + {7'd0,(kernel[2][0] ~^ image[15][1])} + {7'd0,(kernel[2][1] ~^ image[15][2])} + {7'd0,(kernel[2][2] ~^ image[15][3])} + {7'd0,(kernel[2][3] ~^ image[15][4])} + {7'd0,(kernel[2][4] ~^ image[15][5])} + {7'd0,(kernel[3][0] ~^ image[16][1])} + {7'd0,(kernel[3][1] ~^ image[16][2])} + {7'd0,(kernel[3][2] ~^ image[16][3])} + {7'd0,(kernel[3][3] ~^ image[16][4])} + {7'd0,(kernel[3][4] ~^ image[16][5])} + {7'd0,(kernel[4][0] ~^ image[17][1])} + {7'd0,(kernel[4][1] ~^ image[17][2])} + {7'd0,(kernel[4][2] ~^ image[17][3])} + {7'd0,(kernel[4][3] ~^ image[17][4])} + {7'd0,(kernel[4][4] ~^ image[17][5])};
assign out_fmap[13][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[13][2])} + {7'd0,(kernel[0][1] ~^ image[13][3])} + {7'd0,(kernel[0][2] ~^ image[13][4])} + {7'd0,(kernel[0][3] ~^ image[13][5])} + {7'd0,(kernel[0][4] ~^ image[13][6])} + {7'd0,(kernel[1][0] ~^ image[14][2])} + {7'd0,(kernel[1][1] ~^ image[14][3])} + {7'd0,(kernel[1][2] ~^ image[14][4])} + {7'd0,(kernel[1][3] ~^ image[14][5])} + {7'd0,(kernel[1][4] ~^ image[14][6])} + {7'd0,(kernel[2][0] ~^ image[15][2])} + {7'd0,(kernel[2][1] ~^ image[15][3])} + {7'd0,(kernel[2][2] ~^ image[15][4])} + {7'd0,(kernel[2][3] ~^ image[15][5])} + {7'd0,(kernel[2][4] ~^ image[15][6])} + {7'd0,(kernel[3][0] ~^ image[16][2])} + {7'd0,(kernel[3][1] ~^ image[16][3])} + {7'd0,(kernel[3][2] ~^ image[16][4])} + {7'd0,(kernel[3][3] ~^ image[16][5])} + {7'd0,(kernel[3][4] ~^ image[16][6])} + {7'd0,(kernel[4][0] ~^ image[17][2])} + {7'd0,(kernel[4][1] ~^ image[17][3])} + {7'd0,(kernel[4][2] ~^ image[17][4])} + {7'd0,(kernel[4][3] ~^ image[17][5])} + {7'd0,(kernel[4][4] ~^ image[17][6])};
assign out_fmap[13][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[13][3])} + {7'd0,(kernel[0][1] ~^ image[13][4])} + {7'd0,(kernel[0][2] ~^ image[13][5])} + {7'd0,(kernel[0][3] ~^ image[13][6])} + {7'd0,(kernel[0][4] ~^ image[13][7])} + {7'd0,(kernel[1][0] ~^ image[14][3])} + {7'd0,(kernel[1][1] ~^ image[14][4])} + {7'd0,(kernel[1][2] ~^ image[14][5])} + {7'd0,(kernel[1][3] ~^ image[14][6])} + {7'd0,(kernel[1][4] ~^ image[14][7])} + {7'd0,(kernel[2][0] ~^ image[15][3])} + {7'd0,(kernel[2][1] ~^ image[15][4])} + {7'd0,(kernel[2][2] ~^ image[15][5])} + {7'd0,(kernel[2][3] ~^ image[15][6])} + {7'd0,(kernel[2][4] ~^ image[15][7])} + {7'd0,(kernel[3][0] ~^ image[16][3])} + {7'd0,(kernel[3][1] ~^ image[16][4])} + {7'd0,(kernel[3][2] ~^ image[16][5])} + {7'd0,(kernel[3][3] ~^ image[16][6])} + {7'd0,(kernel[3][4] ~^ image[16][7])} + {7'd0,(kernel[4][0] ~^ image[17][3])} + {7'd0,(kernel[4][1] ~^ image[17][4])} + {7'd0,(kernel[4][2] ~^ image[17][5])} + {7'd0,(kernel[4][3] ~^ image[17][6])} + {7'd0,(kernel[4][4] ~^ image[17][7])};
assign out_fmap[13][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[13][4])} + {7'd0,(kernel[0][1] ~^ image[13][5])} + {7'd0,(kernel[0][2] ~^ image[13][6])} + {7'd0,(kernel[0][3] ~^ image[13][7])} + {7'd0,(kernel[0][4] ~^ image[13][8])} + {7'd0,(kernel[1][0] ~^ image[14][4])} + {7'd0,(kernel[1][1] ~^ image[14][5])} + {7'd0,(kernel[1][2] ~^ image[14][6])} + {7'd0,(kernel[1][3] ~^ image[14][7])} + {7'd0,(kernel[1][4] ~^ image[14][8])} + {7'd0,(kernel[2][0] ~^ image[15][4])} + {7'd0,(kernel[2][1] ~^ image[15][5])} + {7'd0,(kernel[2][2] ~^ image[15][6])} + {7'd0,(kernel[2][3] ~^ image[15][7])} + {7'd0,(kernel[2][4] ~^ image[15][8])} + {7'd0,(kernel[3][0] ~^ image[16][4])} + {7'd0,(kernel[3][1] ~^ image[16][5])} + {7'd0,(kernel[3][2] ~^ image[16][6])} + {7'd0,(kernel[3][3] ~^ image[16][7])} + {7'd0,(kernel[3][4] ~^ image[16][8])} + {7'd0,(kernel[4][0] ~^ image[17][4])} + {7'd0,(kernel[4][1] ~^ image[17][5])} + {7'd0,(kernel[4][2] ~^ image[17][6])} + {7'd0,(kernel[4][3] ~^ image[17][7])} + {7'd0,(kernel[4][4] ~^ image[17][8])};
assign out_fmap[13][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[13][5])} + {7'd0,(kernel[0][1] ~^ image[13][6])} + {7'd0,(kernel[0][2] ~^ image[13][7])} + {7'd0,(kernel[0][3] ~^ image[13][8])} + {7'd0,(kernel[0][4] ~^ image[13][9])} + {7'd0,(kernel[1][0] ~^ image[14][5])} + {7'd0,(kernel[1][1] ~^ image[14][6])} + {7'd0,(kernel[1][2] ~^ image[14][7])} + {7'd0,(kernel[1][3] ~^ image[14][8])} + {7'd0,(kernel[1][4] ~^ image[14][9])} + {7'd0,(kernel[2][0] ~^ image[15][5])} + {7'd0,(kernel[2][1] ~^ image[15][6])} + {7'd0,(kernel[2][2] ~^ image[15][7])} + {7'd0,(kernel[2][3] ~^ image[15][8])} + {7'd0,(kernel[2][4] ~^ image[15][9])} + {7'd0,(kernel[3][0] ~^ image[16][5])} + {7'd0,(kernel[3][1] ~^ image[16][6])} + {7'd0,(kernel[3][2] ~^ image[16][7])} + {7'd0,(kernel[3][3] ~^ image[16][8])} + {7'd0,(kernel[3][4] ~^ image[16][9])} + {7'd0,(kernel[4][0] ~^ image[17][5])} + {7'd0,(kernel[4][1] ~^ image[17][6])} + {7'd0,(kernel[4][2] ~^ image[17][7])} + {7'd0,(kernel[4][3] ~^ image[17][8])} + {7'd0,(kernel[4][4] ~^ image[17][9])};
assign out_fmap[13][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[13][6])} + {7'd0,(kernel[0][1] ~^ image[13][7])} + {7'd0,(kernel[0][2] ~^ image[13][8])} + {7'd0,(kernel[0][3] ~^ image[13][9])} + {7'd0,(kernel[0][4] ~^ image[13][10])} + {7'd0,(kernel[1][0] ~^ image[14][6])} + {7'd0,(kernel[1][1] ~^ image[14][7])} + {7'd0,(kernel[1][2] ~^ image[14][8])} + {7'd0,(kernel[1][3] ~^ image[14][9])} + {7'd0,(kernel[1][4] ~^ image[14][10])} + {7'd0,(kernel[2][0] ~^ image[15][6])} + {7'd0,(kernel[2][1] ~^ image[15][7])} + {7'd0,(kernel[2][2] ~^ image[15][8])} + {7'd0,(kernel[2][3] ~^ image[15][9])} + {7'd0,(kernel[2][4] ~^ image[15][10])} + {7'd0,(kernel[3][0] ~^ image[16][6])} + {7'd0,(kernel[3][1] ~^ image[16][7])} + {7'd0,(kernel[3][2] ~^ image[16][8])} + {7'd0,(kernel[3][3] ~^ image[16][9])} + {7'd0,(kernel[3][4] ~^ image[16][10])} + {7'd0,(kernel[4][0] ~^ image[17][6])} + {7'd0,(kernel[4][1] ~^ image[17][7])} + {7'd0,(kernel[4][2] ~^ image[17][8])} + {7'd0,(kernel[4][3] ~^ image[17][9])} + {7'd0,(kernel[4][4] ~^ image[17][10])};
assign out_fmap[13][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[13][7])} + {7'd0,(kernel[0][1] ~^ image[13][8])} + {7'd0,(kernel[0][2] ~^ image[13][9])} + {7'd0,(kernel[0][3] ~^ image[13][10])} + {7'd0,(kernel[0][4] ~^ image[13][11])} + {7'd0,(kernel[1][0] ~^ image[14][7])} + {7'd0,(kernel[1][1] ~^ image[14][8])} + {7'd0,(kernel[1][2] ~^ image[14][9])} + {7'd0,(kernel[1][3] ~^ image[14][10])} + {7'd0,(kernel[1][4] ~^ image[14][11])} + {7'd0,(kernel[2][0] ~^ image[15][7])} + {7'd0,(kernel[2][1] ~^ image[15][8])} + {7'd0,(kernel[2][2] ~^ image[15][9])} + {7'd0,(kernel[2][3] ~^ image[15][10])} + {7'd0,(kernel[2][4] ~^ image[15][11])} + {7'd0,(kernel[3][0] ~^ image[16][7])} + {7'd0,(kernel[3][1] ~^ image[16][8])} + {7'd0,(kernel[3][2] ~^ image[16][9])} + {7'd0,(kernel[3][3] ~^ image[16][10])} + {7'd0,(kernel[3][4] ~^ image[16][11])} + {7'd0,(kernel[4][0] ~^ image[17][7])} + {7'd0,(kernel[4][1] ~^ image[17][8])} + {7'd0,(kernel[4][2] ~^ image[17][9])} + {7'd0,(kernel[4][3] ~^ image[17][10])} + {7'd0,(kernel[4][4] ~^ image[17][11])};
assign out_fmap[13][8][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[13][8])} + {7'd0,(kernel[0][1] ~^ image[13][9])} + {7'd0,(kernel[0][2] ~^ image[13][10])} + {7'd0,(kernel[0][3] ~^ image[13][11])} + {7'd0,(kernel[0][4] ~^ image[13][12])} + {7'd0,(kernel[1][0] ~^ image[14][8])} + {7'd0,(kernel[1][1] ~^ image[14][9])} + {7'd0,(kernel[1][2] ~^ image[14][10])} + {7'd0,(kernel[1][3] ~^ image[14][11])} + {7'd0,(kernel[1][4] ~^ image[14][12])} + {7'd0,(kernel[2][0] ~^ image[15][8])} + {7'd0,(kernel[2][1] ~^ image[15][9])} + {7'd0,(kernel[2][2] ~^ image[15][10])} + {7'd0,(kernel[2][3] ~^ image[15][11])} + {7'd0,(kernel[2][4] ~^ image[15][12])} + {7'd0,(kernel[3][0] ~^ image[16][8])} + {7'd0,(kernel[3][1] ~^ image[16][9])} + {7'd0,(kernel[3][2] ~^ image[16][10])} + {7'd0,(kernel[3][3] ~^ image[16][11])} + {7'd0,(kernel[3][4] ~^ image[16][12])} + {7'd0,(kernel[4][0] ~^ image[17][8])} + {7'd0,(kernel[4][1] ~^ image[17][9])} + {7'd0,(kernel[4][2] ~^ image[17][10])} + {7'd0,(kernel[4][3] ~^ image[17][11])} + {7'd0,(kernel[4][4] ~^ image[17][12])};
assign out_fmap[13][9][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[13][9])} + {7'd0,(kernel[0][1] ~^ image[13][10])} + {7'd0,(kernel[0][2] ~^ image[13][11])} + {7'd0,(kernel[0][3] ~^ image[13][12])} + {7'd0,(kernel[0][4] ~^ image[13][13])} + {7'd0,(kernel[1][0] ~^ image[14][9])} + {7'd0,(kernel[1][1] ~^ image[14][10])} + {7'd0,(kernel[1][2] ~^ image[14][11])} + {7'd0,(kernel[1][3] ~^ image[14][12])} + {7'd0,(kernel[1][4] ~^ image[14][13])} + {7'd0,(kernel[2][0] ~^ image[15][9])} + {7'd0,(kernel[2][1] ~^ image[15][10])} + {7'd0,(kernel[2][2] ~^ image[15][11])} + {7'd0,(kernel[2][3] ~^ image[15][12])} + {7'd0,(kernel[2][4] ~^ image[15][13])} + {7'd0,(kernel[3][0] ~^ image[16][9])} + {7'd0,(kernel[3][1] ~^ image[16][10])} + {7'd0,(kernel[3][2] ~^ image[16][11])} + {7'd0,(kernel[3][3] ~^ image[16][12])} + {7'd0,(kernel[3][4] ~^ image[16][13])} + {7'd0,(kernel[4][0] ~^ image[17][9])} + {7'd0,(kernel[4][1] ~^ image[17][10])} + {7'd0,(kernel[4][2] ~^ image[17][11])} + {7'd0,(kernel[4][3] ~^ image[17][12])} + {7'd0,(kernel[4][4] ~^ image[17][13])};
assign out_fmap[13][10][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[13][10])} + {7'd0,(kernel[0][1] ~^ image[13][11])} + {7'd0,(kernel[0][2] ~^ image[13][12])} + {7'd0,(kernel[0][3] ~^ image[13][13])} + {7'd0,(kernel[0][4] ~^ image[13][14])} + {7'd0,(kernel[1][0] ~^ image[14][10])} + {7'd0,(kernel[1][1] ~^ image[14][11])} + {7'd0,(kernel[1][2] ~^ image[14][12])} + {7'd0,(kernel[1][3] ~^ image[14][13])} + {7'd0,(kernel[1][4] ~^ image[14][14])} + {7'd0,(kernel[2][0] ~^ image[15][10])} + {7'd0,(kernel[2][1] ~^ image[15][11])} + {7'd0,(kernel[2][2] ~^ image[15][12])} + {7'd0,(kernel[2][3] ~^ image[15][13])} + {7'd0,(kernel[2][4] ~^ image[15][14])} + {7'd0,(kernel[3][0] ~^ image[16][10])} + {7'd0,(kernel[3][1] ~^ image[16][11])} + {7'd0,(kernel[3][2] ~^ image[16][12])} + {7'd0,(kernel[3][3] ~^ image[16][13])} + {7'd0,(kernel[3][4] ~^ image[16][14])} + {7'd0,(kernel[4][0] ~^ image[17][10])} + {7'd0,(kernel[4][1] ~^ image[17][11])} + {7'd0,(kernel[4][2] ~^ image[17][12])} + {7'd0,(kernel[4][3] ~^ image[17][13])} + {7'd0,(kernel[4][4] ~^ image[17][14])};
assign out_fmap[13][11][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[13][11])} + {7'd0,(kernel[0][1] ~^ image[13][12])} + {7'd0,(kernel[0][2] ~^ image[13][13])} + {7'd0,(kernel[0][3] ~^ image[13][14])} + {7'd0,(kernel[0][4] ~^ image[13][15])} + {7'd0,(kernel[1][0] ~^ image[14][11])} + {7'd0,(kernel[1][1] ~^ image[14][12])} + {7'd0,(kernel[1][2] ~^ image[14][13])} + {7'd0,(kernel[1][3] ~^ image[14][14])} + {7'd0,(kernel[1][4] ~^ image[14][15])} + {7'd0,(kernel[2][0] ~^ image[15][11])} + {7'd0,(kernel[2][1] ~^ image[15][12])} + {7'd0,(kernel[2][2] ~^ image[15][13])} + {7'd0,(kernel[2][3] ~^ image[15][14])} + {7'd0,(kernel[2][4] ~^ image[15][15])} + {7'd0,(kernel[3][0] ~^ image[16][11])} + {7'd0,(kernel[3][1] ~^ image[16][12])} + {7'd0,(kernel[3][2] ~^ image[16][13])} + {7'd0,(kernel[3][3] ~^ image[16][14])} + {7'd0,(kernel[3][4] ~^ image[16][15])} + {7'd0,(kernel[4][0] ~^ image[17][11])} + {7'd0,(kernel[4][1] ~^ image[17][12])} + {7'd0,(kernel[4][2] ~^ image[17][13])} + {7'd0,(kernel[4][3] ~^ image[17][14])} + {7'd0,(kernel[4][4] ~^ image[17][15])};
assign out_fmap[13][12][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[13][12])} + {7'd0,(kernel[0][1] ~^ image[13][13])} + {7'd0,(kernel[0][2] ~^ image[13][14])} + {7'd0,(kernel[0][3] ~^ image[13][15])} + {7'd0,(kernel[0][4] ~^ image[13][16])} + {7'd0,(kernel[1][0] ~^ image[14][12])} + {7'd0,(kernel[1][1] ~^ image[14][13])} + {7'd0,(kernel[1][2] ~^ image[14][14])} + {7'd0,(kernel[1][3] ~^ image[14][15])} + {7'd0,(kernel[1][4] ~^ image[14][16])} + {7'd0,(kernel[2][0] ~^ image[15][12])} + {7'd0,(kernel[2][1] ~^ image[15][13])} + {7'd0,(kernel[2][2] ~^ image[15][14])} + {7'd0,(kernel[2][3] ~^ image[15][15])} + {7'd0,(kernel[2][4] ~^ image[15][16])} + {7'd0,(kernel[3][0] ~^ image[16][12])} + {7'd0,(kernel[3][1] ~^ image[16][13])} + {7'd0,(kernel[3][2] ~^ image[16][14])} + {7'd0,(kernel[3][3] ~^ image[16][15])} + {7'd0,(kernel[3][4] ~^ image[16][16])} + {7'd0,(kernel[4][0] ~^ image[17][12])} + {7'd0,(kernel[4][1] ~^ image[17][13])} + {7'd0,(kernel[4][2] ~^ image[17][14])} + {7'd0,(kernel[4][3] ~^ image[17][15])} + {7'd0,(kernel[4][4] ~^ image[17][16])};
assign out_fmap[13][13][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[13][13])} + {7'd0,(kernel[0][1] ~^ image[13][14])} + {7'd0,(kernel[0][2] ~^ image[13][15])} + {7'd0,(kernel[0][3] ~^ image[13][16])} + {7'd0,(kernel[0][4] ~^ image[13][17])} + {7'd0,(kernel[1][0] ~^ image[14][13])} + {7'd0,(kernel[1][1] ~^ image[14][14])} + {7'd0,(kernel[1][2] ~^ image[14][15])} + {7'd0,(kernel[1][3] ~^ image[14][16])} + {7'd0,(kernel[1][4] ~^ image[14][17])} + {7'd0,(kernel[2][0] ~^ image[15][13])} + {7'd0,(kernel[2][1] ~^ image[15][14])} + {7'd0,(kernel[2][2] ~^ image[15][15])} + {7'd0,(kernel[2][3] ~^ image[15][16])} + {7'd0,(kernel[2][4] ~^ image[15][17])} + {7'd0,(kernel[3][0] ~^ image[16][13])} + {7'd0,(kernel[3][1] ~^ image[16][14])} + {7'd0,(kernel[3][2] ~^ image[16][15])} + {7'd0,(kernel[3][3] ~^ image[16][16])} + {7'd0,(kernel[3][4] ~^ image[16][17])} + {7'd0,(kernel[4][0] ~^ image[17][13])} + {7'd0,(kernel[4][1] ~^ image[17][14])} + {7'd0,(kernel[4][2] ~^ image[17][15])} + {7'd0,(kernel[4][3] ~^ image[17][16])} + {7'd0,(kernel[4][4] ~^ image[17][17])};
assign out_fmap[13][14][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[13][14])} + {7'd0,(kernel[0][1] ~^ image[13][15])} + {7'd0,(kernel[0][2] ~^ image[13][16])} + {7'd0,(kernel[0][3] ~^ image[13][17])} + {7'd0,(kernel[0][4] ~^ image[13][18])} + {7'd0,(kernel[1][0] ~^ image[14][14])} + {7'd0,(kernel[1][1] ~^ image[14][15])} + {7'd0,(kernel[1][2] ~^ image[14][16])} + {7'd0,(kernel[1][3] ~^ image[14][17])} + {7'd0,(kernel[1][4] ~^ image[14][18])} + {7'd0,(kernel[2][0] ~^ image[15][14])} + {7'd0,(kernel[2][1] ~^ image[15][15])} + {7'd0,(kernel[2][2] ~^ image[15][16])} + {7'd0,(kernel[2][3] ~^ image[15][17])} + {7'd0,(kernel[2][4] ~^ image[15][18])} + {7'd0,(kernel[3][0] ~^ image[16][14])} + {7'd0,(kernel[3][1] ~^ image[16][15])} + {7'd0,(kernel[3][2] ~^ image[16][16])} + {7'd0,(kernel[3][3] ~^ image[16][17])} + {7'd0,(kernel[3][4] ~^ image[16][18])} + {7'd0,(kernel[4][0] ~^ image[17][14])} + {7'd0,(kernel[4][1] ~^ image[17][15])} + {7'd0,(kernel[4][2] ~^ image[17][16])} + {7'd0,(kernel[4][3] ~^ image[17][17])} + {7'd0,(kernel[4][4] ~^ image[17][18])};
assign out_fmap[13][15][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[13][15])} + {7'd0,(kernel[0][1] ~^ image[13][16])} + {7'd0,(kernel[0][2] ~^ image[13][17])} + {7'd0,(kernel[0][3] ~^ image[13][18])} + {7'd0,(kernel[0][4] ~^ image[13][19])} + {7'd0,(kernel[1][0] ~^ image[14][15])} + {7'd0,(kernel[1][1] ~^ image[14][16])} + {7'd0,(kernel[1][2] ~^ image[14][17])} + {7'd0,(kernel[1][3] ~^ image[14][18])} + {7'd0,(kernel[1][4] ~^ image[14][19])} + {7'd0,(kernel[2][0] ~^ image[15][15])} + {7'd0,(kernel[2][1] ~^ image[15][16])} + {7'd0,(kernel[2][2] ~^ image[15][17])} + {7'd0,(kernel[2][3] ~^ image[15][18])} + {7'd0,(kernel[2][4] ~^ image[15][19])} + {7'd0,(kernel[3][0] ~^ image[16][15])} + {7'd0,(kernel[3][1] ~^ image[16][16])} + {7'd0,(kernel[3][2] ~^ image[16][17])} + {7'd0,(kernel[3][3] ~^ image[16][18])} + {7'd0,(kernel[3][4] ~^ image[16][19])} + {7'd0,(kernel[4][0] ~^ image[17][15])} + {7'd0,(kernel[4][1] ~^ image[17][16])} + {7'd0,(kernel[4][2] ~^ image[17][17])} + {7'd0,(kernel[4][3] ~^ image[17][18])} + {7'd0,(kernel[4][4] ~^ image[17][19])};
assign out_fmap[13][16][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[13][16])} + {7'd0,(kernel[0][1] ~^ image[13][17])} + {7'd0,(kernel[0][2] ~^ image[13][18])} + {7'd0,(kernel[0][3] ~^ image[13][19])} + {7'd0,(kernel[0][4] ~^ image[13][20])} + {7'd0,(kernel[1][0] ~^ image[14][16])} + {7'd0,(kernel[1][1] ~^ image[14][17])} + {7'd0,(kernel[1][2] ~^ image[14][18])} + {7'd0,(kernel[1][3] ~^ image[14][19])} + {7'd0,(kernel[1][4] ~^ image[14][20])} + {7'd0,(kernel[2][0] ~^ image[15][16])} + {7'd0,(kernel[2][1] ~^ image[15][17])} + {7'd0,(kernel[2][2] ~^ image[15][18])} + {7'd0,(kernel[2][3] ~^ image[15][19])} + {7'd0,(kernel[2][4] ~^ image[15][20])} + {7'd0,(kernel[3][0] ~^ image[16][16])} + {7'd0,(kernel[3][1] ~^ image[16][17])} + {7'd0,(kernel[3][2] ~^ image[16][18])} + {7'd0,(kernel[3][3] ~^ image[16][19])} + {7'd0,(kernel[3][4] ~^ image[16][20])} + {7'd0,(kernel[4][0] ~^ image[17][16])} + {7'd0,(kernel[4][1] ~^ image[17][17])} + {7'd0,(kernel[4][2] ~^ image[17][18])} + {7'd0,(kernel[4][3] ~^ image[17][19])} + {7'd0,(kernel[4][4] ~^ image[17][20])};
assign out_fmap[13][17][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[13][17])} + {7'd0,(kernel[0][1] ~^ image[13][18])} + {7'd0,(kernel[0][2] ~^ image[13][19])} + {7'd0,(kernel[0][3] ~^ image[13][20])} + {7'd0,(kernel[0][4] ~^ image[13][21])} + {7'd0,(kernel[1][0] ~^ image[14][17])} + {7'd0,(kernel[1][1] ~^ image[14][18])} + {7'd0,(kernel[1][2] ~^ image[14][19])} + {7'd0,(kernel[1][3] ~^ image[14][20])} + {7'd0,(kernel[1][4] ~^ image[14][21])} + {7'd0,(kernel[2][0] ~^ image[15][17])} + {7'd0,(kernel[2][1] ~^ image[15][18])} + {7'd0,(kernel[2][2] ~^ image[15][19])} + {7'd0,(kernel[2][3] ~^ image[15][20])} + {7'd0,(kernel[2][4] ~^ image[15][21])} + {7'd0,(kernel[3][0] ~^ image[16][17])} + {7'd0,(kernel[3][1] ~^ image[16][18])} + {7'd0,(kernel[3][2] ~^ image[16][19])} + {7'd0,(kernel[3][3] ~^ image[16][20])} + {7'd0,(kernel[3][4] ~^ image[16][21])} + {7'd0,(kernel[4][0] ~^ image[17][17])} + {7'd0,(kernel[4][1] ~^ image[17][18])} + {7'd0,(kernel[4][2] ~^ image[17][19])} + {7'd0,(kernel[4][3] ~^ image[17][20])} + {7'd0,(kernel[4][4] ~^ image[17][21])};
assign out_fmap[13][18][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[13][18])} + {7'd0,(kernel[0][1] ~^ image[13][19])} + {7'd0,(kernel[0][2] ~^ image[13][20])} + {7'd0,(kernel[0][3] ~^ image[13][21])} + {7'd0,(kernel[0][4] ~^ image[13][22])} + {7'd0,(kernel[1][0] ~^ image[14][18])} + {7'd0,(kernel[1][1] ~^ image[14][19])} + {7'd0,(kernel[1][2] ~^ image[14][20])} + {7'd0,(kernel[1][3] ~^ image[14][21])} + {7'd0,(kernel[1][4] ~^ image[14][22])} + {7'd0,(kernel[2][0] ~^ image[15][18])} + {7'd0,(kernel[2][1] ~^ image[15][19])} + {7'd0,(kernel[2][2] ~^ image[15][20])} + {7'd0,(kernel[2][3] ~^ image[15][21])} + {7'd0,(kernel[2][4] ~^ image[15][22])} + {7'd0,(kernel[3][0] ~^ image[16][18])} + {7'd0,(kernel[3][1] ~^ image[16][19])} + {7'd0,(kernel[3][2] ~^ image[16][20])} + {7'd0,(kernel[3][3] ~^ image[16][21])} + {7'd0,(kernel[3][4] ~^ image[16][22])} + {7'd0,(kernel[4][0] ~^ image[17][18])} + {7'd0,(kernel[4][1] ~^ image[17][19])} + {7'd0,(kernel[4][2] ~^ image[17][20])} + {7'd0,(kernel[4][3] ~^ image[17][21])} + {7'd0,(kernel[4][4] ~^ image[17][22])};
assign out_fmap[13][19][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[13][19])} + {7'd0,(kernel[0][1] ~^ image[13][20])} + {7'd0,(kernel[0][2] ~^ image[13][21])} + {7'd0,(kernel[0][3] ~^ image[13][22])} + {7'd0,(kernel[0][4] ~^ image[13][23])} + {7'd0,(kernel[1][0] ~^ image[14][19])} + {7'd0,(kernel[1][1] ~^ image[14][20])} + {7'd0,(kernel[1][2] ~^ image[14][21])} + {7'd0,(kernel[1][3] ~^ image[14][22])} + {7'd0,(kernel[1][4] ~^ image[14][23])} + {7'd0,(kernel[2][0] ~^ image[15][19])} + {7'd0,(kernel[2][1] ~^ image[15][20])} + {7'd0,(kernel[2][2] ~^ image[15][21])} + {7'd0,(kernel[2][3] ~^ image[15][22])} + {7'd0,(kernel[2][4] ~^ image[15][23])} + {7'd0,(kernel[3][0] ~^ image[16][19])} + {7'd0,(kernel[3][1] ~^ image[16][20])} + {7'd0,(kernel[3][2] ~^ image[16][21])} + {7'd0,(kernel[3][3] ~^ image[16][22])} + {7'd0,(kernel[3][4] ~^ image[16][23])} + {7'd0,(kernel[4][0] ~^ image[17][19])} + {7'd0,(kernel[4][1] ~^ image[17][20])} + {7'd0,(kernel[4][2] ~^ image[17][21])} + {7'd0,(kernel[4][3] ~^ image[17][22])} + {7'd0,(kernel[4][4] ~^ image[17][23])};
assign out_fmap[13][20][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[13][20])} + {7'd0,(kernel[0][1] ~^ image[13][21])} + {7'd0,(kernel[0][2] ~^ image[13][22])} + {7'd0,(kernel[0][3] ~^ image[13][23])} + {7'd0,(kernel[0][4] ~^ image[13][24])} + {7'd0,(kernel[1][0] ~^ image[14][20])} + {7'd0,(kernel[1][1] ~^ image[14][21])} + {7'd0,(kernel[1][2] ~^ image[14][22])} + {7'd0,(kernel[1][3] ~^ image[14][23])} + {7'd0,(kernel[1][4] ~^ image[14][24])} + {7'd0,(kernel[2][0] ~^ image[15][20])} + {7'd0,(kernel[2][1] ~^ image[15][21])} + {7'd0,(kernel[2][2] ~^ image[15][22])} + {7'd0,(kernel[2][3] ~^ image[15][23])} + {7'd0,(kernel[2][4] ~^ image[15][24])} + {7'd0,(kernel[3][0] ~^ image[16][20])} + {7'd0,(kernel[3][1] ~^ image[16][21])} + {7'd0,(kernel[3][2] ~^ image[16][22])} + {7'd0,(kernel[3][3] ~^ image[16][23])} + {7'd0,(kernel[3][4] ~^ image[16][24])} + {7'd0,(kernel[4][0] ~^ image[17][20])} + {7'd0,(kernel[4][1] ~^ image[17][21])} + {7'd0,(kernel[4][2] ~^ image[17][22])} + {7'd0,(kernel[4][3] ~^ image[17][23])} + {7'd0,(kernel[4][4] ~^ image[17][24])};
assign out_fmap[13][21][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[13][21])} + {7'd0,(kernel[0][1] ~^ image[13][22])} + {7'd0,(kernel[0][2] ~^ image[13][23])} + {7'd0,(kernel[0][3] ~^ image[13][24])} + {7'd0,(kernel[0][4] ~^ image[13][25])} + {7'd0,(kernel[1][0] ~^ image[14][21])} + {7'd0,(kernel[1][1] ~^ image[14][22])} + {7'd0,(kernel[1][2] ~^ image[14][23])} + {7'd0,(kernel[1][3] ~^ image[14][24])} + {7'd0,(kernel[1][4] ~^ image[14][25])} + {7'd0,(kernel[2][0] ~^ image[15][21])} + {7'd0,(kernel[2][1] ~^ image[15][22])} + {7'd0,(kernel[2][2] ~^ image[15][23])} + {7'd0,(kernel[2][3] ~^ image[15][24])} + {7'd0,(kernel[2][4] ~^ image[15][25])} + {7'd0,(kernel[3][0] ~^ image[16][21])} + {7'd0,(kernel[3][1] ~^ image[16][22])} + {7'd0,(kernel[3][2] ~^ image[16][23])} + {7'd0,(kernel[3][3] ~^ image[16][24])} + {7'd0,(kernel[3][4] ~^ image[16][25])} + {7'd0,(kernel[4][0] ~^ image[17][21])} + {7'd0,(kernel[4][1] ~^ image[17][22])} + {7'd0,(kernel[4][2] ~^ image[17][23])} + {7'd0,(kernel[4][3] ~^ image[17][24])} + {7'd0,(kernel[4][4] ~^ image[17][25])};
assign out_fmap[13][22][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[13][22])} + {7'd0,(kernel[0][1] ~^ image[13][23])} + {7'd0,(kernel[0][2] ~^ image[13][24])} + {7'd0,(kernel[0][3] ~^ image[13][25])} + {7'd0,(kernel[0][4] ~^ image[13][26])} + {7'd0,(kernel[1][0] ~^ image[14][22])} + {7'd0,(kernel[1][1] ~^ image[14][23])} + {7'd0,(kernel[1][2] ~^ image[14][24])} + {7'd0,(kernel[1][3] ~^ image[14][25])} + {7'd0,(kernel[1][4] ~^ image[14][26])} + {7'd0,(kernel[2][0] ~^ image[15][22])} + {7'd0,(kernel[2][1] ~^ image[15][23])} + {7'd0,(kernel[2][2] ~^ image[15][24])} + {7'd0,(kernel[2][3] ~^ image[15][25])} + {7'd0,(kernel[2][4] ~^ image[15][26])} + {7'd0,(kernel[3][0] ~^ image[16][22])} + {7'd0,(kernel[3][1] ~^ image[16][23])} + {7'd0,(kernel[3][2] ~^ image[16][24])} + {7'd0,(kernel[3][3] ~^ image[16][25])} + {7'd0,(kernel[3][4] ~^ image[16][26])} + {7'd0,(kernel[4][0] ~^ image[17][22])} + {7'd0,(kernel[4][1] ~^ image[17][23])} + {7'd0,(kernel[4][2] ~^ image[17][24])} + {7'd0,(kernel[4][3] ~^ image[17][25])} + {7'd0,(kernel[4][4] ~^ image[17][26])};
assign out_fmap[13][23][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[13][23])} + {7'd0,(kernel[0][1] ~^ image[13][24])} + {7'd0,(kernel[0][2] ~^ image[13][25])} + {7'd0,(kernel[0][3] ~^ image[13][26])} + {7'd0,(kernel[0][4] ~^ image[13][27])} + {7'd0,(kernel[1][0] ~^ image[14][23])} + {7'd0,(kernel[1][1] ~^ image[14][24])} + {7'd0,(kernel[1][2] ~^ image[14][25])} + {7'd0,(kernel[1][3] ~^ image[14][26])} + {7'd0,(kernel[1][4] ~^ image[14][27])} + {7'd0,(kernel[2][0] ~^ image[15][23])} + {7'd0,(kernel[2][1] ~^ image[15][24])} + {7'd0,(kernel[2][2] ~^ image[15][25])} + {7'd0,(kernel[2][3] ~^ image[15][26])} + {7'd0,(kernel[2][4] ~^ image[15][27])} + {7'd0,(kernel[3][0] ~^ image[16][23])} + {7'd0,(kernel[3][1] ~^ image[16][24])} + {7'd0,(kernel[3][2] ~^ image[16][25])} + {7'd0,(kernel[3][3] ~^ image[16][26])} + {7'd0,(kernel[3][4] ~^ image[16][27])} + {7'd0,(kernel[4][0] ~^ image[17][23])} + {7'd0,(kernel[4][1] ~^ image[17][24])} + {7'd0,(kernel[4][2] ~^ image[17][25])} + {7'd0,(kernel[4][3] ~^ image[17][26])} + {7'd0,(kernel[4][4] ~^ image[17][27])};
assign out_fmap[14][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[14][0])} + {7'd0,(kernel[0][1] ~^ image[14][1])} + {7'd0,(kernel[0][2] ~^ image[14][2])} + {7'd0,(kernel[0][3] ~^ image[14][3])} + {7'd0,(kernel[0][4] ~^ image[14][4])} + {7'd0,(kernel[1][0] ~^ image[15][0])} + {7'd0,(kernel[1][1] ~^ image[15][1])} + {7'd0,(kernel[1][2] ~^ image[15][2])} + {7'd0,(kernel[1][3] ~^ image[15][3])} + {7'd0,(kernel[1][4] ~^ image[15][4])} + {7'd0,(kernel[2][0] ~^ image[16][0])} + {7'd0,(kernel[2][1] ~^ image[16][1])} + {7'd0,(kernel[2][2] ~^ image[16][2])} + {7'd0,(kernel[2][3] ~^ image[16][3])} + {7'd0,(kernel[2][4] ~^ image[16][4])} + {7'd0,(kernel[3][0] ~^ image[17][0])} + {7'd0,(kernel[3][1] ~^ image[17][1])} + {7'd0,(kernel[3][2] ~^ image[17][2])} + {7'd0,(kernel[3][3] ~^ image[17][3])} + {7'd0,(kernel[3][4] ~^ image[17][4])} + {7'd0,(kernel[4][0] ~^ image[18][0])} + {7'd0,(kernel[4][1] ~^ image[18][1])} + {7'd0,(kernel[4][2] ~^ image[18][2])} + {7'd0,(kernel[4][3] ~^ image[18][3])} + {7'd0,(kernel[4][4] ~^ image[18][4])};
assign out_fmap[14][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[14][1])} + {7'd0,(kernel[0][1] ~^ image[14][2])} + {7'd0,(kernel[0][2] ~^ image[14][3])} + {7'd0,(kernel[0][3] ~^ image[14][4])} + {7'd0,(kernel[0][4] ~^ image[14][5])} + {7'd0,(kernel[1][0] ~^ image[15][1])} + {7'd0,(kernel[1][1] ~^ image[15][2])} + {7'd0,(kernel[1][2] ~^ image[15][3])} + {7'd0,(kernel[1][3] ~^ image[15][4])} + {7'd0,(kernel[1][4] ~^ image[15][5])} + {7'd0,(kernel[2][0] ~^ image[16][1])} + {7'd0,(kernel[2][1] ~^ image[16][2])} + {7'd0,(kernel[2][2] ~^ image[16][3])} + {7'd0,(kernel[2][3] ~^ image[16][4])} + {7'd0,(kernel[2][4] ~^ image[16][5])} + {7'd0,(kernel[3][0] ~^ image[17][1])} + {7'd0,(kernel[3][1] ~^ image[17][2])} + {7'd0,(kernel[3][2] ~^ image[17][3])} + {7'd0,(kernel[3][3] ~^ image[17][4])} + {7'd0,(kernel[3][4] ~^ image[17][5])} + {7'd0,(kernel[4][0] ~^ image[18][1])} + {7'd0,(kernel[4][1] ~^ image[18][2])} + {7'd0,(kernel[4][2] ~^ image[18][3])} + {7'd0,(kernel[4][3] ~^ image[18][4])} + {7'd0,(kernel[4][4] ~^ image[18][5])};
assign out_fmap[14][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[14][2])} + {7'd0,(kernel[0][1] ~^ image[14][3])} + {7'd0,(kernel[0][2] ~^ image[14][4])} + {7'd0,(kernel[0][3] ~^ image[14][5])} + {7'd0,(kernel[0][4] ~^ image[14][6])} + {7'd0,(kernel[1][0] ~^ image[15][2])} + {7'd0,(kernel[1][1] ~^ image[15][3])} + {7'd0,(kernel[1][2] ~^ image[15][4])} + {7'd0,(kernel[1][3] ~^ image[15][5])} + {7'd0,(kernel[1][4] ~^ image[15][6])} + {7'd0,(kernel[2][0] ~^ image[16][2])} + {7'd0,(kernel[2][1] ~^ image[16][3])} + {7'd0,(kernel[2][2] ~^ image[16][4])} + {7'd0,(kernel[2][3] ~^ image[16][5])} + {7'd0,(kernel[2][4] ~^ image[16][6])} + {7'd0,(kernel[3][0] ~^ image[17][2])} + {7'd0,(kernel[3][1] ~^ image[17][3])} + {7'd0,(kernel[3][2] ~^ image[17][4])} + {7'd0,(kernel[3][3] ~^ image[17][5])} + {7'd0,(kernel[3][4] ~^ image[17][6])} + {7'd0,(kernel[4][0] ~^ image[18][2])} + {7'd0,(kernel[4][1] ~^ image[18][3])} + {7'd0,(kernel[4][2] ~^ image[18][4])} + {7'd0,(kernel[4][3] ~^ image[18][5])} + {7'd0,(kernel[4][4] ~^ image[18][6])};
assign out_fmap[14][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[14][3])} + {7'd0,(kernel[0][1] ~^ image[14][4])} + {7'd0,(kernel[0][2] ~^ image[14][5])} + {7'd0,(kernel[0][3] ~^ image[14][6])} + {7'd0,(kernel[0][4] ~^ image[14][7])} + {7'd0,(kernel[1][0] ~^ image[15][3])} + {7'd0,(kernel[1][1] ~^ image[15][4])} + {7'd0,(kernel[1][2] ~^ image[15][5])} + {7'd0,(kernel[1][3] ~^ image[15][6])} + {7'd0,(kernel[1][4] ~^ image[15][7])} + {7'd0,(kernel[2][0] ~^ image[16][3])} + {7'd0,(kernel[2][1] ~^ image[16][4])} + {7'd0,(kernel[2][2] ~^ image[16][5])} + {7'd0,(kernel[2][3] ~^ image[16][6])} + {7'd0,(kernel[2][4] ~^ image[16][7])} + {7'd0,(kernel[3][0] ~^ image[17][3])} + {7'd0,(kernel[3][1] ~^ image[17][4])} + {7'd0,(kernel[3][2] ~^ image[17][5])} + {7'd0,(kernel[3][3] ~^ image[17][6])} + {7'd0,(kernel[3][4] ~^ image[17][7])} + {7'd0,(kernel[4][0] ~^ image[18][3])} + {7'd0,(kernel[4][1] ~^ image[18][4])} + {7'd0,(kernel[4][2] ~^ image[18][5])} + {7'd0,(kernel[4][3] ~^ image[18][6])} + {7'd0,(kernel[4][4] ~^ image[18][7])};
assign out_fmap[14][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[14][4])} + {7'd0,(kernel[0][1] ~^ image[14][5])} + {7'd0,(kernel[0][2] ~^ image[14][6])} + {7'd0,(kernel[0][3] ~^ image[14][7])} + {7'd0,(kernel[0][4] ~^ image[14][8])} + {7'd0,(kernel[1][0] ~^ image[15][4])} + {7'd0,(kernel[1][1] ~^ image[15][5])} + {7'd0,(kernel[1][2] ~^ image[15][6])} + {7'd0,(kernel[1][3] ~^ image[15][7])} + {7'd0,(kernel[1][4] ~^ image[15][8])} + {7'd0,(kernel[2][0] ~^ image[16][4])} + {7'd0,(kernel[2][1] ~^ image[16][5])} + {7'd0,(kernel[2][2] ~^ image[16][6])} + {7'd0,(kernel[2][3] ~^ image[16][7])} + {7'd0,(kernel[2][4] ~^ image[16][8])} + {7'd0,(kernel[3][0] ~^ image[17][4])} + {7'd0,(kernel[3][1] ~^ image[17][5])} + {7'd0,(kernel[3][2] ~^ image[17][6])} + {7'd0,(kernel[3][3] ~^ image[17][7])} + {7'd0,(kernel[3][4] ~^ image[17][8])} + {7'd0,(kernel[4][0] ~^ image[18][4])} + {7'd0,(kernel[4][1] ~^ image[18][5])} + {7'd0,(kernel[4][2] ~^ image[18][6])} + {7'd0,(kernel[4][3] ~^ image[18][7])} + {7'd0,(kernel[4][4] ~^ image[18][8])};
assign out_fmap[14][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[14][5])} + {7'd0,(kernel[0][1] ~^ image[14][6])} + {7'd0,(kernel[0][2] ~^ image[14][7])} + {7'd0,(kernel[0][3] ~^ image[14][8])} + {7'd0,(kernel[0][4] ~^ image[14][9])} + {7'd0,(kernel[1][0] ~^ image[15][5])} + {7'd0,(kernel[1][1] ~^ image[15][6])} + {7'd0,(kernel[1][2] ~^ image[15][7])} + {7'd0,(kernel[1][3] ~^ image[15][8])} + {7'd0,(kernel[1][4] ~^ image[15][9])} + {7'd0,(kernel[2][0] ~^ image[16][5])} + {7'd0,(kernel[2][1] ~^ image[16][6])} + {7'd0,(kernel[2][2] ~^ image[16][7])} + {7'd0,(kernel[2][3] ~^ image[16][8])} + {7'd0,(kernel[2][4] ~^ image[16][9])} + {7'd0,(kernel[3][0] ~^ image[17][5])} + {7'd0,(kernel[3][1] ~^ image[17][6])} + {7'd0,(kernel[3][2] ~^ image[17][7])} + {7'd0,(kernel[3][3] ~^ image[17][8])} + {7'd0,(kernel[3][4] ~^ image[17][9])} + {7'd0,(kernel[4][0] ~^ image[18][5])} + {7'd0,(kernel[4][1] ~^ image[18][6])} + {7'd0,(kernel[4][2] ~^ image[18][7])} + {7'd0,(kernel[4][3] ~^ image[18][8])} + {7'd0,(kernel[4][4] ~^ image[18][9])};
assign out_fmap[14][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[14][6])} + {7'd0,(kernel[0][1] ~^ image[14][7])} + {7'd0,(kernel[0][2] ~^ image[14][8])} + {7'd0,(kernel[0][3] ~^ image[14][9])} + {7'd0,(kernel[0][4] ~^ image[14][10])} + {7'd0,(kernel[1][0] ~^ image[15][6])} + {7'd0,(kernel[1][1] ~^ image[15][7])} + {7'd0,(kernel[1][2] ~^ image[15][8])} + {7'd0,(kernel[1][3] ~^ image[15][9])} + {7'd0,(kernel[1][4] ~^ image[15][10])} + {7'd0,(kernel[2][0] ~^ image[16][6])} + {7'd0,(kernel[2][1] ~^ image[16][7])} + {7'd0,(kernel[2][2] ~^ image[16][8])} + {7'd0,(kernel[2][3] ~^ image[16][9])} + {7'd0,(kernel[2][4] ~^ image[16][10])} + {7'd0,(kernel[3][0] ~^ image[17][6])} + {7'd0,(kernel[3][1] ~^ image[17][7])} + {7'd0,(kernel[3][2] ~^ image[17][8])} + {7'd0,(kernel[3][3] ~^ image[17][9])} + {7'd0,(kernel[3][4] ~^ image[17][10])} + {7'd0,(kernel[4][0] ~^ image[18][6])} + {7'd0,(kernel[4][1] ~^ image[18][7])} + {7'd0,(kernel[4][2] ~^ image[18][8])} + {7'd0,(kernel[4][3] ~^ image[18][9])} + {7'd0,(kernel[4][4] ~^ image[18][10])};
assign out_fmap[14][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[14][7])} + {7'd0,(kernel[0][1] ~^ image[14][8])} + {7'd0,(kernel[0][2] ~^ image[14][9])} + {7'd0,(kernel[0][3] ~^ image[14][10])} + {7'd0,(kernel[0][4] ~^ image[14][11])} + {7'd0,(kernel[1][0] ~^ image[15][7])} + {7'd0,(kernel[1][1] ~^ image[15][8])} + {7'd0,(kernel[1][2] ~^ image[15][9])} + {7'd0,(kernel[1][3] ~^ image[15][10])} + {7'd0,(kernel[1][4] ~^ image[15][11])} + {7'd0,(kernel[2][0] ~^ image[16][7])} + {7'd0,(kernel[2][1] ~^ image[16][8])} + {7'd0,(kernel[2][2] ~^ image[16][9])} + {7'd0,(kernel[2][3] ~^ image[16][10])} + {7'd0,(kernel[2][4] ~^ image[16][11])} + {7'd0,(kernel[3][0] ~^ image[17][7])} + {7'd0,(kernel[3][1] ~^ image[17][8])} + {7'd0,(kernel[3][2] ~^ image[17][9])} + {7'd0,(kernel[3][3] ~^ image[17][10])} + {7'd0,(kernel[3][4] ~^ image[17][11])} + {7'd0,(kernel[4][0] ~^ image[18][7])} + {7'd0,(kernel[4][1] ~^ image[18][8])} + {7'd0,(kernel[4][2] ~^ image[18][9])} + {7'd0,(kernel[4][3] ~^ image[18][10])} + {7'd0,(kernel[4][4] ~^ image[18][11])};
assign out_fmap[14][8][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[14][8])} + {7'd0,(kernel[0][1] ~^ image[14][9])} + {7'd0,(kernel[0][2] ~^ image[14][10])} + {7'd0,(kernel[0][3] ~^ image[14][11])} + {7'd0,(kernel[0][4] ~^ image[14][12])} + {7'd0,(kernel[1][0] ~^ image[15][8])} + {7'd0,(kernel[1][1] ~^ image[15][9])} + {7'd0,(kernel[1][2] ~^ image[15][10])} + {7'd0,(kernel[1][3] ~^ image[15][11])} + {7'd0,(kernel[1][4] ~^ image[15][12])} + {7'd0,(kernel[2][0] ~^ image[16][8])} + {7'd0,(kernel[2][1] ~^ image[16][9])} + {7'd0,(kernel[2][2] ~^ image[16][10])} + {7'd0,(kernel[2][3] ~^ image[16][11])} + {7'd0,(kernel[2][4] ~^ image[16][12])} + {7'd0,(kernel[3][0] ~^ image[17][8])} + {7'd0,(kernel[3][1] ~^ image[17][9])} + {7'd0,(kernel[3][2] ~^ image[17][10])} + {7'd0,(kernel[3][3] ~^ image[17][11])} + {7'd0,(kernel[3][4] ~^ image[17][12])} + {7'd0,(kernel[4][0] ~^ image[18][8])} + {7'd0,(kernel[4][1] ~^ image[18][9])} + {7'd0,(kernel[4][2] ~^ image[18][10])} + {7'd0,(kernel[4][3] ~^ image[18][11])} + {7'd0,(kernel[4][4] ~^ image[18][12])};
assign out_fmap[14][9][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[14][9])} + {7'd0,(kernel[0][1] ~^ image[14][10])} + {7'd0,(kernel[0][2] ~^ image[14][11])} + {7'd0,(kernel[0][3] ~^ image[14][12])} + {7'd0,(kernel[0][4] ~^ image[14][13])} + {7'd0,(kernel[1][0] ~^ image[15][9])} + {7'd0,(kernel[1][1] ~^ image[15][10])} + {7'd0,(kernel[1][2] ~^ image[15][11])} + {7'd0,(kernel[1][3] ~^ image[15][12])} + {7'd0,(kernel[1][4] ~^ image[15][13])} + {7'd0,(kernel[2][0] ~^ image[16][9])} + {7'd0,(kernel[2][1] ~^ image[16][10])} + {7'd0,(kernel[2][2] ~^ image[16][11])} + {7'd0,(kernel[2][3] ~^ image[16][12])} + {7'd0,(kernel[2][4] ~^ image[16][13])} + {7'd0,(kernel[3][0] ~^ image[17][9])} + {7'd0,(kernel[3][1] ~^ image[17][10])} + {7'd0,(kernel[3][2] ~^ image[17][11])} + {7'd0,(kernel[3][3] ~^ image[17][12])} + {7'd0,(kernel[3][4] ~^ image[17][13])} + {7'd0,(kernel[4][0] ~^ image[18][9])} + {7'd0,(kernel[4][1] ~^ image[18][10])} + {7'd0,(kernel[4][2] ~^ image[18][11])} + {7'd0,(kernel[4][3] ~^ image[18][12])} + {7'd0,(kernel[4][4] ~^ image[18][13])};
assign out_fmap[14][10][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[14][10])} + {7'd0,(kernel[0][1] ~^ image[14][11])} + {7'd0,(kernel[0][2] ~^ image[14][12])} + {7'd0,(kernel[0][3] ~^ image[14][13])} + {7'd0,(kernel[0][4] ~^ image[14][14])} + {7'd0,(kernel[1][0] ~^ image[15][10])} + {7'd0,(kernel[1][1] ~^ image[15][11])} + {7'd0,(kernel[1][2] ~^ image[15][12])} + {7'd0,(kernel[1][3] ~^ image[15][13])} + {7'd0,(kernel[1][4] ~^ image[15][14])} + {7'd0,(kernel[2][0] ~^ image[16][10])} + {7'd0,(kernel[2][1] ~^ image[16][11])} + {7'd0,(kernel[2][2] ~^ image[16][12])} + {7'd0,(kernel[2][3] ~^ image[16][13])} + {7'd0,(kernel[2][4] ~^ image[16][14])} + {7'd0,(kernel[3][0] ~^ image[17][10])} + {7'd0,(kernel[3][1] ~^ image[17][11])} + {7'd0,(kernel[3][2] ~^ image[17][12])} + {7'd0,(kernel[3][3] ~^ image[17][13])} + {7'd0,(kernel[3][4] ~^ image[17][14])} + {7'd0,(kernel[4][0] ~^ image[18][10])} + {7'd0,(kernel[4][1] ~^ image[18][11])} + {7'd0,(kernel[4][2] ~^ image[18][12])} + {7'd0,(kernel[4][3] ~^ image[18][13])} + {7'd0,(kernel[4][4] ~^ image[18][14])};
assign out_fmap[14][11][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[14][11])} + {7'd0,(kernel[0][1] ~^ image[14][12])} + {7'd0,(kernel[0][2] ~^ image[14][13])} + {7'd0,(kernel[0][3] ~^ image[14][14])} + {7'd0,(kernel[0][4] ~^ image[14][15])} + {7'd0,(kernel[1][0] ~^ image[15][11])} + {7'd0,(kernel[1][1] ~^ image[15][12])} + {7'd0,(kernel[1][2] ~^ image[15][13])} + {7'd0,(kernel[1][3] ~^ image[15][14])} + {7'd0,(kernel[1][4] ~^ image[15][15])} + {7'd0,(kernel[2][0] ~^ image[16][11])} + {7'd0,(kernel[2][1] ~^ image[16][12])} + {7'd0,(kernel[2][2] ~^ image[16][13])} + {7'd0,(kernel[2][3] ~^ image[16][14])} + {7'd0,(kernel[2][4] ~^ image[16][15])} + {7'd0,(kernel[3][0] ~^ image[17][11])} + {7'd0,(kernel[3][1] ~^ image[17][12])} + {7'd0,(kernel[3][2] ~^ image[17][13])} + {7'd0,(kernel[3][3] ~^ image[17][14])} + {7'd0,(kernel[3][4] ~^ image[17][15])} + {7'd0,(kernel[4][0] ~^ image[18][11])} + {7'd0,(kernel[4][1] ~^ image[18][12])} + {7'd0,(kernel[4][2] ~^ image[18][13])} + {7'd0,(kernel[4][3] ~^ image[18][14])} + {7'd0,(kernel[4][4] ~^ image[18][15])};
assign out_fmap[14][12][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[14][12])} + {7'd0,(kernel[0][1] ~^ image[14][13])} + {7'd0,(kernel[0][2] ~^ image[14][14])} + {7'd0,(kernel[0][3] ~^ image[14][15])} + {7'd0,(kernel[0][4] ~^ image[14][16])} + {7'd0,(kernel[1][0] ~^ image[15][12])} + {7'd0,(kernel[1][1] ~^ image[15][13])} + {7'd0,(kernel[1][2] ~^ image[15][14])} + {7'd0,(kernel[1][3] ~^ image[15][15])} + {7'd0,(kernel[1][4] ~^ image[15][16])} + {7'd0,(kernel[2][0] ~^ image[16][12])} + {7'd0,(kernel[2][1] ~^ image[16][13])} + {7'd0,(kernel[2][2] ~^ image[16][14])} + {7'd0,(kernel[2][3] ~^ image[16][15])} + {7'd0,(kernel[2][4] ~^ image[16][16])} + {7'd0,(kernel[3][0] ~^ image[17][12])} + {7'd0,(kernel[3][1] ~^ image[17][13])} + {7'd0,(kernel[3][2] ~^ image[17][14])} + {7'd0,(kernel[3][3] ~^ image[17][15])} + {7'd0,(kernel[3][4] ~^ image[17][16])} + {7'd0,(kernel[4][0] ~^ image[18][12])} + {7'd0,(kernel[4][1] ~^ image[18][13])} + {7'd0,(kernel[4][2] ~^ image[18][14])} + {7'd0,(kernel[4][3] ~^ image[18][15])} + {7'd0,(kernel[4][4] ~^ image[18][16])};
assign out_fmap[14][13][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[14][13])} + {7'd0,(kernel[0][1] ~^ image[14][14])} + {7'd0,(kernel[0][2] ~^ image[14][15])} + {7'd0,(kernel[0][3] ~^ image[14][16])} + {7'd0,(kernel[0][4] ~^ image[14][17])} + {7'd0,(kernel[1][0] ~^ image[15][13])} + {7'd0,(kernel[1][1] ~^ image[15][14])} + {7'd0,(kernel[1][2] ~^ image[15][15])} + {7'd0,(kernel[1][3] ~^ image[15][16])} + {7'd0,(kernel[1][4] ~^ image[15][17])} + {7'd0,(kernel[2][0] ~^ image[16][13])} + {7'd0,(kernel[2][1] ~^ image[16][14])} + {7'd0,(kernel[2][2] ~^ image[16][15])} + {7'd0,(kernel[2][3] ~^ image[16][16])} + {7'd0,(kernel[2][4] ~^ image[16][17])} + {7'd0,(kernel[3][0] ~^ image[17][13])} + {7'd0,(kernel[3][1] ~^ image[17][14])} + {7'd0,(kernel[3][2] ~^ image[17][15])} + {7'd0,(kernel[3][3] ~^ image[17][16])} + {7'd0,(kernel[3][4] ~^ image[17][17])} + {7'd0,(kernel[4][0] ~^ image[18][13])} + {7'd0,(kernel[4][1] ~^ image[18][14])} + {7'd0,(kernel[4][2] ~^ image[18][15])} + {7'd0,(kernel[4][3] ~^ image[18][16])} + {7'd0,(kernel[4][4] ~^ image[18][17])};
assign out_fmap[14][14][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[14][14])} + {7'd0,(kernel[0][1] ~^ image[14][15])} + {7'd0,(kernel[0][2] ~^ image[14][16])} + {7'd0,(kernel[0][3] ~^ image[14][17])} + {7'd0,(kernel[0][4] ~^ image[14][18])} + {7'd0,(kernel[1][0] ~^ image[15][14])} + {7'd0,(kernel[1][1] ~^ image[15][15])} + {7'd0,(kernel[1][2] ~^ image[15][16])} + {7'd0,(kernel[1][3] ~^ image[15][17])} + {7'd0,(kernel[1][4] ~^ image[15][18])} + {7'd0,(kernel[2][0] ~^ image[16][14])} + {7'd0,(kernel[2][1] ~^ image[16][15])} + {7'd0,(kernel[2][2] ~^ image[16][16])} + {7'd0,(kernel[2][3] ~^ image[16][17])} + {7'd0,(kernel[2][4] ~^ image[16][18])} + {7'd0,(kernel[3][0] ~^ image[17][14])} + {7'd0,(kernel[3][1] ~^ image[17][15])} + {7'd0,(kernel[3][2] ~^ image[17][16])} + {7'd0,(kernel[3][3] ~^ image[17][17])} + {7'd0,(kernel[3][4] ~^ image[17][18])} + {7'd0,(kernel[4][0] ~^ image[18][14])} + {7'd0,(kernel[4][1] ~^ image[18][15])} + {7'd0,(kernel[4][2] ~^ image[18][16])} + {7'd0,(kernel[4][3] ~^ image[18][17])} + {7'd0,(kernel[4][4] ~^ image[18][18])};
assign out_fmap[14][15][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[14][15])} + {7'd0,(kernel[0][1] ~^ image[14][16])} + {7'd0,(kernel[0][2] ~^ image[14][17])} + {7'd0,(kernel[0][3] ~^ image[14][18])} + {7'd0,(kernel[0][4] ~^ image[14][19])} + {7'd0,(kernel[1][0] ~^ image[15][15])} + {7'd0,(kernel[1][1] ~^ image[15][16])} + {7'd0,(kernel[1][2] ~^ image[15][17])} + {7'd0,(kernel[1][3] ~^ image[15][18])} + {7'd0,(kernel[1][4] ~^ image[15][19])} + {7'd0,(kernel[2][0] ~^ image[16][15])} + {7'd0,(kernel[2][1] ~^ image[16][16])} + {7'd0,(kernel[2][2] ~^ image[16][17])} + {7'd0,(kernel[2][3] ~^ image[16][18])} + {7'd0,(kernel[2][4] ~^ image[16][19])} + {7'd0,(kernel[3][0] ~^ image[17][15])} + {7'd0,(kernel[3][1] ~^ image[17][16])} + {7'd0,(kernel[3][2] ~^ image[17][17])} + {7'd0,(kernel[3][3] ~^ image[17][18])} + {7'd0,(kernel[3][4] ~^ image[17][19])} + {7'd0,(kernel[4][0] ~^ image[18][15])} + {7'd0,(kernel[4][1] ~^ image[18][16])} + {7'd0,(kernel[4][2] ~^ image[18][17])} + {7'd0,(kernel[4][3] ~^ image[18][18])} + {7'd0,(kernel[4][4] ~^ image[18][19])};
assign out_fmap[14][16][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[14][16])} + {7'd0,(kernel[0][1] ~^ image[14][17])} + {7'd0,(kernel[0][2] ~^ image[14][18])} + {7'd0,(kernel[0][3] ~^ image[14][19])} + {7'd0,(kernel[0][4] ~^ image[14][20])} + {7'd0,(kernel[1][0] ~^ image[15][16])} + {7'd0,(kernel[1][1] ~^ image[15][17])} + {7'd0,(kernel[1][2] ~^ image[15][18])} + {7'd0,(kernel[1][3] ~^ image[15][19])} + {7'd0,(kernel[1][4] ~^ image[15][20])} + {7'd0,(kernel[2][0] ~^ image[16][16])} + {7'd0,(kernel[2][1] ~^ image[16][17])} + {7'd0,(kernel[2][2] ~^ image[16][18])} + {7'd0,(kernel[2][3] ~^ image[16][19])} + {7'd0,(kernel[2][4] ~^ image[16][20])} + {7'd0,(kernel[3][0] ~^ image[17][16])} + {7'd0,(kernel[3][1] ~^ image[17][17])} + {7'd0,(kernel[3][2] ~^ image[17][18])} + {7'd0,(kernel[3][3] ~^ image[17][19])} + {7'd0,(kernel[3][4] ~^ image[17][20])} + {7'd0,(kernel[4][0] ~^ image[18][16])} + {7'd0,(kernel[4][1] ~^ image[18][17])} + {7'd0,(kernel[4][2] ~^ image[18][18])} + {7'd0,(kernel[4][3] ~^ image[18][19])} + {7'd0,(kernel[4][4] ~^ image[18][20])};
assign out_fmap[14][17][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[14][17])} + {7'd0,(kernel[0][1] ~^ image[14][18])} + {7'd0,(kernel[0][2] ~^ image[14][19])} + {7'd0,(kernel[0][3] ~^ image[14][20])} + {7'd0,(kernel[0][4] ~^ image[14][21])} + {7'd0,(kernel[1][0] ~^ image[15][17])} + {7'd0,(kernel[1][1] ~^ image[15][18])} + {7'd0,(kernel[1][2] ~^ image[15][19])} + {7'd0,(kernel[1][3] ~^ image[15][20])} + {7'd0,(kernel[1][4] ~^ image[15][21])} + {7'd0,(kernel[2][0] ~^ image[16][17])} + {7'd0,(kernel[2][1] ~^ image[16][18])} + {7'd0,(kernel[2][2] ~^ image[16][19])} + {7'd0,(kernel[2][3] ~^ image[16][20])} + {7'd0,(kernel[2][4] ~^ image[16][21])} + {7'd0,(kernel[3][0] ~^ image[17][17])} + {7'd0,(kernel[3][1] ~^ image[17][18])} + {7'd0,(kernel[3][2] ~^ image[17][19])} + {7'd0,(kernel[3][3] ~^ image[17][20])} + {7'd0,(kernel[3][4] ~^ image[17][21])} + {7'd0,(kernel[4][0] ~^ image[18][17])} + {7'd0,(kernel[4][1] ~^ image[18][18])} + {7'd0,(kernel[4][2] ~^ image[18][19])} + {7'd0,(kernel[4][3] ~^ image[18][20])} + {7'd0,(kernel[4][4] ~^ image[18][21])};
assign out_fmap[14][18][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[14][18])} + {7'd0,(kernel[0][1] ~^ image[14][19])} + {7'd0,(kernel[0][2] ~^ image[14][20])} + {7'd0,(kernel[0][3] ~^ image[14][21])} + {7'd0,(kernel[0][4] ~^ image[14][22])} + {7'd0,(kernel[1][0] ~^ image[15][18])} + {7'd0,(kernel[1][1] ~^ image[15][19])} + {7'd0,(kernel[1][2] ~^ image[15][20])} + {7'd0,(kernel[1][3] ~^ image[15][21])} + {7'd0,(kernel[1][4] ~^ image[15][22])} + {7'd0,(kernel[2][0] ~^ image[16][18])} + {7'd0,(kernel[2][1] ~^ image[16][19])} + {7'd0,(kernel[2][2] ~^ image[16][20])} + {7'd0,(kernel[2][3] ~^ image[16][21])} + {7'd0,(kernel[2][4] ~^ image[16][22])} + {7'd0,(kernel[3][0] ~^ image[17][18])} + {7'd0,(kernel[3][1] ~^ image[17][19])} + {7'd0,(kernel[3][2] ~^ image[17][20])} + {7'd0,(kernel[3][3] ~^ image[17][21])} + {7'd0,(kernel[3][4] ~^ image[17][22])} + {7'd0,(kernel[4][0] ~^ image[18][18])} + {7'd0,(kernel[4][1] ~^ image[18][19])} + {7'd0,(kernel[4][2] ~^ image[18][20])} + {7'd0,(kernel[4][3] ~^ image[18][21])} + {7'd0,(kernel[4][4] ~^ image[18][22])};
assign out_fmap[14][19][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[14][19])} + {7'd0,(kernel[0][1] ~^ image[14][20])} + {7'd0,(kernel[0][2] ~^ image[14][21])} + {7'd0,(kernel[0][3] ~^ image[14][22])} + {7'd0,(kernel[0][4] ~^ image[14][23])} + {7'd0,(kernel[1][0] ~^ image[15][19])} + {7'd0,(kernel[1][1] ~^ image[15][20])} + {7'd0,(kernel[1][2] ~^ image[15][21])} + {7'd0,(kernel[1][3] ~^ image[15][22])} + {7'd0,(kernel[1][4] ~^ image[15][23])} + {7'd0,(kernel[2][0] ~^ image[16][19])} + {7'd0,(kernel[2][1] ~^ image[16][20])} + {7'd0,(kernel[2][2] ~^ image[16][21])} + {7'd0,(kernel[2][3] ~^ image[16][22])} + {7'd0,(kernel[2][4] ~^ image[16][23])} + {7'd0,(kernel[3][0] ~^ image[17][19])} + {7'd0,(kernel[3][1] ~^ image[17][20])} + {7'd0,(kernel[3][2] ~^ image[17][21])} + {7'd0,(kernel[3][3] ~^ image[17][22])} + {7'd0,(kernel[3][4] ~^ image[17][23])} + {7'd0,(kernel[4][0] ~^ image[18][19])} + {7'd0,(kernel[4][1] ~^ image[18][20])} + {7'd0,(kernel[4][2] ~^ image[18][21])} + {7'd0,(kernel[4][3] ~^ image[18][22])} + {7'd0,(kernel[4][4] ~^ image[18][23])};
assign out_fmap[14][20][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[14][20])} + {7'd0,(kernel[0][1] ~^ image[14][21])} + {7'd0,(kernel[0][2] ~^ image[14][22])} + {7'd0,(kernel[0][3] ~^ image[14][23])} + {7'd0,(kernel[0][4] ~^ image[14][24])} + {7'd0,(kernel[1][0] ~^ image[15][20])} + {7'd0,(kernel[1][1] ~^ image[15][21])} + {7'd0,(kernel[1][2] ~^ image[15][22])} + {7'd0,(kernel[1][3] ~^ image[15][23])} + {7'd0,(kernel[1][4] ~^ image[15][24])} + {7'd0,(kernel[2][0] ~^ image[16][20])} + {7'd0,(kernel[2][1] ~^ image[16][21])} + {7'd0,(kernel[2][2] ~^ image[16][22])} + {7'd0,(kernel[2][3] ~^ image[16][23])} + {7'd0,(kernel[2][4] ~^ image[16][24])} + {7'd0,(kernel[3][0] ~^ image[17][20])} + {7'd0,(kernel[3][1] ~^ image[17][21])} + {7'd0,(kernel[3][2] ~^ image[17][22])} + {7'd0,(kernel[3][3] ~^ image[17][23])} + {7'd0,(kernel[3][4] ~^ image[17][24])} + {7'd0,(kernel[4][0] ~^ image[18][20])} + {7'd0,(kernel[4][1] ~^ image[18][21])} + {7'd0,(kernel[4][2] ~^ image[18][22])} + {7'd0,(kernel[4][3] ~^ image[18][23])} + {7'd0,(kernel[4][4] ~^ image[18][24])};
assign out_fmap[14][21][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[14][21])} + {7'd0,(kernel[0][1] ~^ image[14][22])} + {7'd0,(kernel[0][2] ~^ image[14][23])} + {7'd0,(kernel[0][3] ~^ image[14][24])} + {7'd0,(kernel[0][4] ~^ image[14][25])} + {7'd0,(kernel[1][0] ~^ image[15][21])} + {7'd0,(kernel[1][1] ~^ image[15][22])} + {7'd0,(kernel[1][2] ~^ image[15][23])} + {7'd0,(kernel[1][3] ~^ image[15][24])} + {7'd0,(kernel[1][4] ~^ image[15][25])} + {7'd0,(kernel[2][0] ~^ image[16][21])} + {7'd0,(kernel[2][1] ~^ image[16][22])} + {7'd0,(kernel[2][2] ~^ image[16][23])} + {7'd0,(kernel[2][3] ~^ image[16][24])} + {7'd0,(kernel[2][4] ~^ image[16][25])} + {7'd0,(kernel[3][0] ~^ image[17][21])} + {7'd0,(kernel[3][1] ~^ image[17][22])} + {7'd0,(kernel[3][2] ~^ image[17][23])} + {7'd0,(kernel[3][3] ~^ image[17][24])} + {7'd0,(kernel[3][4] ~^ image[17][25])} + {7'd0,(kernel[4][0] ~^ image[18][21])} + {7'd0,(kernel[4][1] ~^ image[18][22])} + {7'd0,(kernel[4][2] ~^ image[18][23])} + {7'd0,(kernel[4][3] ~^ image[18][24])} + {7'd0,(kernel[4][4] ~^ image[18][25])};
assign out_fmap[14][22][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[14][22])} + {7'd0,(kernel[0][1] ~^ image[14][23])} + {7'd0,(kernel[0][2] ~^ image[14][24])} + {7'd0,(kernel[0][3] ~^ image[14][25])} + {7'd0,(kernel[0][4] ~^ image[14][26])} + {7'd0,(kernel[1][0] ~^ image[15][22])} + {7'd0,(kernel[1][1] ~^ image[15][23])} + {7'd0,(kernel[1][2] ~^ image[15][24])} + {7'd0,(kernel[1][3] ~^ image[15][25])} + {7'd0,(kernel[1][4] ~^ image[15][26])} + {7'd0,(kernel[2][0] ~^ image[16][22])} + {7'd0,(kernel[2][1] ~^ image[16][23])} + {7'd0,(kernel[2][2] ~^ image[16][24])} + {7'd0,(kernel[2][3] ~^ image[16][25])} + {7'd0,(kernel[2][4] ~^ image[16][26])} + {7'd0,(kernel[3][0] ~^ image[17][22])} + {7'd0,(kernel[3][1] ~^ image[17][23])} + {7'd0,(kernel[3][2] ~^ image[17][24])} + {7'd0,(kernel[3][3] ~^ image[17][25])} + {7'd0,(kernel[3][4] ~^ image[17][26])} + {7'd0,(kernel[4][0] ~^ image[18][22])} + {7'd0,(kernel[4][1] ~^ image[18][23])} + {7'd0,(kernel[4][2] ~^ image[18][24])} + {7'd0,(kernel[4][3] ~^ image[18][25])} + {7'd0,(kernel[4][4] ~^ image[18][26])};
assign out_fmap[14][23][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[14][23])} + {7'd0,(kernel[0][1] ~^ image[14][24])} + {7'd0,(kernel[0][2] ~^ image[14][25])} + {7'd0,(kernel[0][3] ~^ image[14][26])} + {7'd0,(kernel[0][4] ~^ image[14][27])} + {7'd0,(kernel[1][0] ~^ image[15][23])} + {7'd0,(kernel[1][1] ~^ image[15][24])} + {7'd0,(kernel[1][2] ~^ image[15][25])} + {7'd0,(kernel[1][3] ~^ image[15][26])} + {7'd0,(kernel[1][4] ~^ image[15][27])} + {7'd0,(kernel[2][0] ~^ image[16][23])} + {7'd0,(kernel[2][1] ~^ image[16][24])} + {7'd0,(kernel[2][2] ~^ image[16][25])} + {7'd0,(kernel[2][3] ~^ image[16][26])} + {7'd0,(kernel[2][4] ~^ image[16][27])} + {7'd0,(kernel[3][0] ~^ image[17][23])} + {7'd0,(kernel[3][1] ~^ image[17][24])} + {7'd0,(kernel[3][2] ~^ image[17][25])} + {7'd0,(kernel[3][3] ~^ image[17][26])} + {7'd0,(kernel[3][4] ~^ image[17][27])} + {7'd0,(kernel[4][0] ~^ image[18][23])} + {7'd0,(kernel[4][1] ~^ image[18][24])} + {7'd0,(kernel[4][2] ~^ image[18][25])} + {7'd0,(kernel[4][3] ~^ image[18][26])} + {7'd0,(kernel[4][4] ~^ image[18][27])};
assign out_fmap[15][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[15][0])} + {7'd0,(kernel[0][1] ~^ image[15][1])} + {7'd0,(kernel[0][2] ~^ image[15][2])} + {7'd0,(kernel[0][3] ~^ image[15][3])} + {7'd0,(kernel[0][4] ~^ image[15][4])} + {7'd0,(kernel[1][0] ~^ image[16][0])} + {7'd0,(kernel[1][1] ~^ image[16][1])} + {7'd0,(kernel[1][2] ~^ image[16][2])} + {7'd0,(kernel[1][3] ~^ image[16][3])} + {7'd0,(kernel[1][4] ~^ image[16][4])} + {7'd0,(kernel[2][0] ~^ image[17][0])} + {7'd0,(kernel[2][1] ~^ image[17][1])} + {7'd0,(kernel[2][2] ~^ image[17][2])} + {7'd0,(kernel[2][3] ~^ image[17][3])} + {7'd0,(kernel[2][4] ~^ image[17][4])} + {7'd0,(kernel[3][0] ~^ image[18][0])} + {7'd0,(kernel[3][1] ~^ image[18][1])} + {7'd0,(kernel[3][2] ~^ image[18][2])} + {7'd0,(kernel[3][3] ~^ image[18][3])} + {7'd0,(kernel[3][4] ~^ image[18][4])} + {7'd0,(kernel[4][0] ~^ image[19][0])} + {7'd0,(kernel[4][1] ~^ image[19][1])} + {7'd0,(kernel[4][2] ~^ image[19][2])} + {7'd0,(kernel[4][3] ~^ image[19][3])} + {7'd0,(kernel[4][4] ~^ image[19][4])};
assign out_fmap[15][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[15][1])} + {7'd0,(kernel[0][1] ~^ image[15][2])} + {7'd0,(kernel[0][2] ~^ image[15][3])} + {7'd0,(kernel[0][3] ~^ image[15][4])} + {7'd0,(kernel[0][4] ~^ image[15][5])} + {7'd0,(kernel[1][0] ~^ image[16][1])} + {7'd0,(kernel[1][1] ~^ image[16][2])} + {7'd0,(kernel[1][2] ~^ image[16][3])} + {7'd0,(kernel[1][3] ~^ image[16][4])} + {7'd0,(kernel[1][4] ~^ image[16][5])} + {7'd0,(kernel[2][0] ~^ image[17][1])} + {7'd0,(kernel[2][1] ~^ image[17][2])} + {7'd0,(kernel[2][2] ~^ image[17][3])} + {7'd0,(kernel[2][3] ~^ image[17][4])} + {7'd0,(kernel[2][4] ~^ image[17][5])} + {7'd0,(kernel[3][0] ~^ image[18][1])} + {7'd0,(kernel[3][1] ~^ image[18][2])} + {7'd0,(kernel[3][2] ~^ image[18][3])} + {7'd0,(kernel[3][3] ~^ image[18][4])} + {7'd0,(kernel[3][4] ~^ image[18][5])} + {7'd0,(kernel[4][0] ~^ image[19][1])} + {7'd0,(kernel[4][1] ~^ image[19][2])} + {7'd0,(kernel[4][2] ~^ image[19][3])} + {7'd0,(kernel[4][3] ~^ image[19][4])} + {7'd0,(kernel[4][4] ~^ image[19][5])};
assign out_fmap[15][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[15][2])} + {7'd0,(kernel[0][1] ~^ image[15][3])} + {7'd0,(kernel[0][2] ~^ image[15][4])} + {7'd0,(kernel[0][3] ~^ image[15][5])} + {7'd0,(kernel[0][4] ~^ image[15][6])} + {7'd0,(kernel[1][0] ~^ image[16][2])} + {7'd0,(kernel[1][1] ~^ image[16][3])} + {7'd0,(kernel[1][2] ~^ image[16][4])} + {7'd0,(kernel[1][3] ~^ image[16][5])} + {7'd0,(kernel[1][4] ~^ image[16][6])} + {7'd0,(kernel[2][0] ~^ image[17][2])} + {7'd0,(kernel[2][1] ~^ image[17][3])} + {7'd0,(kernel[2][2] ~^ image[17][4])} + {7'd0,(kernel[2][3] ~^ image[17][5])} + {7'd0,(kernel[2][4] ~^ image[17][6])} + {7'd0,(kernel[3][0] ~^ image[18][2])} + {7'd0,(kernel[3][1] ~^ image[18][3])} + {7'd0,(kernel[3][2] ~^ image[18][4])} + {7'd0,(kernel[3][3] ~^ image[18][5])} + {7'd0,(kernel[3][4] ~^ image[18][6])} + {7'd0,(kernel[4][0] ~^ image[19][2])} + {7'd0,(kernel[4][1] ~^ image[19][3])} + {7'd0,(kernel[4][2] ~^ image[19][4])} + {7'd0,(kernel[4][3] ~^ image[19][5])} + {7'd0,(kernel[4][4] ~^ image[19][6])};
assign out_fmap[15][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[15][3])} + {7'd0,(kernel[0][1] ~^ image[15][4])} + {7'd0,(kernel[0][2] ~^ image[15][5])} + {7'd0,(kernel[0][3] ~^ image[15][6])} + {7'd0,(kernel[0][4] ~^ image[15][7])} + {7'd0,(kernel[1][0] ~^ image[16][3])} + {7'd0,(kernel[1][1] ~^ image[16][4])} + {7'd0,(kernel[1][2] ~^ image[16][5])} + {7'd0,(kernel[1][3] ~^ image[16][6])} + {7'd0,(kernel[1][4] ~^ image[16][7])} + {7'd0,(kernel[2][0] ~^ image[17][3])} + {7'd0,(kernel[2][1] ~^ image[17][4])} + {7'd0,(kernel[2][2] ~^ image[17][5])} + {7'd0,(kernel[2][3] ~^ image[17][6])} + {7'd0,(kernel[2][4] ~^ image[17][7])} + {7'd0,(kernel[3][0] ~^ image[18][3])} + {7'd0,(kernel[3][1] ~^ image[18][4])} + {7'd0,(kernel[3][2] ~^ image[18][5])} + {7'd0,(kernel[3][3] ~^ image[18][6])} + {7'd0,(kernel[3][4] ~^ image[18][7])} + {7'd0,(kernel[4][0] ~^ image[19][3])} + {7'd0,(kernel[4][1] ~^ image[19][4])} + {7'd0,(kernel[4][2] ~^ image[19][5])} + {7'd0,(kernel[4][3] ~^ image[19][6])} + {7'd0,(kernel[4][4] ~^ image[19][7])};
assign out_fmap[15][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[15][4])} + {7'd0,(kernel[0][1] ~^ image[15][5])} + {7'd0,(kernel[0][2] ~^ image[15][6])} + {7'd0,(kernel[0][3] ~^ image[15][7])} + {7'd0,(kernel[0][4] ~^ image[15][8])} + {7'd0,(kernel[1][0] ~^ image[16][4])} + {7'd0,(kernel[1][1] ~^ image[16][5])} + {7'd0,(kernel[1][2] ~^ image[16][6])} + {7'd0,(kernel[1][3] ~^ image[16][7])} + {7'd0,(kernel[1][4] ~^ image[16][8])} + {7'd0,(kernel[2][0] ~^ image[17][4])} + {7'd0,(kernel[2][1] ~^ image[17][5])} + {7'd0,(kernel[2][2] ~^ image[17][6])} + {7'd0,(kernel[2][3] ~^ image[17][7])} + {7'd0,(kernel[2][4] ~^ image[17][8])} + {7'd0,(kernel[3][0] ~^ image[18][4])} + {7'd0,(kernel[3][1] ~^ image[18][5])} + {7'd0,(kernel[3][2] ~^ image[18][6])} + {7'd0,(kernel[3][3] ~^ image[18][7])} + {7'd0,(kernel[3][4] ~^ image[18][8])} + {7'd0,(kernel[4][0] ~^ image[19][4])} + {7'd0,(kernel[4][1] ~^ image[19][5])} + {7'd0,(kernel[4][2] ~^ image[19][6])} + {7'd0,(kernel[4][3] ~^ image[19][7])} + {7'd0,(kernel[4][4] ~^ image[19][8])};
assign out_fmap[15][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[15][5])} + {7'd0,(kernel[0][1] ~^ image[15][6])} + {7'd0,(kernel[0][2] ~^ image[15][7])} + {7'd0,(kernel[0][3] ~^ image[15][8])} + {7'd0,(kernel[0][4] ~^ image[15][9])} + {7'd0,(kernel[1][0] ~^ image[16][5])} + {7'd0,(kernel[1][1] ~^ image[16][6])} + {7'd0,(kernel[1][2] ~^ image[16][7])} + {7'd0,(kernel[1][3] ~^ image[16][8])} + {7'd0,(kernel[1][4] ~^ image[16][9])} + {7'd0,(kernel[2][0] ~^ image[17][5])} + {7'd0,(kernel[2][1] ~^ image[17][6])} + {7'd0,(kernel[2][2] ~^ image[17][7])} + {7'd0,(kernel[2][3] ~^ image[17][8])} + {7'd0,(kernel[2][4] ~^ image[17][9])} + {7'd0,(kernel[3][0] ~^ image[18][5])} + {7'd0,(kernel[3][1] ~^ image[18][6])} + {7'd0,(kernel[3][2] ~^ image[18][7])} + {7'd0,(kernel[3][3] ~^ image[18][8])} + {7'd0,(kernel[3][4] ~^ image[18][9])} + {7'd0,(kernel[4][0] ~^ image[19][5])} + {7'd0,(kernel[4][1] ~^ image[19][6])} + {7'd0,(kernel[4][2] ~^ image[19][7])} + {7'd0,(kernel[4][3] ~^ image[19][8])} + {7'd0,(kernel[4][4] ~^ image[19][9])};
assign out_fmap[15][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[15][6])} + {7'd0,(kernel[0][1] ~^ image[15][7])} + {7'd0,(kernel[0][2] ~^ image[15][8])} + {7'd0,(kernel[0][3] ~^ image[15][9])} + {7'd0,(kernel[0][4] ~^ image[15][10])} + {7'd0,(kernel[1][0] ~^ image[16][6])} + {7'd0,(kernel[1][1] ~^ image[16][7])} + {7'd0,(kernel[1][2] ~^ image[16][8])} + {7'd0,(kernel[1][3] ~^ image[16][9])} + {7'd0,(kernel[1][4] ~^ image[16][10])} + {7'd0,(kernel[2][0] ~^ image[17][6])} + {7'd0,(kernel[2][1] ~^ image[17][7])} + {7'd0,(kernel[2][2] ~^ image[17][8])} + {7'd0,(kernel[2][3] ~^ image[17][9])} + {7'd0,(kernel[2][4] ~^ image[17][10])} + {7'd0,(kernel[3][0] ~^ image[18][6])} + {7'd0,(kernel[3][1] ~^ image[18][7])} + {7'd0,(kernel[3][2] ~^ image[18][8])} + {7'd0,(kernel[3][3] ~^ image[18][9])} + {7'd0,(kernel[3][4] ~^ image[18][10])} + {7'd0,(kernel[4][0] ~^ image[19][6])} + {7'd0,(kernel[4][1] ~^ image[19][7])} + {7'd0,(kernel[4][2] ~^ image[19][8])} + {7'd0,(kernel[4][3] ~^ image[19][9])} + {7'd0,(kernel[4][4] ~^ image[19][10])};
assign out_fmap[15][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[15][7])} + {7'd0,(kernel[0][1] ~^ image[15][8])} + {7'd0,(kernel[0][2] ~^ image[15][9])} + {7'd0,(kernel[0][3] ~^ image[15][10])} + {7'd0,(kernel[0][4] ~^ image[15][11])} + {7'd0,(kernel[1][0] ~^ image[16][7])} + {7'd0,(kernel[1][1] ~^ image[16][8])} + {7'd0,(kernel[1][2] ~^ image[16][9])} + {7'd0,(kernel[1][3] ~^ image[16][10])} + {7'd0,(kernel[1][4] ~^ image[16][11])} + {7'd0,(kernel[2][0] ~^ image[17][7])} + {7'd0,(kernel[2][1] ~^ image[17][8])} + {7'd0,(kernel[2][2] ~^ image[17][9])} + {7'd0,(kernel[2][3] ~^ image[17][10])} + {7'd0,(kernel[2][4] ~^ image[17][11])} + {7'd0,(kernel[3][0] ~^ image[18][7])} + {7'd0,(kernel[3][1] ~^ image[18][8])} + {7'd0,(kernel[3][2] ~^ image[18][9])} + {7'd0,(kernel[3][3] ~^ image[18][10])} + {7'd0,(kernel[3][4] ~^ image[18][11])} + {7'd0,(kernel[4][0] ~^ image[19][7])} + {7'd0,(kernel[4][1] ~^ image[19][8])} + {7'd0,(kernel[4][2] ~^ image[19][9])} + {7'd0,(kernel[4][3] ~^ image[19][10])} + {7'd0,(kernel[4][4] ~^ image[19][11])};
assign out_fmap[15][8][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[15][8])} + {7'd0,(kernel[0][1] ~^ image[15][9])} + {7'd0,(kernel[0][2] ~^ image[15][10])} + {7'd0,(kernel[0][3] ~^ image[15][11])} + {7'd0,(kernel[0][4] ~^ image[15][12])} + {7'd0,(kernel[1][0] ~^ image[16][8])} + {7'd0,(kernel[1][1] ~^ image[16][9])} + {7'd0,(kernel[1][2] ~^ image[16][10])} + {7'd0,(kernel[1][3] ~^ image[16][11])} + {7'd0,(kernel[1][4] ~^ image[16][12])} + {7'd0,(kernel[2][0] ~^ image[17][8])} + {7'd0,(kernel[2][1] ~^ image[17][9])} + {7'd0,(kernel[2][2] ~^ image[17][10])} + {7'd0,(kernel[2][3] ~^ image[17][11])} + {7'd0,(kernel[2][4] ~^ image[17][12])} + {7'd0,(kernel[3][0] ~^ image[18][8])} + {7'd0,(kernel[3][1] ~^ image[18][9])} + {7'd0,(kernel[3][2] ~^ image[18][10])} + {7'd0,(kernel[3][3] ~^ image[18][11])} + {7'd0,(kernel[3][4] ~^ image[18][12])} + {7'd0,(kernel[4][0] ~^ image[19][8])} + {7'd0,(kernel[4][1] ~^ image[19][9])} + {7'd0,(kernel[4][2] ~^ image[19][10])} + {7'd0,(kernel[4][3] ~^ image[19][11])} + {7'd0,(kernel[4][4] ~^ image[19][12])};
assign out_fmap[15][9][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[15][9])} + {7'd0,(kernel[0][1] ~^ image[15][10])} + {7'd0,(kernel[0][2] ~^ image[15][11])} + {7'd0,(kernel[0][3] ~^ image[15][12])} + {7'd0,(kernel[0][4] ~^ image[15][13])} + {7'd0,(kernel[1][0] ~^ image[16][9])} + {7'd0,(kernel[1][1] ~^ image[16][10])} + {7'd0,(kernel[1][2] ~^ image[16][11])} + {7'd0,(kernel[1][3] ~^ image[16][12])} + {7'd0,(kernel[1][4] ~^ image[16][13])} + {7'd0,(kernel[2][0] ~^ image[17][9])} + {7'd0,(kernel[2][1] ~^ image[17][10])} + {7'd0,(kernel[2][2] ~^ image[17][11])} + {7'd0,(kernel[2][3] ~^ image[17][12])} + {7'd0,(kernel[2][4] ~^ image[17][13])} + {7'd0,(kernel[3][0] ~^ image[18][9])} + {7'd0,(kernel[3][1] ~^ image[18][10])} + {7'd0,(kernel[3][2] ~^ image[18][11])} + {7'd0,(kernel[3][3] ~^ image[18][12])} + {7'd0,(kernel[3][4] ~^ image[18][13])} + {7'd0,(kernel[4][0] ~^ image[19][9])} + {7'd0,(kernel[4][1] ~^ image[19][10])} + {7'd0,(kernel[4][2] ~^ image[19][11])} + {7'd0,(kernel[4][3] ~^ image[19][12])} + {7'd0,(kernel[4][4] ~^ image[19][13])};
assign out_fmap[15][10][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[15][10])} + {7'd0,(kernel[0][1] ~^ image[15][11])} + {7'd0,(kernel[0][2] ~^ image[15][12])} + {7'd0,(kernel[0][3] ~^ image[15][13])} + {7'd0,(kernel[0][4] ~^ image[15][14])} + {7'd0,(kernel[1][0] ~^ image[16][10])} + {7'd0,(kernel[1][1] ~^ image[16][11])} + {7'd0,(kernel[1][2] ~^ image[16][12])} + {7'd0,(kernel[1][3] ~^ image[16][13])} + {7'd0,(kernel[1][4] ~^ image[16][14])} + {7'd0,(kernel[2][0] ~^ image[17][10])} + {7'd0,(kernel[2][1] ~^ image[17][11])} + {7'd0,(kernel[2][2] ~^ image[17][12])} + {7'd0,(kernel[2][3] ~^ image[17][13])} + {7'd0,(kernel[2][4] ~^ image[17][14])} + {7'd0,(kernel[3][0] ~^ image[18][10])} + {7'd0,(kernel[3][1] ~^ image[18][11])} + {7'd0,(kernel[3][2] ~^ image[18][12])} + {7'd0,(kernel[3][3] ~^ image[18][13])} + {7'd0,(kernel[3][4] ~^ image[18][14])} + {7'd0,(kernel[4][0] ~^ image[19][10])} + {7'd0,(kernel[4][1] ~^ image[19][11])} + {7'd0,(kernel[4][2] ~^ image[19][12])} + {7'd0,(kernel[4][3] ~^ image[19][13])} + {7'd0,(kernel[4][4] ~^ image[19][14])};
assign out_fmap[15][11][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[15][11])} + {7'd0,(kernel[0][1] ~^ image[15][12])} + {7'd0,(kernel[0][2] ~^ image[15][13])} + {7'd0,(kernel[0][3] ~^ image[15][14])} + {7'd0,(kernel[0][4] ~^ image[15][15])} + {7'd0,(kernel[1][0] ~^ image[16][11])} + {7'd0,(kernel[1][1] ~^ image[16][12])} + {7'd0,(kernel[1][2] ~^ image[16][13])} + {7'd0,(kernel[1][3] ~^ image[16][14])} + {7'd0,(kernel[1][4] ~^ image[16][15])} + {7'd0,(kernel[2][0] ~^ image[17][11])} + {7'd0,(kernel[2][1] ~^ image[17][12])} + {7'd0,(kernel[2][2] ~^ image[17][13])} + {7'd0,(kernel[2][3] ~^ image[17][14])} + {7'd0,(kernel[2][4] ~^ image[17][15])} + {7'd0,(kernel[3][0] ~^ image[18][11])} + {7'd0,(kernel[3][1] ~^ image[18][12])} + {7'd0,(kernel[3][2] ~^ image[18][13])} + {7'd0,(kernel[3][3] ~^ image[18][14])} + {7'd0,(kernel[3][4] ~^ image[18][15])} + {7'd0,(kernel[4][0] ~^ image[19][11])} + {7'd0,(kernel[4][1] ~^ image[19][12])} + {7'd0,(kernel[4][2] ~^ image[19][13])} + {7'd0,(kernel[4][3] ~^ image[19][14])} + {7'd0,(kernel[4][4] ~^ image[19][15])};
assign out_fmap[15][12][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[15][12])} + {7'd0,(kernel[0][1] ~^ image[15][13])} + {7'd0,(kernel[0][2] ~^ image[15][14])} + {7'd0,(kernel[0][3] ~^ image[15][15])} + {7'd0,(kernel[0][4] ~^ image[15][16])} + {7'd0,(kernel[1][0] ~^ image[16][12])} + {7'd0,(kernel[1][1] ~^ image[16][13])} + {7'd0,(kernel[1][2] ~^ image[16][14])} + {7'd0,(kernel[1][3] ~^ image[16][15])} + {7'd0,(kernel[1][4] ~^ image[16][16])} + {7'd0,(kernel[2][0] ~^ image[17][12])} + {7'd0,(kernel[2][1] ~^ image[17][13])} + {7'd0,(kernel[2][2] ~^ image[17][14])} + {7'd0,(kernel[2][3] ~^ image[17][15])} + {7'd0,(kernel[2][4] ~^ image[17][16])} + {7'd0,(kernel[3][0] ~^ image[18][12])} + {7'd0,(kernel[3][1] ~^ image[18][13])} + {7'd0,(kernel[3][2] ~^ image[18][14])} + {7'd0,(kernel[3][3] ~^ image[18][15])} + {7'd0,(kernel[3][4] ~^ image[18][16])} + {7'd0,(kernel[4][0] ~^ image[19][12])} + {7'd0,(kernel[4][1] ~^ image[19][13])} + {7'd0,(kernel[4][2] ~^ image[19][14])} + {7'd0,(kernel[4][3] ~^ image[19][15])} + {7'd0,(kernel[4][4] ~^ image[19][16])};
assign out_fmap[15][13][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[15][13])} + {7'd0,(kernel[0][1] ~^ image[15][14])} + {7'd0,(kernel[0][2] ~^ image[15][15])} + {7'd0,(kernel[0][3] ~^ image[15][16])} + {7'd0,(kernel[0][4] ~^ image[15][17])} + {7'd0,(kernel[1][0] ~^ image[16][13])} + {7'd0,(kernel[1][1] ~^ image[16][14])} + {7'd0,(kernel[1][2] ~^ image[16][15])} + {7'd0,(kernel[1][3] ~^ image[16][16])} + {7'd0,(kernel[1][4] ~^ image[16][17])} + {7'd0,(kernel[2][0] ~^ image[17][13])} + {7'd0,(kernel[2][1] ~^ image[17][14])} + {7'd0,(kernel[2][2] ~^ image[17][15])} + {7'd0,(kernel[2][3] ~^ image[17][16])} + {7'd0,(kernel[2][4] ~^ image[17][17])} + {7'd0,(kernel[3][0] ~^ image[18][13])} + {7'd0,(kernel[3][1] ~^ image[18][14])} + {7'd0,(kernel[3][2] ~^ image[18][15])} + {7'd0,(kernel[3][3] ~^ image[18][16])} + {7'd0,(kernel[3][4] ~^ image[18][17])} + {7'd0,(kernel[4][0] ~^ image[19][13])} + {7'd0,(kernel[4][1] ~^ image[19][14])} + {7'd0,(kernel[4][2] ~^ image[19][15])} + {7'd0,(kernel[4][3] ~^ image[19][16])} + {7'd0,(kernel[4][4] ~^ image[19][17])};
assign out_fmap[15][14][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[15][14])} + {7'd0,(kernel[0][1] ~^ image[15][15])} + {7'd0,(kernel[0][2] ~^ image[15][16])} + {7'd0,(kernel[0][3] ~^ image[15][17])} + {7'd0,(kernel[0][4] ~^ image[15][18])} + {7'd0,(kernel[1][0] ~^ image[16][14])} + {7'd0,(kernel[1][1] ~^ image[16][15])} + {7'd0,(kernel[1][2] ~^ image[16][16])} + {7'd0,(kernel[1][3] ~^ image[16][17])} + {7'd0,(kernel[1][4] ~^ image[16][18])} + {7'd0,(kernel[2][0] ~^ image[17][14])} + {7'd0,(kernel[2][1] ~^ image[17][15])} + {7'd0,(kernel[2][2] ~^ image[17][16])} + {7'd0,(kernel[2][3] ~^ image[17][17])} + {7'd0,(kernel[2][4] ~^ image[17][18])} + {7'd0,(kernel[3][0] ~^ image[18][14])} + {7'd0,(kernel[3][1] ~^ image[18][15])} + {7'd0,(kernel[3][2] ~^ image[18][16])} + {7'd0,(kernel[3][3] ~^ image[18][17])} + {7'd0,(kernel[3][4] ~^ image[18][18])} + {7'd0,(kernel[4][0] ~^ image[19][14])} + {7'd0,(kernel[4][1] ~^ image[19][15])} + {7'd0,(kernel[4][2] ~^ image[19][16])} + {7'd0,(kernel[4][3] ~^ image[19][17])} + {7'd0,(kernel[4][4] ~^ image[19][18])};
assign out_fmap[15][15][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[15][15])} + {7'd0,(kernel[0][1] ~^ image[15][16])} + {7'd0,(kernel[0][2] ~^ image[15][17])} + {7'd0,(kernel[0][3] ~^ image[15][18])} + {7'd0,(kernel[0][4] ~^ image[15][19])} + {7'd0,(kernel[1][0] ~^ image[16][15])} + {7'd0,(kernel[1][1] ~^ image[16][16])} + {7'd0,(kernel[1][2] ~^ image[16][17])} + {7'd0,(kernel[1][3] ~^ image[16][18])} + {7'd0,(kernel[1][4] ~^ image[16][19])} + {7'd0,(kernel[2][0] ~^ image[17][15])} + {7'd0,(kernel[2][1] ~^ image[17][16])} + {7'd0,(kernel[2][2] ~^ image[17][17])} + {7'd0,(kernel[2][3] ~^ image[17][18])} + {7'd0,(kernel[2][4] ~^ image[17][19])} + {7'd0,(kernel[3][0] ~^ image[18][15])} + {7'd0,(kernel[3][1] ~^ image[18][16])} + {7'd0,(kernel[3][2] ~^ image[18][17])} + {7'd0,(kernel[3][3] ~^ image[18][18])} + {7'd0,(kernel[3][4] ~^ image[18][19])} + {7'd0,(kernel[4][0] ~^ image[19][15])} + {7'd0,(kernel[4][1] ~^ image[19][16])} + {7'd0,(kernel[4][2] ~^ image[19][17])} + {7'd0,(kernel[4][3] ~^ image[19][18])} + {7'd0,(kernel[4][4] ~^ image[19][19])};
assign out_fmap[15][16][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[15][16])} + {7'd0,(kernel[0][1] ~^ image[15][17])} + {7'd0,(kernel[0][2] ~^ image[15][18])} + {7'd0,(kernel[0][3] ~^ image[15][19])} + {7'd0,(kernel[0][4] ~^ image[15][20])} + {7'd0,(kernel[1][0] ~^ image[16][16])} + {7'd0,(kernel[1][1] ~^ image[16][17])} + {7'd0,(kernel[1][2] ~^ image[16][18])} + {7'd0,(kernel[1][3] ~^ image[16][19])} + {7'd0,(kernel[1][4] ~^ image[16][20])} + {7'd0,(kernel[2][0] ~^ image[17][16])} + {7'd0,(kernel[2][1] ~^ image[17][17])} + {7'd0,(kernel[2][2] ~^ image[17][18])} + {7'd0,(kernel[2][3] ~^ image[17][19])} + {7'd0,(kernel[2][4] ~^ image[17][20])} + {7'd0,(kernel[3][0] ~^ image[18][16])} + {7'd0,(kernel[3][1] ~^ image[18][17])} + {7'd0,(kernel[3][2] ~^ image[18][18])} + {7'd0,(kernel[3][3] ~^ image[18][19])} + {7'd0,(kernel[3][4] ~^ image[18][20])} + {7'd0,(kernel[4][0] ~^ image[19][16])} + {7'd0,(kernel[4][1] ~^ image[19][17])} + {7'd0,(kernel[4][2] ~^ image[19][18])} + {7'd0,(kernel[4][3] ~^ image[19][19])} + {7'd0,(kernel[4][4] ~^ image[19][20])};
assign out_fmap[15][17][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[15][17])} + {7'd0,(kernel[0][1] ~^ image[15][18])} + {7'd0,(kernel[0][2] ~^ image[15][19])} + {7'd0,(kernel[0][3] ~^ image[15][20])} + {7'd0,(kernel[0][4] ~^ image[15][21])} + {7'd0,(kernel[1][0] ~^ image[16][17])} + {7'd0,(kernel[1][1] ~^ image[16][18])} + {7'd0,(kernel[1][2] ~^ image[16][19])} + {7'd0,(kernel[1][3] ~^ image[16][20])} + {7'd0,(kernel[1][4] ~^ image[16][21])} + {7'd0,(kernel[2][0] ~^ image[17][17])} + {7'd0,(kernel[2][1] ~^ image[17][18])} + {7'd0,(kernel[2][2] ~^ image[17][19])} + {7'd0,(kernel[2][3] ~^ image[17][20])} + {7'd0,(kernel[2][4] ~^ image[17][21])} + {7'd0,(kernel[3][0] ~^ image[18][17])} + {7'd0,(kernel[3][1] ~^ image[18][18])} + {7'd0,(kernel[3][2] ~^ image[18][19])} + {7'd0,(kernel[3][3] ~^ image[18][20])} + {7'd0,(kernel[3][4] ~^ image[18][21])} + {7'd0,(kernel[4][0] ~^ image[19][17])} + {7'd0,(kernel[4][1] ~^ image[19][18])} + {7'd0,(kernel[4][2] ~^ image[19][19])} + {7'd0,(kernel[4][3] ~^ image[19][20])} + {7'd0,(kernel[4][4] ~^ image[19][21])};
assign out_fmap[15][18][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[15][18])} + {7'd0,(kernel[0][1] ~^ image[15][19])} + {7'd0,(kernel[0][2] ~^ image[15][20])} + {7'd0,(kernel[0][3] ~^ image[15][21])} + {7'd0,(kernel[0][4] ~^ image[15][22])} + {7'd0,(kernel[1][0] ~^ image[16][18])} + {7'd0,(kernel[1][1] ~^ image[16][19])} + {7'd0,(kernel[1][2] ~^ image[16][20])} + {7'd0,(kernel[1][3] ~^ image[16][21])} + {7'd0,(kernel[1][4] ~^ image[16][22])} + {7'd0,(kernel[2][0] ~^ image[17][18])} + {7'd0,(kernel[2][1] ~^ image[17][19])} + {7'd0,(kernel[2][2] ~^ image[17][20])} + {7'd0,(kernel[2][3] ~^ image[17][21])} + {7'd0,(kernel[2][4] ~^ image[17][22])} + {7'd0,(kernel[3][0] ~^ image[18][18])} + {7'd0,(kernel[3][1] ~^ image[18][19])} + {7'd0,(kernel[3][2] ~^ image[18][20])} + {7'd0,(kernel[3][3] ~^ image[18][21])} + {7'd0,(kernel[3][4] ~^ image[18][22])} + {7'd0,(kernel[4][0] ~^ image[19][18])} + {7'd0,(kernel[4][1] ~^ image[19][19])} + {7'd0,(kernel[4][2] ~^ image[19][20])} + {7'd0,(kernel[4][3] ~^ image[19][21])} + {7'd0,(kernel[4][4] ~^ image[19][22])};
assign out_fmap[15][19][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[15][19])} + {7'd0,(kernel[0][1] ~^ image[15][20])} + {7'd0,(kernel[0][2] ~^ image[15][21])} + {7'd0,(kernel[0][3] ~^ image[15][22])} + {7'd0,(kernel[0][4] ~^ image[15][23])} + {7'd0,(kernel[1][0] ~^ image[16][19])} + {7'd0,(kernel[1][1] ~^ image[16][20])} + {7'd0,(kernel[1][2] ~^ image[16][21])} + {7'd0,(kernel[1][3] ~^ image[16][22])} + {7'd0,(kernel[1][4] ~^ image[16][23])} + {7'd0,(kernel[2][0] ~^ image[17][19])} + {7'd0,(kernel[2][1] ~^ image[17][20])} + {7'd0,(kernel[2][2] ~^ image[17][21])} + {7'd0,(kernel[2][3] ~^ image[17][22])} + {7'd0,(kernel[2][4] ~^ image[17][23])} + {7'd0,(kernel[3][0] ~^ image[18][19])} + {7'd0,(kernel[3][1] ~^ image[18][20])} + {7'd0,(kernel[3][2] ~^ image[18][21])} + {7'd0,(kernel[3][3] ~^ image[18][22])} + {7'd0,(kernel[3][4] ~^ image[18][23])} + {7'd0,(kernel[4][0] ~^ image[19][19])} + {7'd0,(kernel[4][1] ~^ image[19][20])} + {7'd0,(kernel[4][2] ~^ image[19][21])} + {7'd0,(kernel[4][3] ~^ image[19][22])} + {7'd0,(kernel[4][4] ~^ image[19][23])};
assign out_fmap[15][20][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[15][20])} + {7'd0,(kernel[0][1] ~^ image[15][21])} + {7'd0,(kernel[0][2] ~^ image[15][22])} + {7'd0,(kernel[0][3] ~^ image[15][23])} + {7'd0,(kernel[0][4] ~^ image[15][24])} + {7'd0,(kernel[1][0] ~^ image[16][20])} + {7'd0,(kernel[1][1] ~^ image[16][21])} + {7'd0,(kernel[1][2] ~^ image[16][22])} + {7'd0,(kernel[1][3] ~^ image[16][23])} + {7'd0,(kernel[1][4] ~^ image[16][24])} + {7'd0,(kernel[2][0] ~^ image[17][20])} + {7'd0,(kernel[2][1] ~^ image[17][21])} + {7'd0,(kernel[2][2] ~^ image[17][22])} + {7'd0,(kernel[2][3] ~^ image[17][23])} + {7'd0,(kernel[2][4] ~^ image[17][24])} + {7'd0,(kernel[3][0] ~^ image[18][20])} + {7'd0,(kernel[3][1] ~^ image[18][21])} + {7'd0,(kernel[3][2] ~^ image[18][22])} + {7'd0,(kernel[3][3] ~^ image[18][23])} + {7'd0,(kernel[3][4] ~^ image[18][24])} + {7'd0,(kernel[4][0] ~^ image[19][20])} + {7'd0,(kernel[4][1] ~^ image[19][21])} + {7'd0,(kernel[4][2] ~^ image[19][22])} + {7'd0,(kernel[4][3] ~^ image[19][23])} + {7'd0,(kernel[4][4] ~^ image[19][24])};
assign out_fmap[15][21][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[15][21])} + {7'd0,(kernel[0][1] ~^ image[15][22])} + {7'd0,(kernel[0][2] ~^ image[15][23])} + {7'd0,(kernel[0][3] ~^ image[15][24])} + {7'd0,(kernel[0][4] ~^ image[15][25])} + {7'd0,(kernel[1][0] ~^ image[16][21])} + {7'd0,(kernel[1][1] ~^ image[16][22])} + {7'd0,(kernel[1][2] ~^ image[16][23])} + {7'd0,(kernel[1][3] ~^ image[16][24])} + {7'd0,(kernel[1][4] ~^ image[16][25])} + {7'd0,(kernel[2][0] ~^ image[17][21])} + {7'd0,(kernel[2][1] ~^ image[17][22])} + {7'd0,(kernel[2][2] ~^ image[17][23])} + {7'd0,(kernel[2][3] ~^ image[17][24])} + {7'd0,(kernel[2][4] ~^ image[17][25])} + {7'd0,(kernel[3][0] ~^ image[18][21])} + {7'd0,(kernel[3][1] ~^ image[18][22])} + {7'd0,(kernel[3][2] ~^ image[18][23])} + {7'd0,(kernel[3][3] ~^ image[18][24])} + {7'd0,(kernel[3][4] ~^ image[18][25])} + {7'd0,(kernel[4][0] ~^ image[19][21])} + {7'd0,(kernel[4][1] ~^ image[19][22])} + {7'd0,(kernel[4][2] ~^ image[19][23])} + {7'd0,(kernel[4][3] ~^ image[19][24])} + {7'd0,(kernel[4][4] ~^ image[19][25])};
assign out_fmap[15][22][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[15][22])} + {7'd0,(kernel[0][1] ~^ image[15][23])} + {7'd0,(kernel[0][2] ~^ image[15][24])} + {7'd0,(kernel[0][3] ~^ image[15][25])} + {7'd0,(kernel[0][4] ~^ image[15][26])} + {7'd0,(kernel[1][0] ~^ image[16][22])} + {7'd0,(kernel[1][1] ~^ image[16][23])} + {7'd0,(kernel[1][2] ~^ image[16][24])} + {7'd0,(kernel[1][3] ~^ image[16][25])} + {7'd0,(kernel[1][4] ~^ image[16][26])} + {7'd0,(kernel[2][0] ~^ image[17][22])} + {7'd0,(kernel[2][1] ~^ image[17][23])} + {7'd0,(kernel[2][2] ~^ image[17][24])} + {7'd0,(kernel[2][3] ~^ image[17][25])} + {7'd0,(kernel[2][4] ~^ image[17][26])} + {7'd0,(kernel[3][0] ~^ image[18][22])} + {7'd0,(kernel[3][1] ~^ image[18][23])} + {7'd0,(kernel[3][2] ~^ image[18][24])} + {7'd0,(kernel[3][3] ~^ image[18][25])} + {7'd0,(kernel[3][4] ~^ image[18][26])} + {7'd0,(kernel[4][0] ~^ image[19][22])} + {7'd0,(kernel[4][1] ~^ image[19][23])} + {7'd0,(kernel[4][2] ~^ image[19][24])} + {7'd0,(kernel[4][3] ~^ image[19][25])} + {7'd0,(kernel[4][4] ~^ image[19][26])};
assign out_fmap[15][23][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[15][23])} + {7'd0,(kernel[0][1] ~^ image[15][24])} + {7'd0,(kernel[0][2] ~^ image[15][25])} + {7'd0,(kernel[0][3] ~^ image[15][26])} + {7'd0,(kernel[0][4] ~^ image[15][27])} + {7'd0,(kernel[1][0] ~^ image[16][23])} + {7'd0,(kernel[1][1] ~^ image[16][24])} + {7'd0,(kernel[1][2] ~^ image[16][25])} + {7'd0,(kernel[1][3] ~^ image[16][26])} + {7'd0,(kernel[1][4] ~^ image[16][27])} + {7'd0,(kernel[2][0] ~^ image[17][23])} + {7'd0,(kernel[2][1] ~^ image[17][24])} + {7'd0,(kernel[2][2] ~^ image[17][25])} + {7'd0,(kernel[2][3] ~^ image[17][26])} + {7'd0,(kernel[2][4] ~^ image[17][27])} + {7'd0,(kernel[3][0] ~^ image[18][23])} + {7'd0,(kernel[3][1] ~^ image[18][24])} + {7'd0,(kernel[3][2] ~^ image[18][25])} + {7'd0,(kernel[3][3] ~^ image[18][26])} + {7'd0,(kernel[3][4] ~^ image[18][27])} + {7'd0,(kernel[4][0] ~^ image[19][23])} + {7'd0,(kernel[4][1] ~^ image[19][24])} + {7'd0,(kernel[4][2] ~^ image[19][25])} + {7'd0,(kernel[4][3] ~^ image[19][26])} + {7'd0,(kernel[4][4] ~^ image[19][27])};
assign out_fmap[16][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[16][0])} + {7'd0,(kernel[0][1] ~^ image[16][1])} + {7'd0,(kernel[0][2] ~^ image[16][2])} + {7'd0,(kernel[0][3] ~^ image[16][3])} + {7'd0,(kernel[0][4] ~^ image[16][4])} + {7'd0,(kernel[1][0] ~^ image[17][0])} + {7'd0,(kernel[1][1] ~^ image[17][1])} + {7'd0,(kernel[1][2] ~^ image[17][2])} + {7'd0,(kernel[1][3] ~^ image[17][3])} + {7'd0,(kernel[1][4] ~^ image[17][4])} + {7'd0,(kernel[2][0] ~^ image[18][0])} + {7'd0,(kernel[2][1] ~^ image[18][1])} + {7'd0,(kernel[2][2] ~^ image[18][2])} + {7'd0,(kernel[2][3] ~^ image[18][3])} + {7'd0,(kernel[2][4] ~^ image[18][4])} + {7'd0,(kernel[3][0] ~^ image[19][0])} + {7'd0,(kernel[3][1] ~^ image[19][1])} + {7'd0,(kernel[3][2] ~^ image[19][2])} + {7'd0,(kernel[3][3] ~^ image[19][3])} + {7'd0,(kernel[3][4] ~^ image[19][4])} + {7'd0,(kernel[4][0] ~^ image[20][0])} + {7'd0,(kernel[4][1] ~^ image[20][1])} + {7'd0,(kernel[4][2] ~^ image[20][2])} + {7'd0,(kernel[4][3] ~^ image[20][3])} + {7'd0,(kernel[4][4] ~^ image[20][4])};
assign out_fmap[16][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[16][1])} + {7'd0,(kernel[0][1] ~^ image[16][2])} + {7'd0,(kernel[0][2] ~^ image[16][3])} + {7'd0,(kernel[0][3] ~^ image[16][4])} + {7'd0,(kernel[0][4] ~^ image[16][5])} + {7'd0,(kernel[1][0] ~^ image[17][1])} + {7'd0,(kernel[1][1] ~^ image[17][2])} + {7'd0,(kernel[1][2] ~^ image[17][3])} + {7'd0,(kernel[1][3] ~^ image[17][4])} + {7'd0,(kernel[1][4] ~^ image[17][5])} + {7'd0,(kernel[2][0] ~^ image[18][1])} + {7'd0,(kernel[2][1] ~^ image[18][2])} + {7'd0,(kernel[2][2] ~^ image[18][3])} + {7'd0,(kernel[2][3] ~^ image[18][4])} + {7'd0,(kernel[2][4] ~^ image[18][5])} + {7'd0,(kernel[3][0] ~^ image[19][1])} + {7'd0,(kernel[3][1] ~^ image[19][2])} + {7'd0,(kernel[3][2] ~^ image[19][3])} + {7'd0,(kernel[3][3] ~^ image[19][4])} + {7'd0,(kernel[3][4] ~^ image[19][5])} + {7'd0,(kernel[4][0] ~^ image[20][1])} + {7'd0,(kernel[4][1] ~^ image[20][2])} + {7'd0,(kernel[4][2] ~^ image[20][3])} + {7'd0,(kernel[4][3] ~^ image[20][4])} + {7'd0,(kernel[4][4] ~^ image[20][5])};
assign out_fmap[16][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[16][2])} + {7'd0,(kernel[0][1] ~^ image[16][3])} + {7'd0,(kernel[0][2] ~^ image[16][4])} + {7'd0,(kernel[0][3] ~^ image[16][5])} + {7'd0,(kernel[0][4] ~^ image[16][6])} + {7'd0,(kernel[1][0] ~^ image[17][2])} + {7'd0,(kernel[1][1] ~^ image[17][3])} + {7'd0,(kernel[1][2] ~^ image[17][4])} + {7'd0,(kernel[1][3] ~^ image[17][5])} + {7'd0,(kernel[1][4] ~^ image[17][6])} + {7'd0,(kernel[2][0] ~^ image[18][2])} + {7'd0,(kernel[2][1] ~^ image[18][3])} + {7'd0,(kernel[2][2] ~^ image[18][4])} + {7'd0,(kernel[2][3] ~^ image[18][5])} + {7'd0,(kernel[2][4] ~^ image[18][6])} + {7'd0,(kernel[3][0] ~^ image[19][2])} + {7'd0,(kernel[3][1] ~^ image[19][3])} + {7'd0,(kernel[3][2] ~^ image[19][4])} + {7'd0,(kernel[3][3] ~^ image[19][5])} + {7'd0,(kernel[3][4] ~^ image[19][6])} + {7'd0,(kernel[4][0] ~^ image[20][2])} + {7'd0,(kernel[4][1] ~^ image[20][3])} + {7'd0,(kernel[4][2] ~^ image[20][4])} + {7'd0,(kernel[4][3] ~^ image[20][5])} + {7'd0,(kernel[4][4] ~^ image[20][6])};
assign out_fmap[16][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[16][3])} + {7'd0,(kernel[0][1] ~^ image[16][4])} + {7'd0,(kernel[0][2] ~^ image[16][5])} + {7'd0,(kernel[0][3] ~^ image[16][6])} + {7'd0,(kernel[0][4] ~^ image[16][7])} + {7'd0,(kernel[1][0] ~^ image[17][3])} + {7'd0,(kernel[1][1] ~^ image[17][4])} + {7'd0,(kernel[1][2] ~^ image[17][5])} + {7'd0,(kernel[1][3] ~^ image[17][6])} + {7'd0,(kernel[1][4] ~^ image[17][7])} + {7'd0,(kernel[2][0] ~^ image[18][3])} + {7'd0,(kernel[2][1] ~^ image[18][4])} + {7'd0,(kernel[2][2] ~^ image[18][5])} + {7'd0,(kernel[2][3] ~^ image[18][6])} + {7'd0,(kernel[2][4] ~^ image[18][7])} + {7'd0,(kernel[3][0] ~^ image[19][3])} + {7'd0,(kernel[3][1] ~^ image[19][4])} + {7'd0,(kernel[3][2] ~^ image[19][5])} + {7'd0,(kernel[3][3] ~^ image[19][6])} + {7'd0,(kernel[3][4] ~^ image[19][7])} + {7'd0,(kernel[4][0] ~^ image[20][3])} + {7'd0,(kernel[4][1] ~^ image[20][4])} + {7'd0,(kernel[4][2] ~^ image[20][5])} + {7'd0,(kernel[4][3] ~^ image[20][6])} + {7'd0,(kernel[4][4] ~^ image[20][7])};
assign out_fmap[16][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[16][4])} + {7'd0,(kernel[0][1] ~^ image[16][5])} + {7'd0,(kernel[0][2] ~^ image[16][6])} + {7'd0,(kernel[0][3] ~^ image[16][7])} + {7'd0,(kernel[0][4] ~^ image[16][8])} + {7'd0,(kernel[1][0] ~^ image[17][4])} + {7'd0,(kernel[1][1] ~^ image[17][5])} + {7'd0,(kernel[1][2] ~^ image[17][6])} + {7'd0,(kernel[1][3] ~^ image[17][7])} + {7'd0,(kernel[1][4] ~^ image[17][8])} + {7'd0,(kernel[2][0] ~^ image[18][4])} + {7'd0,(kernel[2][1] ~^ image[18][5])} + {7'd0,(kernel[2][2] ~^ image[18][6])} + {7'd0,(kernel[2][3] ~^ image[18][7])} + {7'd0,(kernel[2][4] ~^ image[18][8])} + {7'd0,(kernel[3][0] ~^ image[19][4])} + {7'd0,(kernel[3][1] ~^ image[19][5])} + {7'd0,(kernel[3][2] ~^ image[19][6])} + {7'd0,(kernel[3][3] ~^ image[19][7])} + {7'd0,(kernel[3][4] ~^ image[19][8])} + {7'd0,(kernel[4][0] ~^ image[20][4])} + {7'd0,(kernel[4][1] ~^ image[20][5])} + {7'd0,(kernel[4][2] ~^ image[20][6])} + {7'd0,(kernel[4][3] ~^ image[20][7])} + {7'd0,(kernel[4][4] ~^ image[20][8])};
assign out_fmap[16][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[16][5])} + {7'd0,(kernel[0][1] ~^ image[16][6])} + {7'd0,(kernel[0][2] ~^ image[16][7])} + {7'd0,(kernel[0][3] ~^ image[16][8])} + {7'd0,(kernel[0][4] ~^ image[16][9])} + {7'd0,(kernel[1][0] ~^ image[17][5])} + {7'd0,(kernel[1][1] ~^ image[17][6])} + {7'd0,(kernel[1][2] ~^ image[17][7])} + {7'd0,(kernel[1][3] ~^ image[17][8])} + {7'd0,(kernel[1][4] ~^ image[17][9])} + {7'd0,(kernel[2][0] ~^ image[18][5])} + {7'd0,(kernel[2][1] ~^ image[18][6])} + {7'd0,(kernel[2][2] ~^ image[18][7])} + {7'd0,(kernel[2][3] ~^ image[18][8])} + {7'd0,(kernel[2][4] ~^ image[18][9])} + {7'd0,(kernel[3][0] ~^ image[19][5])} + {7'd0,(kernel[3][1] ~^ image[19][6])} + {7'd0,(kernel[3][2] ~^ image[19][7])} + {7'd0,(kernel[3][3] ~^ image[19][8])} + {7'd0,(kernel[3][4] ~^ image[19][9])} + {7'd0,(kernel[4][0] ~^ image[20][5])} + {7'd0,(kernel[4][1] ~^ image[20][6])} + {7'd0,(kernel[4][2] ~^ image[20][7])} + {7'd0,(kernel[4][3] ~^ image[20][8])} + {7'd0,(kernel[4][4] ~^ image[20][9])};
assign out_fmap[16][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[16][6])} + {7'd0,(kernel[0][1] ~^ image[16][7])} + {7'd0,(kernel[0][2] ~^ image[16][8])} + {7'd0,(kernel[0][3] ~^ image[16][9])} + {7'd0,(kernel[0][4] ~^ image[16][10])} + {7'd0,(kernel[1][0] ~^ image[17][6])} + {7'd0,(kernel[1][1] ~^ image[17][7])} + {7'd0,(kernel[1][2] ~^ image[17][8])} + {7'd0,(kernel[1][3] ~^ image[17][9])} + {7'd0,(kernel[1][4] ~^ image[17][10])} + {7'd0,(kernel[2][0] ~^ image[18][6])} + {7'd0,(kernel[2][1] ~^ image[18][7])} + {7'd0,(kernel[2][2] ~^ image[18][8])} + {7'd0,(kernel[2][3] ~^ image[18][9])} + {7'd0,(kernel[2][4] ~^ image[18][10])} + {7'd0,(kernel[3][0] ~^ image[19][6])} + {7'd0,(kernel[3][1] ~^ image[19][7])} + {7'd0,(kernel[3][2] ~^ image[19][8])} + {7'd0,(kernel[3][3] ~^ image[19][9])} + {7'd0,(kernel[3][4] ~^ image[19][10])} + {7'd0,(kernel[4][0] ~^ image[20][6])} + {7'd0,(kernel[4][1] ~^ image[20][7])} + {7'd0,(kernel[4][2] ~^ image[20][8])} + {7'd0,(kernel[4][3] ~^ image[20][9])} + {7'd0,(kernel[4][4] ~^ image[20][10])};
assign out_fmap[16][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[16][7])} + {7'd0,(kernel[0][1] ~^ image[16][8])} + {7'd0,(kernel[0][2] ~^ image[16][9])} + {7'd0,(kernel[0][3] ~^ image[16][10])} + {7'd0,(kernel[0][4] ~^ image[16][11])} + {7'd0,(kernel[1][0] ~^ image[17][7])} + {7'd0,(kernel[1][1] ~^ image[17][8])} + {7'd0,(kernel[1][2] ~^ image[17][9])} + {7'd0,(kernel[1][3] ~^ image[17][10])} + {7'd0,(kernel[1][4] ~^ image[17][11])} + {7'd0,(kernel[2][0] ~^ image[18][7])} + {7'd0,(kernel[2][1] ~^ image[18][8])} + {7'd0,(kernel[2][2] ~^ image[18][9])} + {7'd0,(kernel[2][3] ~^ image[18][10])} + {7'd0,(kernel[2][4] ~^ image[18][11])} + {7'd0,(kernel[3][0] ~^ image[19][7])} + {7'd0,(kernel[3][1] ~^ image[19][8])} + {7'd0,(kernel[3][2] ~^ image[19][9])} + {7'd0,(kernel[3][3] ~^ image[19][10])} + {7'd0,(kernel[3][4] ~^ image[19][11])} + {7'd0,(kernel[4][0] ~^ image[20][7])} + {7'd0,(kernel[4][1] ~^ image[20][8])} + {7'd0,(kernel[4][2] ~^ image[20][9])} + {7'd0,(kernel[4][3] ~^ image[20][10])} + {7'd0,(kernel[4][4] ~^ image[20][11])};
assign out_fmap[16][8][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[16][8])} + {7'd0,(kernel[0][1] ~^ image[16][9])} + {7'd0,(kernel[0][2] ~^ image[16][10])} + {7'd0,(kernel[0][3] ~^ image[16][11])} + {7'd0,(kernel[0][4] ~^ image[16][12])} + {7'd0,(kernel[1][0] ~^ image[17][8])} + {7'd0,(kernel[1][1] ~^ image[17][9])} + {7'd0,(kernel[1][2] ~^ image[17][10])} + {7'd0,(kernel[1][3] ~^ image[17][11])} + {7'd0,(kernel[1][4] ~^ image[17][12])} + {7'd0,(kernel[2][0] ~^ image[18][8])} + {7'd0,(kernel[2][1] ~^ image[18][9])} + {7'd0,(kernel[2][2] ~^ image[18][10])} + {7'd0,(kernel[2][3] ~^ image[18][11])} + {7'd0,(kernel[2][4] ~^ image[18][12])} + {7'd0,(kernel[3][0] ~^ image[19][8])} + {7'd0,(kernel[3][1] ~^ image[19][9])} + {7'd0,(kernel[3][2] ~^ image[19][10])} + {7'd0,(kernel[3][3] ~^ image[19][11])} + {7'd0,(kernel[3][4] ~^ image[19][12])} + {7'd0,(kernel[4][0] ~^ image[20][8])} + {7'd0,(kernel[4][1] ~^ image[20][9])} + {7'd0,(kernel[4][2] ~^ image[20][10])} + {7'd0,(kernel[4][3] ~^ image[20][11])} + {7'd0,(kernel[4][4] ~^ image[20][12])};
assign out_fmap[16][9][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[16][9])} + {7'd0,(kernel[0][1] ~^ image[16][10])} + {7'd0,(kernel[0][2] ~^ image[16][11])} + {7'd0,(kernel[0][3] ~^ image[16][12])} + {7'd0,(kernel[0][4] ~^ image[16][13])} + {7'd0,(kernel[1][0] ~^ image[17][9])} + {7'd0,(kernel[1][1] ~^ image[17][10])} + {7'd0,(kernel[1][2] ~^ image[17][11])} + {7'd0,(kernel[1][3] ~^ image[17][12])} + {7'd0,(kernel[1][4] ~^ image[17][13])} + {7'd0,(kernel[2][0] ~^ image[18][9])} + {7'd0,(kernel[2][1] ~^ image[18][10])} + {7'd0,(kernel[2][2] ~^ image[18][11])} + {7'd0,(kernel[2][3] ~^ image[18][12])} + {7'd0,(kernel[2][4] ~^ image[18][13])} + {7'd0,(kernel[3][0] ~^ image[19][9])} + {7'd0,(kernel[3][1] ~^ image[19][10])} + {7'd0,(kernel[3][2] ~^ image[19][11])} + {7'd0,(kernel[3][3] ~^ image[19][12])} + {7'd0,(kernel[3][4] ~^ image[19][13])} + {7'd0,(kernel[4][0] ~^ image[20][9])} + {7'd0,(kernel[4][1] ~^ image[20][10])} + {7'd0,(kernel[4][2] ~^ image[20][11])} + {7'd0,(kernel[4][3] ~^ image[20][12])} + {7'd0,(kernel[4][4] ~^ image[20][13])};
assign out_fmap[16][10][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[16][10])} + {7'd0,(kernel[0][1] ~^ image[16][11])} + {7'd0,(kernel[0][2] ~^ image[16][12])} + {7'd0,(kernel[0][3] ~^ image[16][13])} + {7'd0,(kernel[0][4] ~^ image[16][14])} + {7'd0,(kernel[1][0] ~^ image[17][10])} + {7'd0,(kernel[1][1] ~^ image[17][11])} + {7'd0,(kernel[1][2] ~^ image[17][12])} + {7'd0,(kernel[1][3] ~^ image[17][13])} + {7'd0,(kernel[1][4] ~^ image[17][14])} + {7'd0,(kernel[2][0] ~^ image[18][10])} + {7'd0,(kernel[2][1] ~^ image[18][11])} + {7'd0,(kernel[2][2] ~^ image[18][12])} + {7'd0,(kernel[2][3] ~^ image[18][13])} + {7'd0,(kernel[2][4] ~^ image[18][14])} + {7'd0,(kernel[3][0] ~^ image[19][10])} + {7'd0,(kernel[3][1] ~^ image[19][11])} + {7'd0,(kernel[3][2] ~^ image[19][12])} + {7'd0,(kernel[3][3] ~^ image[19][13])} + {7'd0,(kernel[3][4] ~^ image[19][14])} + {7'd0,(kernel[4][0] ~^ image[20][10])} + {7'd0,(kernel[4][1] ~^ image[20][11])} + {7'd0,(kernel[4][2] ~^ image[20][12])} + {7'd0,(kernel[4][3] ~^ image[20][13])} + {7'd0,(kernel[4][4] ~^ image[20][14])};
assign out_fmap[16][11][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[16][11])} + {7'd0,(kernel[0][1] ~^ image[16][12])} + {7'd0,(kernel[0][2] ~^ image[16][13])} + {7'd0,(kernel[0][3] ~^ image[16][14])} + {7'd0,(kernel[0][4] ~^ image[16][15])} + {7'd0,(kernel[1][0] ~^ image[17][11])} + {7'd0,(kernel[1][1] ~^ image[17][12])} + {7'd0,(kernel[1][2] ~^ image[17][13])} + {7'd0,(kernel[1][3] ~^ image[17][14])} + {7'd0,(kernel[1][4] ~^ image[17][15])} + {7'd0,(kernel[2][0] ~^ image[18][11])} + {7'd0,(kernel[2][1] ~^ image[18][12])} + {7'd0,(kernel[2][2] ~^ image[18][13])} + {7'd0,(kernel[2][3] ~^ image[18][14])} + {7'd0,(kernel[2][4] ~^ image[18][15])} + {7'd0,(kernel[3][0] ~^ image[19][11])} + {7'd0,(kernel[3][1] ~^ image[19][12])} + {7'd0,(kernel[3][2] ~^ image[19][13])} + {7'd0,(kernel[3][3] ~^ image[19][14])} + {7'd0,(kernel[3][4] ~^ image[19][15])} + {7'd0,(kernel[4][0] ~^ image[20][11])} + {7'd0,(kernel[4][1] ~^ image[20][12])} + {7'd0,(kernel[4][2] ~^ image[20][13])} + {7'd0,(kernel[4][3] ~^ image[20][14])} + {7'd0,(kernel[4][4] ~^ image[20][15])};
assign out_fmap[16][12][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[16][12])} + {7'd0,(kernel[0][1] ~^ image[16][13])} + {7'd0,(kernel[0][2] ~^ image[16][14])} + {7'd0,(kernel[0][3] ~^ image[16][15])} + {7'd0,(kernel[0][4] ~^ image[16][16])} + {7'd0,(kernel[1][0] ~^ image[17][12])} + {7'd0,(kernel[1][1] ~^ image[17][13])} + {7'd0,(kernel[1][2] ~^ image[17][14])} + {7'd0,(kernel[1][3] ~^ image[17][15])} + {7'd0,(kernel[1][4] ~^ image[17][16])} + {7'd0,(kernel[2][0] ~^ image[18][12])} + {7'd0,(kernel[2][1] ~^ image[18][13])} + {7'd0,(kernel[2][2] ~^ image[18][14])} + {7'd0,(kernel[2][3] ~^ image[18][15])} + {7'd0,(kernel[2][4] ~^ image[18][16])} + {7'd0,(kernel[3][0] ~^ image[19][12])} + {7'd0,(kernel[3][1] ~^ image[19][13])} + {7'd0,(kernel[3][2] ~^ image[19][14])} + {7'd0,(kernel[3][3] ~^ image[19][15])} + {7'd0,(kernel[3][4] ~^ image[19][16])} + {7'd0,(kernel[4][0] ~^ image[20][12])} + {7'd0,(kernel[4][1] ~^ image[20][13])} + {7'd0,(kernel[4][2] ~^ image[20][14])} + {7'd0,(kernel[4][3] ~^ image[20][15])} + {7'd0,(kernel[4][4] ~^ image[20][16])};
assign out_fmap[16][13][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[16][13])} + {7'd0,(kernel[0][1] ~^ image[16][14])} + {7'd0,(kernel[0][2] ~^ image[16][15])} + {7'd0,(kernel[0][3] ~^ image[16][16])} + {7'd0,(kernel[0][4] ~^ image[16][17])} + {7'd0,(kernel[1][0] ~^ image[17][13])} + {7'd0,(kernel[1][1] ~^ image[17][14])} + {7'd0,(kernel[1][2] ~^ image[17][15])} + {7'd0,(kernel[1][3] ~^ image[17][16])} + {7'd0,(kernel[1][4] ~^ image[17][17])} + {7'd0,(kernel[2][0] ~^ image[18][13])} + {7'd0,(kernel[2][1] ~^ image[18][14])} + {7'd0,(kernel[2][2] ~^ image[18][15])} + {7'd0,(kernel[2][3] ~^ image[18][16])} + {7'd0,(kernel[2][4] ~^ image[18][17])} + {7'd0,(kernel[3][0] ~^ image[19][13])} + {7'd0,(kernel[3][1] ~^ image[19][14])} + {7'd0,(kernel[3][2] ~^ image[19][15])} + {7'd0,(kernel[3][3] ~^ image[19][16])} + {7'd0,(kernel[3][4] ~^ image[19][17])} + {7'd0,(kernel[4][0] ~^ image[20][13])} + {7'd0,(kernel[4][1] ~^ image[20][14])} + {7'd0,(kernel[4][2] ~^ image[20][15])} + {7'd0,(kernel[4][3] ~^ image[20][16])} + {7'd0,(kernel[4][4] ~^ image[20][17])};
assign out_fmap[16][14][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[16][14])} + {7'd0,(kernel[0][1] ~^ image[16][15])} + {7'd0,(kernel[0][2] ~^ image[16][16])} + {7'd0,(kernel[0][3] ~^ image[16][17])} + {7'd0,(kernel[0][4] ~^ image[16][18])} + {7'd0,(kernel[1][0] ~^ image[17][14])} + {7'd0,(kernel[1][1] ~^ image[17][15])} + {7'd0,(kernel[1][2] ~^ image[17][16])} + {7'd0,(kernel[1][3] ~^ image[17][17])} + {7'd0,(kernel[1][4] ~^ image[17][18])} + {7'd0,(kernel[2][0] ~^ image[18][14])} + {7'd0,(kernel[2][1] ~^ image[18][15])} + {7'd0,(kernel[2][2] ~^ image[18][16])} + {7'd0,(kernel[2][3] ~^ image[18][17])} + {7'd0,(kernel[2][4] ~^ image[18][18])} + {7'd0,(kernel[3][0] ~^ image[19][14])} + {7'd0,(kernel[3][1] ~^ image[19][15])} + {7'd0,(kernel[3][2] ~^ image[19][16])} + {7'd0,(kernel[3][3] ~^ image[19][17])} + {7'd0,(kernel[3][4] ~^ image[19][18])} + {7'd0,(kernel[4][0] ~^ image[20][14])} + {7'd0,(kernel[4][1] ~^ image[20][15])} + {7'd0,(kernel[4][2] ~^ image[20][16])} + {7'd0,(kernel[4][3] ~^ image[20][17])} + {7'd0,(kernel[4][4] ~^ image[20][18])};
assign out_fmap[16][15][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[16][15])} + {7'd0,(kernel[0][1] ~^ image[16][16])} + {7'd0,(kernel[0][2] ~^ image[16][17])} + {7'd0,(kernel[0][3] ~^ image[16][18])} + {7'd0,(kernel[0][4] ~^ image[16][19])} + {7'd0,(kernel[1][0] ~^ image[17][15])} + {7'd0,(kernel[1][1] ~^ image[17][16])} + {7'd0,(kernel[1][2] ~^ image[17][17])} + {7'd0,(kernel[1][3] ~^ image[17][18])} + {7'd0,(kernel[1][4] ~^ image[17][19])} + {7'd0,(kernel[2][0] ~^ image[18][15])} + {7'd0,(kernel[2][1] ~^ image[18][16])} + {7'd0,(kernel[2][2] ~^ image[18][17])} + {7'd0,(kernel[2][3] ~^ image[18][18])} + {7'd0,(kernel[2][4] ~^ image[18][19])} + {7'd0,(kernel[3][0] ~^ image[19][15])} + {7'd0,(kernel[3][1] ~^ image[19][16])} + {7'd0,(kernel[3][2] ~^ image[19][17])} + {7'd0,(kernel[3][3] ~^ image[19][18])} + {7'd0,(kernel[3][4] ~^ image[19][19])} + {7'd0,(kernel[4][0] ~^ image[20][15])} + {7'd0,(kernel[4][1] ~^ image[20][16])} + {7'd0,(kernel[4][2] ~^ image[20][17])} + {7'd0,(kernel[4][3] ~^ image[20][18])} + {7'd0,(kernel[4][4] ~^ image[20][19])};
assign out_fmap[16][16][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[16][16])} + {7'd0,(kernel[0][1] ~^ image[16][17])} + {7'd0,(kernel[0][2] ~^ image[16][18])} + {7'd0,(kernel[0][3] ~^ image[16][19])} + {7'd0,(kernel[0][4] ~^ image[16][20])} + {7'd0,(kernel[1][0] ~^ image[17][16])} + {7'd0,(kernel[1][1] ~^ image[17][17])} + {7'd0,(kernel[1][2] ~^ image[17][18])} + {7'd0,(kernel[1][3] ~^ image[17][19])} + {7'd0,(kernel[1][4] ~^ image[17][20])} + {7'd0,(kernel[2][0] ~^ image[18][16])} + {7'd0,(kernel[2][1] ~^ image[18][17])} + {7'd0,(kernel[2][2] ~^ image[18][18])} + {7'd0,(kernel[2][3] ~^ image[18][19])} + {7'd0,(kernel[2][4] ~^ image[18][20])} + {7'd0,(kernel[3][0] ~^ image[19][16])} + {7'd0,(kernel[3][1] ~^ image[19][17])} + {7'd0,(kernel[3][2] ~^ image[19][18])} + {7'd0,(kernel[3][3] ~^ image[19][19])} + {7'd0,(kernel[3][4] ~^ image[19][20])} + {7'd0,(kernel[4][0] ~^ image[20][16])} + {7'd0,(kernel[4][1] ~^ image[20][17])} + {7'd0,(kernel[4][2] ~^ image[20][18])} + {7'd0,(kernel[4][3] ~^ image[20][19])} + {7'd0,(kernel[4][4] ~^ image[20][20])};
assign out_fmap[16][17][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[16][17])} + {7'd0,(kernel[0][1] ~^ image[16][18])} + {7'd0,(kernel[0][2] ~^ image[16][19])} + {7'd0,(kernel[0][3] ~^ image[16][20])} + {7'd0,(kernel[0][4] ~^ image[16][21])} + {7'd0,(kernel[1][0] ~^ image[17][17])} + {7'd0,(kernel[1][1] ~^ image[17][18])} + {7'd0,(kernel[1][2] ~^ image[17][19])} + {7'd0,(kernel[1][3] ~^ image[17][20])} + {7'd0,(kernel[1][4] ~^ image[17][21])} + {7'd0,(kernel[2][0] ~^ image[18][17])} + {7'd0,(kernel[2][1] ~^ image[18][18])} + {7'd0,(kernel[2][2] ~^ image[18][19])} + {7'd0,(kernel[2][3] ~^ image[18][20])} + {7'd0,(kernel[2][4] ~^ image[18][21])} + {7'd0,(kernel[3][0] ~^ image[19][17])} + {7'd0,(kernel[3][1] ~^ image[19][18])} + {7'd0,(kernel[3][2] ~^ image[19][19])} + {7'd0,(kernel[3][3] ~^ image[19][20])} + {7'd0,(kernel[3][4] ~^ image[19][21])} + {7'd0,(kernel[4][0] ~^ image[20][17])} + {7'd0,(kernel[4][1] ~^ image[20][18])} + {7'd0,(kernel[4][2] ~^ image[20][19])} + {7'd0,(kernel[4][3] ~^ image[20][20])} + {7'd0,(kernel[4][4] ~^ image[20][21])};
assign out_fmap[16][18][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[16][18])} + {7'd0,(kernel[0][1] ~^ image[16][19])} + {7'd0,(kernel[0][2] ~^ image[16][20])} + {7'd0,(kernel[0][3] ~^ image[16][21])} + {7'd0,(kernel[0][4] ~^ image[16][22])} + {7'd0,(kernel[1][0] ~^ image[17][18])} + {7'd0,(kernel[1][1] ~^ image[17][19])} + {7'd0,(kernel[1][2] ~^ image[17][20])} + {7'd0,(kernel[1][3] ~^ image[17][21])} + {7'd0,(kernel[1][4] ~^ image[17][22])} + {7'd0,(kernel[2][0] ~^ image[18][18])} + {7'd0,(kernel[2][1] ~^ image[18][19])} + {7'd0,(kernel[2][2] ~^ image[18][20])} + {7'd0,(kernel[2][3] ~^ image[18][21])} + {7'd0,(kernel[2][4] ~^ image[18][22])} + {7'd0,(kernel[3][0] ~^ image[19][18])} + {7'd0,(kernel[3][1] ~^ image[19][19])} + {7'd0,(kernel[3][2] ~^ image[19][20])} + {7'd0,(kernel[3][3] ~^ image[19][21])} + {7'd0,(kernel[3][4] ~^ image[19][22])} + {7'd0,(kernel[4][0] ~^ image[20][18])} + {7'd0,(kernel[4][1] ~^ image[20][19])} + {7'd0,(kernel[4][2] ~^ image[20][20])} + {7'd0,(kernel[4][3] ~^ image[20][21])} + {7'd0,(kernel[4][4] ~^ image[20][22])};
assign out_fmap[16][19][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[16][19])} + {7'd0,(kernel[0][1] ~^ image[16][20])} + {7'd0,(kernel[0][2] ~^ image[16][21])} + {7'd0,(kernel[0][3] ~^ image[16][22])} + {7'd0,(kernel[0][4] ~^ image[16][23])} + {7'd0,(kernel[1][0] ~^ image[17][19])} + {7'd0,(kernel[1][1] ~^ image[17][20])} + {7'd0,(kernel[1][2] ~^ image[17][21])} + {7'd0,(kernel[1][3] ~^ image[17][22])} + {7'd0,(kernel[1][4] ~^ image[17][23])} + {7'd0,(kernel[2][0] ~^ image[18][19])} + {7'd0,(kernel[2][1] ~^ image[18][20])} + {7'd0,(kernel[2][2] ~^ image[18][21])} + {7'd0,(kernel[2][3] ~^ image[18][22])} + {7'd0,(kernel[2][4] ~^ image[18][23])} + {7'd0,(kernel[3][0] ~^ image[19][19])} + {7'd0,(kernel[3][1] ~^ image[19][20])} + {7'd0,(kernel[3][2] ~^ image[19][21])} + {7'd0,(kernel[3][3] ~^ image[19][22])} + {7'd0,(kernel[3][4] ~^ image[19][23])} + {7'd0,(kernel[4][0] ~^ image[20][19])} + {7'd0,(kernel[4][1] ~^ image[20][20])} + {7'd0,(kernel[4][2] ~^ image[20][21])} + {7'd0,(kernel[4][3] ~^ image[20][22])} + {7'd0,(kernel[4][4] ~^ image[20][23])};
assign out_fmap[16][20][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[16][20])} + {7'd0,(kernel[0][1] ~^ image[16][21])} + {7'd0,(kernel[0][2] ~^ image[16][22])} + {7'd0,(kernel[0][3] ~^ image[16][23])} + {7'd0,(kernel[0][4] ~^ image[16][24])} + {7'd0,(kernel[1][0] ~^ image[17][20])} + {7'd0,(kernel[1][1] ~^ image[17][21])} + {7'd0,(kernel[1][2] ~^ image[17][22])} + {7'd0,(kernel[1][3] ~^ image[17][23])} + {7'd0,(kernel[1][4] ~^ image[17][24])} + {7'd0,(kernel[2][0] ~^ image[18][20])} + {7'd0,(kernel[2][1] ~^ image[18][21])} + {7'd0,(kernel[2][2] ~^ image[18][22])} + {7'd0,(kernel[2][3] ~^ image[18][23])} + {7'd0,(kernel[2][4] ~^ image[18][24])} + {7'd0,(kernel[3][0] ~^ image[19][20])} + {7'd0,(kernel[3][1] ~^ image[19][21])} + {7'd0,(kernel[3][2] ~^ image[19][22])} + {7'd0,(kernel[3][3] ~^ image[19][23])} + {7'd0,(kernel[3][4] ~^ image[19][24])} + {7'd0,(kernel[4][0] ~^ image[20][20])} + {7'd0,(kernel[4][1] ~^ image[20][21])} + {7'd0,(kernel[4][2] ~^ image[20][22])} + {7'd0,(kernel[4][3] ~^ image[20][23])} + {7'd0,(kernel[4][4] ~^ image[20][24])};
assign out_fmap[16][21][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[16][21])} + {7'd0,(kernel[0][1] ~^ image[16][22])} + {7'd0,(kernel[0][2] ~^ image[16][23])} + {7'd0,(kernel[0][3] ~^ image[16][24])} + {7'd0,(kernel[0][4] ~^ image[16][25])} + {7'd0,(kernel[1][0] ~^ image[17][21])} + {7'd0,(kernel[1][1] ~^ image[17][22])} + {7'd0,(kernel[1][2] ~^ image[17][23])} + {7'd0,(kernel[1][3] ~^ image[17][24])} + {7'd0,(kernel[1][4] ~^ image[17][25])} + {7'd0,(kernel[2][0] ~^ image[18][21])} + {7'd0,(kernel[2][1] ~^ image[18][22])} + {7'd0,(kernel[2][2] ~^ image[18][23])} + {7'd0,(kernel[2][3] ~^ image[18][24])} + {7'd0,(kernel[2][4] ~^ image[18][25])} + {7'd0,(kernel[3][0] ~^ image[19][21])} + {7'd0,(kernel[3][1] ~^ image[19][22])} + {7'd0,(kernel[3][2] ~^ image[19][23])} + {7'd0,(kernel[3][3] ~^ image[19][24])} + {7'd0,(kernel[3][4] ~^ image[19][25])} + {7'd0,(kernel[4][0] ~^ image[20][21])} + {7'd0,(kernel[4][1] ~^ image[20][22])} + {7'd0,(kernel[4][2] ~^ image[20][23])} + {7'd0,(kernel[4][3] ~^ image[20][24])} + {7'd0,(kernel[4][4] ~^ image[20][25])};
assign out_fmap[16][22][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[16][22])} + {7'd0,(kernel[0][1] ~^ image[16][23])} + {7'd0,(kernel[0][2] ~^ image[16][24])} + {7'd0,(kernel[0][3] ~^ image[16][25])} + {7'd0,(kernel[0][4] ~^ image[16][26])} + {7'd0,(kernel[1][0] ~^ image[17][22])} + {7'd0,(kernel[1][1] ~^ image[17][23])} + {7'd0,(kernel[1][2] ~^ image[17][24])} + {7'd0,(kernel[1][3] ~^ image[17][25])} + {7'd0,(kernel[1][4] ~^ image[17][26])} + {7'd0,(kernel[2][0] ~^ image[18][22])} + {7'd0,(kernel[2][1] ~^ image[18][23])} + {7'd0,(kernel[2][2] ~^ image[18][24])} + {7'd0,(kernel[2][3] ~^ image[18][25])} + {7'd0,(kernel[2][4] ~^ image[18][26])} + {7'd0,(kernel[3][0] ~^ image[19][22])} + {7'd0,(kernel[3][1] ~^ image[19][23])} + {7'd0,(kernel[3][2] ~^ image[19][24])} + {7'd0,(kernel[3][3] ~^ image[19][25])} + {7'd0,(kernel[3][4] ~^ image[19][26])} + {7'd0,(kernel[4][0] ~^ image[20][22])} + {7'd0,(kernel[4][1] ~^ image[20][23])} + {7'd0,(kernel[4][2] ~^ image[20][24])} + {7'd0,(kernel[4][3] ~^ image[20][25])} + {7'd0,(kernel[4][4] ~^ image[20][26])};
assign out_fmap[16][23][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[16][23])} + {7'd0,(kernel[0][1] ~^ image[16][24])} + {7'd0,(kernel[0][2] ~^ image[16][25])} + {7'd0,(kernel[0][3] ~^ image[16][26])} + {7'd0,(kernel[0][4] ~^ image[16][27])} + {7'd0,(kernel[1][0] ~^ image[17][23])} + {7'd0,(kernel[1][1] ~^ image[17][24])} + {7'd0,(kernel[1][2] ~^ image[17][25])} + {7'd0,(kernel[1][3] ~^ image[17][26])} + {7'd0,(kernel[1][4] ~^ image[17][27])} + {7'd0,(kernel[2][0] ~^ image[18][23])} + {7'd0,(kernel[2][1] ~^ image[18][24])} + {7'd0,(kernel[2][2] ~^ image[18][25])} + {7'd0,(kernel[2][3] ~^ image[18][26])} + {7'd0,(kernel[2][4] ~^ image[18][27])} + {7'd0,(kernel[3][0] ~^ image[19][23])} + {7'd0,(kernel[3][1] ~^ image[19][24])} + {7'd0,(kernel[3][2] ~^ image[19][25])} + {7'd0,(kernel[3][3] ~^ image[19][26])} + {7'd0,(kernel[3][4] ~^ image[19][27])} + {7'd0,(kernel[4][0] ~^ image[20][23])} + {7'd0,(kernel[4][1] ~^ image[20][24])} + {7'd0,(kernel[4][2] ~^ image[20][25])} + {7'd0,(kernel[4][3] ~^ image[20][26])} + {7'd0,(kernel[4][4] ~^ image[20][27])};
assign out_fmap[17][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[17][0])} + {7'd0,(kernel[0][1] ~^ image[17][1])} + {7'd0,(kernel[0][2] ~^ image[17][2])} + {7'd0,(kernel[0][3] ~^ image[17][3])} + {7'd0,(kernel[0][4] ~^ image[17][4])} + {7'd0,(kernel[1][0] ~^ image[18][0])} + {7'd0,(kernel[1][1] ~^ image[18][1])} + {7'd0,(kernel[1][2] ~^ image[18][2])} + {7'd0,(kernel[1][3] ~^ image[18][3])} + {7'd0,(kernel[1][4] ~^ image[18][4])} + {7'd0,(kernel[2][0] ~^ image[19][0])} + {7'd0,(kernel[2][1] ~^ image[19][1])} + {7'd0,(kernel[2][2] ~^ image[19][2])} + {7'd0,(kernel[2][3] ~^ image[19][3])} + {7'd0,(kernel[2][4] ~^ image[19][4])} + {7'd0,(kernel[3][0] ~^ image[20][0])} + {7'd0,(kernel[3][1] ~^ image[20][1])} + {7'd0,(kernel[3][2] ~^ image[20][2])} + {7'd0,(kernel[3][3] ~^ image[20][3])} + {7'd0,(kernel[3][4] ~^ image[20][4])} + {7'd0,(kernel[4][0] ~^ image[21][0])} + {7'd0,(kernel[4][1] ~^ image[21][1])} + {7'd0,(kernel[4][2] ~^ image[21][2])} + {7'd0,(kernel[4][3] ~^ image[21][3])} + {7'd0,(kernel[4][4] ~^ image[21][4])};
assign out_fmap[17][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[17][1])} + {7'd0,(kernel[0][1] ~^ image[17][2])} + {7'd0,(kernel[0][2] ~^ image[17][3])} + {7'd0,(kernel[0][3] ~^ image[17][4])} + {7'd0,(kernel[0][4] ~^ image[17][5])} + {7'd0,(kernel[1][0] ~^ image[18][1])} + {7'd0,(kernel[1][1] ~^ image[18][2])} + {7'd0,(kernel[1][2] ~^ image[18][3])} + {7'd0,(kernel[1][3] ~^ image[18][4])} + {7'd0,(kernel[1][4] ~^ image[18][5])} + {7'd0,(kernel[2][0] ~^ image[19][1])} + {7'd0,(kernel[2][1] ~^ image[19][2])} + {7'd0,(kernel[2][2] ~^ image[19][3])} + {7'd0,(kernel[2][3] ~^ image[19][4])} + {7'd0,(kernel[2][4] ~^ image[19][5])} + {7'd0,(kernel[3][0] ~^ image[20][1])} + {7'd0,(kernel[3][1] ~^ image[20][2])} + {7'd0,(kernel[3][2] ~^ image[20][3])} + {7'd0,(kernel[3][3] ~^ image[20][4])} + {7'd0,(kernel[3][4] ~^ image[20][5])} + {7'd0,(kernel[4][0] ~^ image[21][1])} + {7'd0,(kernel[4][1] ~^ image[21][2])} + {7'd0,(kernel[4][2] ~^ image[21][3])} + {7'd0,(kernel[4][3] ~^ image[21][4])} + {7'd0,(kernel[4][4] ~^ image[21][5])};
assign out_fmap[17][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[17][2])} + {7'd0,(kernel[0][1] ~^ image[17][3])} + {7'd0,(kernel[0][2] ~^ image[17][4])} + {7'd0,(kernel[0][3] ~^ image[17][5])} + {7'd0,(kernel[0][4] ~^ image[17][6])} + {7'd0,(kernel[1][0] ~^ image[18][2])} + {7'd0,(kernel[1][1] ~^ image[18][3])} + {7'd0,(kernel[1][2] ~^ image[18][4])} + {7'd0,(kernel[1][3] ~^ image[18][5])} + {7'd0,(kernel[1][4] ~^ image[18][6])} + {7'd0,(kernel[2][0] ~^ image[19][2])} + {7'd0,(kernel[2][1] ~^ image[19][3])} + {7'd0,(kernel[2][2] ~^ image[19][4])} + {7'd0,(kernel[2][3] ~^ image[19][5])} + {7'd0,(kernel[2][4] ~^ image[19][6])} + {7'd0,(kernel[3][0] ~^ image[20][2])} + {7'd0,(kernel[3][1] ~^ image[20][3])} + {7'd0,(kernel[3][2] ~^ image[20][4])} + {7'd0,(kernel[3][3] ~^ image[20][5])} + {7'd0,(kernel[3][4] ~^ image[20][6])} + {7'd0,(kernel[4][0] ~^ image[21][2])} + {7'd0,(kernel[4][1] ~^ image[21][3])} + {7'd0,(kernel[4][2] ~^ image[21][4])} + {7'd0,(kernel[4][3] ~^ image[21][5])} + {7'd0,(kernel[4][4] ~^ image[21][6])};
assign out_fmap[17][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[17][3])} + {7'd0,(kernel[0][1] ~^ image[17][4])} + {7'd0,(kernel[0][2] ~^ image[17][5])} + {7'd0,(kernel[0][3] ~^ image[17][6])} + {7'd0,(kernel[0][4] ~^ image[17][7])} + {7'd0,(kernel[1][0] ~^ image[18][3])} + {7'd0,(kernel[1][1] ~^ image[18][4])} + {7'd0,(kernel[1][2] ~^ image[18][5])} + {7'd0,(kernel[1][3] ~^ image[18][6])} + {7'd0,(kernel[1][4] ~^ image[18][7])} + {7'd0,(kernel[2][0] ~^ image[19][3])} + {7'd0,(kernel[2][1] ~^ image[19][4])} + {7'd0,(kernel[2][2] ~^ image[19][5])} + {7'd0,(kernel[2][3] ~^ image[19][6])} + {7'd0,(kernel[2][4] ~^ image[19][7])} + {7'd0,(kernel[3][0] ~^ image[20][3])} + {7'd0,(kernel[3][1] ~^ image[20][4])} + {7'd0,(kernel[3][2] ~^ image[20][5])} + {7'd0,(kernel[3][3] ~^ image[20][6])} + {7'd0,(kernel[3][4] ~^ image[20][7])} + {7'd0,(kernel[4][0] ~^ image[21][3])} + {7'd0,(kernel[4][1] ~^ image[21][4])} + {7'd0,(kernel[4][2] ~^ image[21][5])} + {7'd0,(kernel[4][3] ~^ image[21][6])} + {7'd0,(kernel[4][4] ~^ image[21][7])};
assign out_fmap[17][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[17][4])} + {7'd0,(kernel[0][1] ~^ image[17][5])} + {7'd0,(kernel[0][2] ~^ image[17][6])} + {7'd0,(kernel[0][3] ~^ image[17][7])} + {7'd0,(kernel[0][4] ~^ image[17][8])} + {7'd0,(kernel[1][0] ~^ image[18][4])} + {7'd0,(kernel[1][1] ~^ image[18][5])} + {7'd0,(kernel[1][2] ~^ image[18][6])} + {7'd0,(kernel[1][3] ~^ image[18][7])} + {7'd0,(kernel[1][4] ~^ image[18][8])} + {7'd0,(kernel[2][0] ~^ image[19][4])} + {7'd0,(kernel[2][1] ~^ image[19][5])} + {7'd0,(kernel[2][2] ~^ image[19][6])} + {7'd0,(kernel[2][3] ~^ image[19][7])} + {7'd0,(kernel[2][4] ~^ image[19][8])} + {7'd0,(kernel[3][0] ~^ image[20][4])} + {7'd0,(kernel[3][1] ~^ image[20][5])} + {7'd0,(kernel[3][2] ~^ image[20][6])} + {7'd0,(kernel[3][3] ~^ image[20][7])} + {7'd0,(kernel[3][4] ~^ image[20][8])} + {7'd0,(kernel[4][0] ~^ image[21][4])} + {7'd0,(kernel[4][1] ~^ image[21][5])} + {7'd0,(kernel[4][2] ~^ image[21][6])} + {7'd0,(kernel[4][3] ~^ image[21][7])} + {7'd0,(kernel[4][4] ~^ image[21][8])};
assign out_fmap[17][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[17][5])} + {7'd0,(kernel[0][1] ~^ image[17][6])} + {7'd0,(kernel[0][2] ~^ image[17][7])} + {7'd0,(kernel[0][3] ~^ image[17][8])} + {7'd0,(kernel[0][4] ~^ image[17][9])} + {7'd0,(kernel[1][0] ~^ image[18][5])} + {7'd0,(kernel[1][1] ~^ image[18][6])} + {7'd0,(kernel[1][2] ~^ image[18][7])} + {7'd0,(kernel[1][3] ~^ image[18][8])} + {7'd0,(kernel[1][4] ~^ image[18][9])} + {7'd0,(kernel[2][0] ~^ image[19][5])} + {7'd0,(kernel[2][1] ~^ image[19][6])} + {7'd0,(kernel[2][2] ~^ image[19][7])} + {7'd0,(kernel[2][3] ~^ image[19][8])} + {7'd0,(kernel[2][4] ~^ image[19][9])} + {7'd0,(kernel[3][0] ~^ image[20][5])} + {7'd0,(kernel[3][1] ~^ image[20][6])} + {7'd0,(kernel[3][2] ~^ image[20][7])} + {7'd0,(kernel[3][3] ~^ image[20][8])} + {7'd0,(kernel[3][4] ~^ image[20][9])} + {7'd0,(kernel[4][0] ~^ image[21][5])} + {7'd0,(kernel[4][1] ~^ image[21][6])} + {7'd0,(kernel[4][2] ~^ image[21][7])} + {7'd0,(kernel[4][3] ~^ image[21][8])} + {7'd0,(kernel[4][4] ~^ image[21][9])};
assign out_fmap[17][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[17][6])} + {7'd0,(kernel[0][1] ~^ image[17][7])} + {7'd0,(kernel[0][2] ~^ image[17][8])} + {7'd0,(kernel[0][3] ~^ image[17][9])} + {7'd0,(kernel[0][4] ~^ image[17][10])} + {7'd0,(kernel[1][0] ~^ image[18][6])} + {7'd0,(kernel[1][1] ~^ image[18][7])} + {7'd0,(kernel[1][2] ~^ image[18][8])} + {7'd0,(kernel[1][3] ~^ image[18][9])} + {7'd0,(kernel[1][4] ~^ image[18][10])} + {7'd0,(kernel[2][0] ~^ image[19][6])} + {7'd0,(kernel[2][1] ~^ image[19][7])} + {7'd0,(kernel[2][2] ~^ image[19][8])} + {7'd0,(kernel[2][3] ~^ image[19][9])} + {7'd0,(kernel[2][4] ~^ image[19][10])} + {7'd0,(kernel[3][0] ~^ image[20][6])} + {7'd0,(kernel[3][1] ~^ image[20][7])} + {7'd0,(kernel[3][2] ~^ image[20][8])} + {7'd0,(kernel[3][3] ~^ image[20][9])} + {7'd0,(kernel[3][4] ~^ image[20][10])} + {7'd0,(kernel[4][0] ~^ image[21][6])} + {7'd0,(kernel[4][1] ~^ image[21][7])} + {7'd0,(kernel[4][2] ~^ image[21][8])} + {7'd0,(kernel[4][3] ~^ image[21][9])} + {7'd0,(kernel[4][4] ~^ image[21][10])};
assign out_fmap[17][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[17][7])} + {7'd0,(kernel[0][1] ~^ image[17][8])} + {7'd0,(kernel[0][2] ~^ image[17][9])} + {7'd0,(kernel[0][3] ~^ image[17][10])} + {7'd0,(kernel[0][4] ~^ image[17][11])} + {7'd0,(kernel[1][0] ~^ image[18][7])} + {7'd0,(kernel[1][1] ~^ image[18][8])} + {7'd0,(kernel[1][2] ~^ image[18][9])} + {7'd0,(kernel[1][3] ~^ image[18][10])} + {7'd0,(kernel[1][4] ~^ image[18][11])} + {7'd0,(kernel[2][0] ~^ image[19][7])} + {7'd0,(kernel[2][1] ~^ image[19][8])} + {7'd0,(kernel[2][2] ~^ image[19][9])} + {7'd0,(kernel[2][3] ~^ image[19][10])} + {7'd0,(kernel[2][4] ~^ image[19][11])} + {7'd0,(kernel[3][0] ~^ image[20][7])} + {7'd0,(kernel[3][1] ~^ image[20][8])} + {7'd0,(kernel[3][2] ~^ image[20][9])} + {7'd0,(kernel[3][3] ~^ image[20][10])} + {7'd0,(kernel[3][4] ~^ image[20][11])} + {7'd0,(kernel[4][0] ~^ image[21][7])} + {7'd0,(kernel[4][1] ~^ image[21][8])} + {7'd0,(kernel[4][2] ~^ image[21][9])} + {7'd0,(kernel[4][3] ~^ image[21][10])} + {7'd0,(kernel[4][4] ~^ image[21][11])};
assign out_fmap[17][8][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[17][8])} + {7'd0,(kernel[0][1] ~^ image[17][9])} + {7'd0,(kernel[0][2] ~^ image[17][10])} + {7'd0,(kernel[0][3] ~^ image[17][11])} + {7'd0,(kernel[0][4] ~^ image[17][12])} + {7'd0,(kernel[1][0] ~^ image[18][8])} + {7'd0,(kernel[1][1] ~^ image[18][9])} + {7'd0,(kernel[1][2] ~^ image[18][10])} + {7'd0,(kernel[1][3] ~^ image[18][11])} + {7'd0,(kernel[1][4] ~^ image[18][12])} + {7'd0,(kernel[2][0] ~^ image[19][8])} + {7'd0,(kernel[2][1] ~^ image[19][9])} + {7'd0,(kernel[2][2] ~^ image[19][10])} + {7'd0,(kernel[2][3] ~^ image[19][11])} + {7'd0,(kernel[2][4] ~^ image[19][12])} + {7'd0,(kernel[3][0] ~^ image[20][8])} + {7'd0,(kernel[3][1] ~^ image[20][9])} + {7'd0,(kernel[3][2] ~^ image[20][10])} + {7'd0,(kernel[3][3] ~^ image[20][11])} + {7'd0,(kernel[3][4] ~^ image[20][12])} + {7'd0,(kernel[4][0] ~^ image[21][8])} + {7'd0,(kernel[4][1] ~^ image[21][9])} + {7'd0,(kernel[4][2] ~^ image[21][10])} + {7'd0,(kernel[4][3] ~^ image[21][11])} + {7'd0,(kernel[4][4] ~^ image[21][12])};
assign out_fmap[17][9][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[17][9])} + {7'd0,(kernel[0][1] ~^ image[17][10])} + {7'd0,(kernel[0][2] ~^ image[17][11])} + {7'd0,(kernel[0][3] ~^ image[17][12])} + {7'd0,(kernel[0][4] ~^ image[17][13])} + {7'd0,(kernel[1][0] ~^ image[18][9])} + {7'd0,(kernel[1][1] ~^ image[18][10])} + {7'd0,(kernel[1][2] ~^ image[18][11])} + {7'd0,(kernel[1][3] ~^ image[18][12])} + {7'd0,(kernel[1][4] ~^ image[18][13])} + {7'd0,(kernel[2][0] ~^ image[19][9])} + {7'd0,(kernel[2][1] ~^ image[19][10])} + {7'd0,(kernel[2][2] ~^ image[19][11])} + {7'd0,(kernel[2][3] ~^ image[19][12])} + {7'd0,(kernel[2][4] ~^ image[19][13])} + {7'd0,(kernel[3][0] ~^ image[20][9])} + {7'd0,(kernel[3][1] ~^ image[20][10])} + {7'd0,(kernel[3][2] ~^ image[20][11])} + {7'd0,(kernel[3][3] ~^ image[20][12])} + {7'd0,(kernel[3][4] ~^ image[20][13])} + {7'd0,(kernel[4][0] ~^ image[21][9])} + {7'd0,(kernel[4][1] ~^ image[21][10])} + {7'd0,(kernel[4][2] ~^ image[21][11])} + {7'd0,(kernel[4][3] ~^ image[21][12])} + {7'd0,(kernel[4][4] ~^ image[21][13])};
assign out_fmap[17][10][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[17][10])} + {7'd0,(kernel[0][1] ~^ image[17][11])} + {7'd0,(kernel[0][2] ~^ image[17][12])} + {7'd0,(kernel[0][3] ~^ image[17][13])} + {7'd0,(kernel[0][4] ~^ image[17][14])} + {7'd0,(kernel[1][0] ~^ image[18][10])} + {7'd0,(kernel[1][1] ~^ image[18][11])} + {7'd0,(kernel[1][2] ~^ image[18][12])} + {7'd0,(kernel[1][3] ~^ image[18][13])} + {7'd0,(kernel[1][4] ~^ image[18][14])} + {7'd0,(kernel[2][0] ~^ image[19][10])} + {7'd0,(kernel[2][1] ~^ image[19][11])} + {7'd0,(kernel[2][2] ~^ image[19][12])} + {7'd0,(kernel[2][3] ~^ image[19][13])} + {7'd0,(kernel[2][4] ~^ image[19][14])} + {7'd0,(kernel[3][0] ~^ image[20][10])} + {7'd0,(kernel[3][1] ~^ image[20][11])} + {7'd0,(kernel[3][2] ~^ image[20][12])} + {7'd0,(kernel[3][3] ~^ image[20][13])} + {7'd0,(kernel[3][4] ~^ image[20][14])} + {7'd0,(kernel[4][0] ~^ image[21][10])} + {7'd0,(kernel[4][1] ~^ image[21][11])} + {7'd0,(kernel[4][2] ~^ image[21][12])} + {7'd0,(kernel[4][3] ~^ image[21][13])} + {7'd0,(kernel[4][4] ~^ image[21][14])};
assign out_fmap[17][11][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[17][11])} + {7'd0,(kernel[0][1] ~^ image[17][12])} + {7'd0,(kernel[0][2] ~^ image[17][13])} + {7'd0,(kernel[0][3] ~^ image[17][14])} + {7'd0,(kernel[0][4] ~^ image[17][15])} + {7'd0,(kernel[1][0] ~^ image[18][11])} + {7'd0,(kernel[1][1] ~^ image[18][12])} + {7'd0,(kernel[1][2] ~^ image[18][13])} + {7'd0,(kernel[1][3] ~^ image[18][14])} + {7'd0,(kernel[1][4] ~^ image[18][15])} + {7'd0,(kernel[2][0] ~^ image[19][11])} + {7'd0,(kernel[2][1] ~^ image[19][12])} + {7'd0,(kernel[2][2] ~^ image[19][13])} + {7'd0,(kernel[2][3] ~^ image[19][14])} + {7'd0,(kernel[2][4] ~^ image[19][15])} + {7'd0,(kernel[3][0] ~^ image[20][11])} + {7'd0,(kernel[3][1] ~^ image[20][12])} + {7'd0,(kernel[3][2] ~^ image[20][13])} + {7'd0,(kernel[3][3] ~^ image[20][14])} + {7'd0,(kernel[3][4] ~^ image[20][15])} + {7'd0,(kernel[4][0] ~^ image[21][11])} + {7'd0,(kernel[4][1] ~^ image[21][12])} + {7'd0,(kernel[4][2] ~^ image[21][13])} + {7'd0,(kernel[4][3] ~^ image[21][14])} + {7'd0,(kernel[4][4] ~^ image[21][15])};
assign out_fmap[17][12][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[17][12])} + {7'd0,(kernel[0][1] ~^ image[17][13])} + {7'd0,(kernel[0][2] ~^ image[17][14])} + {7'd0,(kernel[0][3] ~^ image[17][15])} + {7'd0,(kernel[0][4] ~^ image[17][16])} + {7'd0,(kernel[1][0] ~^ image[18][12])} + {7'd0,(kernel[1][1] ~^ image[18][13])} + {7'd0,(kernel[1][2] ~^ image[18][14])} + {7'd0,(kernel[1][3] ~^ image[18][15])} + {7'd0,(kernel[1][4] ~^ image[18][16])} + {7'd0,(kernel[2][0] ~^ image[19][12])} + {7'd0,(kernel[2][1] ~^ image[19][13])} + {7'd0,(kernel[2][2] ~^ image[19][14])} + {7'd0,(kernel[2][3] ~^ image[19][15])} + {7'd0,(kernel[2][4] ~^ image[19][16])} + {7'd0,(kernel[3][0] ~^ image[20][12])} + {7'd0,(kernel[3][1] ~^ image[20][13])} + {7'd0,(kernel[3][2] ~^ image[20][14])} + {7'd0,(kernel[3][3] ~^ image[20][15])} + {7'd0,(kernel[3][4] ~^ image[20][16])} + {7'd0,(kernel[4][0] ~^ image[21][12])} + {7'd0,(kernel[4][1] ~^ image[21][13])} + {7'd0,(kernel[4][2] ~^ image[21][14])} + {7'd0,(kernel[4][3] ~^ image[21][15])} + {7'd0,(kernel[4][4] ~^ image[21][16])};
assign out_fmap[17][13][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[17][13])} + {7'd0,(kernel[0][1] ~^ image[17][14])} + {7'd0,(kernel[0][2] ~^ image[17][15])} + {7'd0,(kernel[0][3] ~^ image[17][16])} + {7'd0,(kernel[0][4] ~^ image[17][17])} + {7'd0,(kernel[1][0] ~^ image[18][13])} + {7'd0,(kernel[1][1] ~^ image[18][14])} + {7'd0,(kernel[1][2] ~^ image[18][15])} + {7'd0,(kernel[1][3] ~^ image[18][16])} + {7'd0,(kernel[1][4] ~^ image[18][17])} + {7'd0,(kernel[2][0] ~^ image[19][13])} + {7'd0,(kernel[2][1] ~^ image[19][14])} + {7'd0,(kernel[2][2] ~^ image[19][15])} + {7'd0,(kernel[2][3] ~^ image[19][16])} + {7'd0,(kernel[2][4] ~^ image[19][17])} + {7'd0,(kernel[3][0] ~^ image[20][13])} + {7'd0,(kernel[3][1] ~^ image[20][14])} + {7'd0,(kernel[3][2] ~^ image[20][15])} + {7'd0,(kernel[3][3] ~^ image[20][16])} + {7'd0,(kernel[3][4] ~^ image[20][17])} + {7'd0,(kernel[4][0] ~^ image[21][13])} + {7'd0,(kernel[4][1] ~^ image[21][14])} + {7'd0,(kernel[4][2] ~^ image[21][15])} + {7'd0,(kernel[4][3] ~^ image[21][16])} + {7'd0,(kernel[4][4] ~^ image[21][17])};
assign out_fmap[17][14][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[17][14])} + {7'd0,(kernel[0][1] ~^ image[17][15])} + {7'd0,(kernel[0][2] ~^ image[17][16])} + {7'd0,(kernel[0][3] ~^ image[17][17])} + {7'd0,(kernel[0][4] ~^ image[17][18])} + {7'd0,(kernel[1][0] ~^ image[18][14])} + {7'd0,(kernel[1][1] ~^ image[18][15])} + {7'd0,(kernel[1][2] ~^ image[18][16])} + {7'd0,(kernel[1][3] ~^ image[18][17])} + {7'd0,(kernel[1][4] ~^ image[18][18])} + {7'd0,(kernel[2][0] ~^ image[19][14])} + {7'd0,(kernel[2][1] ~^ image[19][15])} + {7'd0,(kernel[2][2] ~^ image[19][16])} + {7'd0,(kernel[2][3] ~^ image[19][17])} + {7'd0,(kernel[2][4] ~^ image[19][18])} + {7'd0,(kernel[3][0] ~^ image[20][14])} + {7'd0,(kernel[3][1] ~^ image[20][15])} + {7'd0,(kernel[3][2] ~^ image[20][16])} + {7'd0,(kernel[3][3] ~^ image[20][17])} + {7'd0,(kernel[3][4] ~^ image[20][18])} + {7'd0,(kernel[4][0] ~^ image[21][14])} + {7'd0,(kernel[4][1] ~^ image[21][15])} + {7'd0,(kernel[4][2] ~^ image[21][16])} + {7'd0,(kernel[4][3] ~^ image[21][17])} + {7'd0,(kernel[4][4] ~^ image[21][18])};
assign out_fmap[17][15][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[17][15])} + {7'd0,(kernel[0][1] ~^ image[17][16])} + {7'd0,(kernel[0][2] ~^ image[17][17])} + {7'd0,(kernel[0][3] ~^ image[17][18])} + {7'd0,(kernel[0][4] ~^ image[17][19])} + {7'd0,(kernel[1][0] ~^ image[18][15])} + {7'd0,(kernel[1][1] ~^ image[18][16])} + {7'd0,(kernel[1][2] ~^ image[18][17])} + {7'd0,(kernel[1][3] ~^ image[18][18])} + {7'd0,(kernel[1][4] ~^ image[18][19])} + {7'd0,(kernel[2][0] ~^ image[19][15])} + {7'd0,(kernel[2][1] ~^ image[19][16])} + {7'd0,(kernel[2][2] ~^ image[19][17])} + {7'd0,(kernel[2][3] ~^ image[19][18])} + {7'd0,(kernel[2][4] ~^ image[19][19])} + {7'd0,(kernel[3][0] ~^ image[20][15])} + {7'd0,(kernel[3][1] ~^ image[20][16])} + {7'd0,(kernel[3][2] ~^ image[20][17])} + {7'd0,(kernel[3][3] ~^ image[20][18])} + {7'd0,(kernel[3][4] ~^ image[20][19])} + {7'd0,(kernel[4][0] ~^ image[21][15])} + {7'd0,(kernel[4][1] ~^ image[21][16])} + {7'd0,(kernel[4][2] ~^ image[21][17])} + {7'd0,(kernel[4][3] ~^ image[21][18])} + {7'd0,(kernel[4][4] ~^ image[21][19])};
assign out_fmap[17][16][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[17][16])} + {7'd0,(kernel[0][1] ~^ image[17][17])} + {7'd0,(kernel[0][2] ~^ image[17][18])} + {7'd0,(kernel[0][3] ~^ image[17][19])} + {7'd0,(kernel[0][4] ~^ image[17][20])} + {7'd0,(kernel[1][0] ~^ image[18][16])} + {7'd0,(kernel[1][1] ~^ image[18][17])} + {7'd0,(kernel[1][2] ~^ image[18][18])} + {7'd0,(kernel[1][3] ~^ image[18][19])} + {7'd0,(kernel[1][4] ~^ image[18][20])} + {7'd0,(kernel[2][0] ~^ image[19][16])} + {7'd0,(kernel[2][1] ~^ image[19][17])} + {7'd0,(kernel[2][2] ~^ image[19][18])} + {7'd0,(kernel[2][3] ~^ image[19][19])} + {7'd0,(kernel[2][4] ~^ image[19][20])} + {7'd0,(kernel[3][0] ~^ image[20][16])} + {7'd0,(kernel[3][1] ~^ image[20][17])} + {7'd0,(kernel[3][2] ~^ image[20][18])} + {7'd0,(kernel[3][3] ~^ image[20][19])} + {7'd0,(kernel[3][4] ~^ image[20][20])} + {7'd0,(kernel[4][0] ~^ image[21][16])} + {7'd0,(kernel[4][1] ~^ image[21][17])} + {7'd0,(kernel[4][2] ~^ image[21][18])} + {7'd0,(kernel[4][3] ~^ image[21][19])} + {7'd0,(kernel[4][4] ~^ image[21][20])};
assign out_fmap[17][17][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[17][17])} + {7'd0,(kernel[0][1] ~^ image[17][18])} + {7'd0,(kernel[0][2] ~^ image[17][19])} + {7'd0,(kernel[0][3] ~^ image[17][20])} + {7'd0,(kernel[0][4] ~^ image[17][21])} + {7'd0,(kernel[1][0] ~^ image[18][17])} + {7'd0,(kernel[1][1] ~^ image[18][18])} + {7'd0,(kernel[1][2] ~^ image[18][19])} + {7'd0,(kernel[1][3] ~^ image[18][20])} + {7'd0,(kernel[1][4] ~^ image[18][21])} + {7'd0,(kernel[2][0] ~^ image[19][17])} + {7'd0,(kernel[2][1] ~^ image[19][18])} + {7'd0,(kernel[2][2] ~^ image[19][19])} + {7'd0,(kernel[2][3] ~^ image[19][20])} + {7'd0,(kernel[2][4] ~^ image[19][21])} + {7'd0,(kernel[3][0] ~^ image[20][17])} + {7'd0,(kernel[3][1] ~^ image[20][18])} + {7'd0,(kernel[3][2] ~^ image[20][19])} + {7'd0,(kernel[3][3] ~^ image[20][20])} + {7'd0,(kernel[3][4] ~^ image[20][21])} + {7'd0,(kernel[4][0] ~^ image[21][17])} + {7'd0,(kernel[4][1] ~^ image[21][18])} + {7'd0,(kernel[4][2] ~^ image[21][19])} + {7'd0,(kernel[4][3] ~^ image[21][20])} + {7'd0,(kernel[4][4] ~^ image[21][21])};
assign out_fmap[17][18][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[17][18])} + {7'd0,(kernel[0][1] ~^ image[17][19])} + {7'd0,(kernel[0][2] ~^ image[17][20])} + {7'd0,(kernel[0][3] ~^ image[17][21])} + {7'd0,(kernel[0][4] ~^ image[17][22])} + {7'd0,(kernel[1][0] ~^ image[18][18])} + {7'd0,(kernel[1][1] ~^ image[18][19])} + {7'd0,(kernel[1][2] ~^ image[18][20])} + {7'd0,(kernel[1][3] ~^ image[18][21])} + {7'd0,(kernel[1][4] ~^ image[18][22])} + {7'd0,(kernel[2][0] ~^ image[19][18])} + {7'd0,(kernel[2][1] ~^ image[19][19])} + {7'd0,(kernel[2][2] ~^ image[19][20])} + {7'd0,(kernel[2][3] ~^ image[19][21])} + {7'd0,(kernel[2][4] ~^ image[19][22])} + {7'd0,(kernel[3][0] ~^ image[20][18])} + {7'd0,(kernel[3][1] ~^ image[20][19])} + {7'd0,(kernel[3][2] ~^ image[20][20])} + {7'd0,(kernel[3][3] ~^ image[20][21])} + {7'd0,(kernel[3][4] ~^ image[20][22])} + {7'd0,(kernel[4][0] ~^ image[21][18])} + {7'd0,(kernel[4][1] ~^ image[21][19])} + {7'd0,(kernel[4][2] ~^ image[21][20])} + {7'd0,(kernel[4][3] ~^ image[21][21])} + {7'd0,(kernel[4][4] ~^ image[21][22])};
assign out_fmap[17][19][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[17][19])} + {7'd0,(kernel[0][1] ~^ image[17][20])} + {7'd0,(kernel[0][2] ~^ image[17][21])} + {7'd0,(kernel[0][3] ~^ image[17][22])} + {7'd0,(kernel[0][4] ~^ image[17][23])} + {7'd0,(kernel[1][0] ~^ image[18][19])} + {7'd0,(kernel[1][1] ~^ image[18][20])} + {7'd0,(kernel[1][2] ~^ image[18][21])} + {7'd0,(kernel[1][3] ~^ image[18][22])} + {7'd0,(kernel[1][4] ~^ image[18][23])} + {7'd0,(kernel[2][0] ~^ image[19][19])} + {7'd0,(kernel[2][1] ~^ image[19][20])} + {7'd0,(kernel[2][2] ~^ image[19][21])} + {7'd0,(kernel[2][3] ~^ image[19][22])} + {7'd0,(kernel[2][4] ~^ image[19][23])} + {7'd0,(kernel[3][0] ~^ image[20][19])} + {7'd0,(kernel[3][1] ~^ image[20][20])} + {7'd0,(kernel[3][2] ~^ image[20][21])} + {7'd0,(kernel[3][3] ~^ image[20][22])} + {7'd0,(kernel[3][4] ~^ image[20][23])} + {7'd0,(kernel[4][0] ~^ image[21][19])} + {7'd0,(kernel[4][1] ~^ image[21][20])} + {7'd0,(kernel[4][2] ~^ image[21][21])} + {7'd0,(kernel[4][3] ~^ image[21][22])} + {7'd0,(kernel[4][4] ~^ image[21][23])};
assign out_fmap[17][20][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[17][20])} + {7'd0,(kernel[0][1] ~^ image[17][21])} + {7'd0,(kernel[0][2] ~^ image[17][22])} + {7'd0,(kernel[0][3] ~^ image[17][23])} + {7'd0,(kernel[0][4] ~^ image[17][24])} + {7'd0,(kernel[1][0] ~^ image[18][20])} + {7'd0,(kernel[1][1] ~^ image[18][21])} + {7'd0,(kernel[1][2] ~^ image[18][22])} + {7'd0,(kernel[1][3] ~^ image[18][23])} + {7'd0,(kernel[1][4] ~^ image[18][24])} + {7'd0,(kernel[2][0] ~^ image[19][20])} + {7'd0,(kernel[2][1] ~^ image[19][21])} + {7'd0,(kernel[2][2] ~^ image[19][22])} + {7'd0,(kernel[2][3] ~^ image[19][23])} + {7'd0,(kernel[2][4] ~^ image[19][24])} + {7'd0,(kernel[3][0] ~^ image[20][20])} + {7'd0,(kernel[3][1] ~^ image[20][21])} + {7'd0,(kernel[3][2] ~^ image[20][22])} + {7'd0,(kernel[3][3] ~^ image[20][23])} + {7'd0,(kernel[3][4] ~^ image[20][24])} + {7'd0,(kernel[4][0] ~^ image[21][20])} + {7'd0,(kernel[4][1] ~^ image[21][21])} + {7'd0,(kernel[4][2] ~^ image[21][22])} + {7'd0,(kernel[4][3] ~^ image[21][23])} + {7'd0,(kernel[4][4] ~^ image[21][24])};
assign out_fmap[17][21][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[17][21])} + {7'd0,(kernel[0][1] ~^ image[17][22])} + {7'd0,(kernel[0][2] ~^ image[17][23])} + {7'd0,(kernel[0][3] ~^ image[17][24])} + {7'd0,(kernel[0][4] ~^ image[17][25])} + {7'd0,(kernel[1][0] ~^ image[18][21])} + {7'd0,(kernel[1][1] ~^ image[18][22])} + {7'd0,(kernel[1][2] ~^ image[18][23])} + {7'd0,(kernel[1][3] ~^ image[18][24])} + {7'd0,(kernel[1][4] ~^ image[18][25])} + {7'd0,(kernel[2][0] ~^ image[19][21])} + {7'd0,(kernel[2][1] ~^ image[19][22])} + {7'd0,(kernel[2][2] ~^ image[19][23])} + {7'd0,(kernel[2][3] ~^ image[19][24])} + {7'd0,(kernel[2][4] ~^ image[19][25])} + {7'd0,(kernel[3][0] ~^ image[20][21])} + {7'd0,(kernel[3][1] ~^ image[20][22])} + {7'd0,(kernel[3][2] ~^ image[20][23])} + {7'd0,(kernel[3][3] ~^ image[20][24])} + {7'd0,(kernel[3][4] ~^ image[20][25])} + {7'd0,(kernel[4][0] ~^ image[21][21])} + {7'd0,(kernel[4][1] ~^ image[21][22])} + {7'd0,(kernel[4][2] ~^ image[21][23])} + {7'd0,(kernel[4][3] ~^ image[21][24])} + {7'd0,(kernel[4][4] ~^ image[21][25])};
assign out_fmap[17][22][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[17][22])} + {7'd0,(kernel[0][1] ~^ image[17][23])} + {7'd0,(kernel[0][2] ~^ image[17][24])} + {7'd0,(kernel[0][3] ~^ image[17][25])} + {7'd0,(kernel[0][4] ~^ image[17][26])} + {7'd0,(kernel[1][0] ~^ image[18][22])} + {7'd0,(kernel[1][1] ~^ image[18][23])} + {7'd0,(kernel[1][2] ~^ image[18][24])} + {7'd0,(kernel[1][3] ~^ image[18][25])} + {7'd0,(kernel[1][4] ~^ image[18][26])} + {7'd0,(kernel[2][0] ~^ image[19][22])} + {7'd0,(kernel[2][1] ~^ image[19][23])} + {7'd0,(kernel[2][2] ~^ image[19][24])} + {7'd0,(kernel[2][3] ~^ image[19][25])} + {7'd0,(kernel[2][4] ~^ image[19][26])} + {7'd0,(kernel[3][0] ~^ image[20][22])} + {7'd0,(kernel[3][1] ~^ image[20][23])} + {7'd0,(kernel[3][2] ~^ image[20][24])} + {7'd0,(kernel[3][3] ~^ image[20][25])} + {7'd0,(kernel[3][4] ~^ image[20][26])} + {7'd0,(kernel[4][0] ~^ image[21][22])} + {7'd0,(kernel[4][1] ~^ image[21][23])} + {7'd0,(kernel[4][2] ~^ image[21][24])} + {7'd0,(kernel[4][3] ~^ image[21][25])} + {7'd0,(kernel[4][4] ~^ image[21][26])};
assign out_fmap[17][23][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[17][23])} + {7'd0,(kernel[0][1] ~^ image[17][24])} + {7'd0,(kernel[0][2] ~^ image[17][25])} + {7'd0,(kernel[0][3] ~^ image[17][26])} + {7'd0,(kernel[0][4] ~^ image[17][27])} + {7'd0,(kernel[1][0] ~^ image[18][23])} + {7'd0,(kernel[1][1] ~^ image[18][24])} + {7'd0,(kernel[1][2] ~^ image[18][25])} + {7'd0,(kernel[1][3] ~^ image[18][26])} + {7'd0,(kernel[1][4] ~^ image[18][27])} + {7'd0,(kernel[2][0] ~^ image[19][23])} + {7'd0,(kernel[2][1] ~^ image[19][24])} + {7'd0,(kernel[2][2] ~^ image[19][25])} + {7'd0,(kernel[2][3] ~^ image[19][26])} + {7'd0,(kernel[2][4] ~^ image[19][27])} + {7'd0,(kernel[3][0] ~^ image[20][23])} + {7'd0,(kernel[3][1] ~^ image[20][24])} + {7'd0,(kernel[3][2] ~^ image[20][25])} + {7'd0,(kernel[3][3] ~^ image[20][26])} + {7'd0,(kernel[3][4] ~^ image[20][27])} + {7'd0,(kernel[4][0] ~^ image[21][23])} + {7'd0,(kernel[4][1] ~^ image[21][24])} + {7'd0,(kernel[4][2] ~^ image[21][25])} + {7'd0,(kernel[4][3] ~^ image[21][26])} + {7'd0,(kernel[4][4] ~^ image[21][27])};
assign out_fmap[18][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[18][0])} + {7'd0,(kernel[0][1] ~^ image[18][1])} + {7'd0,(kernel[0][2] ~^ image[18][2])} + {7'd0,(kernel[0][3] ~^ image[18][3])} + {7'd0,(kernel[0][4] ~^ image[18][4])} + {7'd0,(kernel[1][0] ~^ image[19][0])} + {7'd0,(kernel[1][1] ~^ image[19][1])} + {7'd0,(kernel[1][2] ~^ image[19][2])} + {7'd0,(kernel[1][3] ~^ image[19][3])} + {7'd0,(kernel[1][4] ~^ image[19][4])} + {7'd0,(kernel[2][0] ~^ image[20][0])} + {7'd0,(kernel[2][1] ~^ image[20][1])} + {7'd0,(kernel[2][2] ~^ image[20][2])} + {7'd0,(kernel[2][3] ~^ image[20][3])} + {7'd0,(kernel[2][4] ~^ image[20][4])} + {7'd0,(kernel[3][0] ~^ image[21][0])} + {7'd0,(kernel[3][1] ~^ image[21][1])} + {7'd0,(kernel[3][2] ~^ image[21][2])} + {7'd0,(kernel[3][3] ~^ image[21][3])} + {7'd0,(kernel[3][4] ~^ image[21][4])} + {7'd0,(kernel[4][0] ~^ image[22][0])} + {7'd0,(kernel[4][1] ~^ image[22][1])} + {7'd0,(kernel[4][2] ~^ image[22][2])} + {7'd0,(kernel[4][3] ~^ image[22][3])} + {7'd0,(kernel[4][4] ~^ image[22][4])};
assign out_fmap[18][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[18][1])} + {7'd0,(kernel[0][1] ~^ image[18][2])} + {7'd0,(kernel[0][2] ~^ image[18][3])} + {7'd0,(kernel[0][3] ~^ image[18][4])} + {7'd0,(kernel[0][4] ~^ image[18][5])} + {7'd0,(kernel[1][0] ~^ image[19][1])} + {7'd0,(kernel[1][1] ~^ image[19][2])} + {7'd0,(kernel[1][2] ~^ image[19][3])} + {7'd0,(kernel[1][3] ~^ image[19][4])} + {7'd0,(kernel[1][4] ~^ image[19][5])} + {7'd0,(kernel[2][0] ~^ image[20][1])} + {7'd0,(kernel[2][1] ~^ image[20][2])} + {7'd0,(kernel[2][2] ~^ image[20][3])} + {7'd0,(kernel[2][3] ~^ image[20][4])} + {7'd0,(kernel[2][4] ~^ image[20][5])} + {7'd0,(kernel[3][0] ~^ image[21][1])} + {7'd0,(kernel[3][1] ~^ image[21][2])} + {7'd0,(kernel[3][2] ~^ image[21][3])} + {7'd0,(kernel[3][3] ~^ image[21][4])} + {7'd0,(kernel[3][4] ~^ image[21][5])} + {7'd0,(kernel[4][0] ~^ image[22][1])} + {7'd0,(kernel[4][1] ~^ image[22][2])} + {7'd0,(kernel[4][2] ~^ image[22][3])} + {7'd0,(kernel[4][3] ~^ image[22][4])} + {7'd0,(kernel[4][4] ~^ image[22][5])};
assign out_fmap[18][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[18][2])} + {7'd0,(kernel[0][1] ~^ image[18][3])} + {7'd0,(kernel[0][2] ~^ image[18][4])} + {7'd0,(kernel[0][3] ~^ image[18][5])} + {7'd0,(kernel[0][4] ~^ image[18][6])} + {7'd0,(kernel[1][0] ~^ image[19][2])} + {7'd0,(kernel[1][1] ~^ image[19][3])} + {7'd0,(kernel[1][2] ~^ image[19][4])} + {7'd0,(kernel[1][3] ~^ image[19][5])} + {7'd0,(kernel[1][4] ~^ image[19][6])} + {7'd0,(kernel[2][0] ~^ image[20][2])} + {7'd0,(kernel[2][1] ~^ image[20][3])} + {7'd0,(kernel[2][2] ~^ image[20][4])} + {7'd0,(kernel[2][3] ~^ image[20][5])} + {7'd0,(kernel[2][4] ~^ image[20][6])} + {7'd0,(kernel[3][0] ~^ image[21][2])} + {7'd0,(kernel[3][1] ~^ image[21][3])} + {7'd0,(kernel[3][2] ~^ image[21][4])} + {7'd0,(kernel[3][3] ~^ image[21][5])} + {7'd0,(kernel[3][4] ~^ image[21][6])} + {7'd0,(kernel[4][0] ~^ image[22][2])} + {7'd0,(kernel[4][1] ~^ image[22][3])} + {7'd0,(kernel[4][2] ~^ image[22][4])} + {7'd0,(kernel[4][3] ~^ image[22][5])} + {7'd0,(kernel[4][4] ~^ image[22][6])};
assign out_fmap[18][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[18][3])} + {7'd0,(kernel[0][1] ~^ image[18][4])} + {7'd0,(kernel[0][2] ~^ image[18][5])} + {7'd0,(kernel[0][3] ~^ image[18][6])} + {7'd0,(kernel[0][4] ~^ image[18][7])} + {7'd0,(kernel[1][0] ~^ image[19][3])} + {7'd0,(kernel[1][1] ~^ image[19][4])} + {7'd0,(kernel[1][2] ~^ image[19][5])} + {7'd0,(kernel[1][3] ~^ image[19][6])} + {7'd0,(kernel[1][4] ~^ image[19][7])} + {7'd0,(kernel[2][0] ~^ image[20][3])} + {7'd0,(kernel[2][1] ~^ image[20][4])} + {7'd0,(kernel[2][2] ~^ image[20][5])} + {7'd0,(kernel[2][3] ~^ image[20][6])} + {7'd0,(kernel[2][4] ~^ image[20][7])} + {7'd0,(kernel[3][0] ~^ image[21][3])} + {7'd0,(kernel[3][1] ~^ image[21][4])} + {7'd0,(kernel[3][2] ~^ image[21][5])} + {7'd0,(kernel[3][3] ~^ image[21][6])} + {7'd0,(kernel[3][4] ~^ image[21][7])} + {7'd0,(kernel[4][0] ~^ image[22][3])} + {7'd0,(kernel[4][1] ~^ image[22][4])} + {7'd0,(kernel[4][2] ~^ image[22][5])} + {7'd0,(kernel[4][3] ~^ image[22][6])} + {7'd0,(kernel[4][4] ~^ image[22][7])};
assign out_fmap[18][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[18][4])} + {7'd0,(kernel[0][1] ~^ image[18][5])} + {7'd0,(kernel[0][2] ~^ image[18][6])} + {7'd0,(kernel[0][3] ~^ image[18][7])} + {7'd0,(kernel[0][4] ~^ image[18][8])} + {7'd0,(kernel[1][0] ~^ image[19][4])} + {7'd0,(kernel[1][1] ~^ image[19][5])} + {7'd0,(kernel[1][2] ~^ image[19][6])} + {7'd0,(kernel[1][3] ~^ image[19][7])} + {7'd0,(kernel[1][4] ~^ image[19][8])} + {7'd0,(kernel[2][0] ~^ image[20][4])} + {7'd0,(kernel[2][1] ~^ image[20][5])} + {7'd0,(kernel[2][2] ~^ image[20][6])} + {7'd0,(kernel[2][3] ~^ image[20][7])} + {7'd0,(kernel[2][4] ~^ image[20][8])} + {7'd0,(kernel[3][0] ~^ image[21][4])} + {7'd0,(kernel[3][1] ~^ image[21][5])} + {7'd0,(kernel[3][2] ~^ image[21][6])} + {7'd0,(kernel[3][3] ~^ image[21][7])} + {7'd0,(kernel[3][4] ~^ image[21][8])} + {7'd0,(kernel[4][0] ~^ image[22][4])} + {7'd0,(kernel[4][1] ~^ image[22][5])} + {7'd0,(kernel[4][2] ~^ image[22][6])} + {7'd0,(kernel[4][3] ~^ image[22][7])} + {7'd0,(kernel[4][4] ~^ image[22][8])};
assign out_fmap[18][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[18][5])} + {7'd0,(kernel[0][1] ~^ image[18][6])} + {7'd0,(kernel[0][2] ~^ image[18][7])} + {7'd0,(kernel[0][3] ~^ image[18][8])} + {7'd0,(kernel[0][4] ~^ image[18][9])} + {7'd0,(kernel[1][0] ~^ image[19][5])} + {7'd0,(kernel[1][1] ~^ image[19][6])} + {7'd0,(kernel[1][2] ~^ image[19][7])} + {7'd0,(kernel[1][3] ~^ image[19][8])} + {7'd0,(kernel[1][4] ~^ image[19][9])} + {7'd0,(kernel[2][0] ~^ image[20][5])} + {7'd0,(kernel[2][1] ~^ image[20][6])} + {7'd0,(kernel[2][2] ~^ image[20][7])} + {7'd0,(kernel[2][3] ~^ image[20][8])} + {7'd0,(kernel[2][4] ~^ image[20][9])} + {7'd0,(kernel[3][0] ~^ image[21][5])} + {7'd0,(kernel[3][1] ~^ image[21][6])} + {7'd0,(kernel[3][2] ~^ image[21][7])} + {7'd0,(kernel[3][3] ~^ image[21][8])} + {7'd0,(kernel[3][4] ~^ image[21][9])} + {7'd0,(kernel[4][0] ~^ image[22][5])} + {7'd0,(kernel[4][1] ~^ image[22][6])} + {7'd0,(kernel[4][2] ~^ image[22][7])} + {7'd0,(kernel[4][3] ~^ image[22][8])} + {7'd0,(kernel[4][4] ~^ image[22][9])};
assign out_fmap[18][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[18][6])} + {7'd0,(kernel[0][1] ~^ image[18][7])} + {7'd0,(kernel[0][2] ~^ image[18][8])} + {7'd0,(kernel[0][3] ~^ image[18][9])} + {7'd0,(kernel[0][4] ~^ image[18][10])} + {7'd0,(kernel[1][0] ~^ image[19][6])} + {7'd0,(kernel[1][1] ~^ image[19][7])} + {7'd0,(kernel[1][2] ~^ image[19][8])} + {7'd0,(kernel[1][3] ~^ image[19][9])} + {7'd0,(kernel[1][4] ~^ image[19][10])} + {7'd0,(kernel[2][0] ~^ image[20][6])} + {7'd0,(kernel[2][1] ~^ image[20][7])} + {7'd0,(kernel[2][2] ~^ image[20][8])} + {7'd0,(kernel[2][3] ~^ image[20][9])} + {7'd0,(kernel[2][4] ~^ image[20][10])} + {7'd0,(kernel[3][0] ~^ image[21][6])} + {7'd0,(kernel[3][1] ~^ image[21][7])} + {7'd0,(kernel[3][2] ~^ image[21][8])} + {7'd0,(kernel[3][3] ~^ image[21][9])} + {7'd0,(kernel[3][4] ~^ image[21][10])} + {7'd0,(kernel[4][0] ~^ image[22][6])} + {7'd0,(kernel[4][1] ~^ image[22][7])} + {7'd0,(kernel[4][2] ~^ image[22][8])} + {7'd0,(kernel[4][3] ~^ image[22][9])} + {7'd0,(kernel[4][4] ~^ image[22][10])};
assign out_fmap[18][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[18][7])} + {7'd0,(kernel[0][1] ~^ image[18][8])} + {7'd0,(kernel[0][2] ~^ image[18][9])} + {7'd0,(kernel[0][3] ~^ image[18][10])} + {7'd0,(kernel[0][4] ~^ image[18][11])} + {7'd0,(kernel[1][0] ~^ image[19][7])} + {7'd0,(kernel[1][1] ~^ image[19][8])} + {7'd0,(kernel[1][2] ~^ image[19][9])} + {7'd0,(kernel[1][3] ~^ image[19][10])} + {7'd0,(kernel[1][4] ~^ image[19][11])} + {7'd0,(kernel[2][0] ~^ image[20][7])} + {7'd0,(kernel[2][1] ~^ image[20][8])} + {7'd0,(kernel[2][2] ~^ image[20][9])} + {7'd0,(kernel[2][3] ~^ image[20][10])} + {7'd0,(kernel[2][4] ~^ image[20][11])} + {7'd0,(kernel[3][0] ~^ image[21][7])} + {7'd0,(kernel[3][1] ~^ image[21][8])} + {7'd0,(kernel[3][2] ~^ image[21][9])} + {7'd0,(kernel[3][3] ~^ image[21][10])} + {7'd0,(kernel[3][4] ~^ image[21][11])} + {7'd0,(kernel[4][0] ~^ image[22][7])} + {7'd0,(kernel[4][1] ~^ image[22][8])} + {7'd0,(kernel[4][2] ~^ image[22][9])} + {7'd0,(kernel[4][3] ~^ image[22][10])} + {7'd0,(kernel[4][4] ~^ image[22][11])};
assign out_fmap[18][8][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[18][8])} + {7'd0,(kernel[0][1] ~^ image[18][9])} + {7'd0,(kernel[0][2] ~^ image[18][10])} + {7'd0,(kernel[0][3] ~^ image[18][11])} + {7'd0,(kernel[0][4] ~^ image[18][12])} + {7'd0,(kernel[1][0] ~^ image[19][8])} + {7'd0,(kernel[1][1] ~^ image[19][9])} + {7'd0,(kernel[1][2] ~^ image[19][10])} + {7'd0,(kernel[1][3] ~^ image[19][11])} + {7'd0,(kernel[1][4] ~^ image[19][12])} + {7'd0,(kernel[2][0] ~^ image[20][8])} + {7'd0,(kernel[2][1] ~^ image[20][9])} + {7'd0,(kernel[2][2] ~^ image[20][10])} + {7'd0,(kernel[2][3] ~^ image[20][11])} + {7'd0,(kernel[2][4] ~^ image[20][12])} + {7'd0,(kernel[3][0] ~^ image[21][8])} + {7'd0,(kernel[3][1] ~^ image[21][9])} + {7'd0,(kernel[3][2] ~^ image[21][10])} + {7'd0,(kernel[3][3] ~^ image[21][11])} + {7'd0,(kernel[3][4] ~^ image[21][12])} + {7'd0,(kernel[4][0] ~^ image[22][8])} + {7'd0,(kernel[4][1] ~^ image[22][9])} + {7'd0,(kernel[4][2] ~^ image[22][10])} + {7'd0,(kernel[4][3] ~^ image[22][11])} + {7'd0,(kernel[4][4] ~^ image[22][12])};
assign out_fmap[18][9][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[18][9])} + {7'd0,(kernel[0][1] ~^ image[18][10])} + {7'd0,(kernel[0][2] ~^ image[18][11])} + {7'd0,(kernel[0][3] ~^ image[18][12])} + {7'd0,(kernel[0][4] ~^ image[18][13])} + {7'd0,(kernel[1][0] ~^ image[19][9])} + {7'd0,(kernel[1][1] ~^ image[19][10])} + {7'd0,(kernel[1][2] ~^ image[19][11])} + {7'd0,(kernel[1][3] ~^ image[19][12])} + {7'd0,(kernel[1][4] ~^ image[19][13])} + {7'd0,(kernel[2][0] ~^ image[20][9])} + {7'd0,(kernel[2][1] ~^ image[20][10])} + {7'd0,(kernel[2][2] ~^ image[20][11])} + {7'd0,(kernel[2][3] ~^ image[20][12])} + {7'd0,(kernel[2][4] ~^ image[20][13])} + {7'd0,(kernel[3][0] ~^ image[21][9])} + {7'd0,(kernel[3][1] ~^ image[21][10])} + {7'd0,(kernel[3][2] ~^ image[21][11])} + {7'd0,(kernel[3][3] ~^ image[21][12])} + {7'd0,(kernel[3][4] ~^ image[21][13])} + {7'd0,(kernel[4][0] ~^ image[22][9])} + {7'd0,(kernel[4][1] ~^ image[22][10])} + {7'd0,(kernel[4][2] ~^ image[22][11])} + {7'd0,(kernel[4][3] ~^ image[22][12])} + {7'd0,(kernel[4][4] ~^ image[22][13])};
assign out_fmap[18][10][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[18][10])} + {7'd0,(kernel[0][1] ~^ image[18][11])} + {7'd0,(kernel[0][2] ~^ image[18][12])} + {7'd0,(kernel[0][3] ~^ image[18][13])} + {7'd0,(kernel[0][4] ~^ image[18][14])} + {7'd0,(kernel[1][0] ~^ image[19][10])} + {7'd0,(kernel[1][1] ~^ image[19][11])} + {7'd0,(kernel[1][2] ~^ image[19][12])} + {7'd0,(kernel[1][3] ~^ image[19][13])} + {7'd0,(kernel[1][4] ~^ image[19][14])} + {7'd0,(kernel[2][0] ~^ image[20][10])} + {7'd0,(kernel[2][1] ~^ image[20][11])} + {7'd0,(kernel[2][2] ~^ image[20][12])} + {7'd0,(kernel[2][3] ~^ image[20][13])} + {7'd0,(kernel[2][4] ~^ image[20][14])} + {7'd0,(kernel[3][0] ~^ image[21][10])} + {7'd0,(kernel[3][1] ~^ image[21][11])} + {7'd0,(kernel[3][2] ~^ image[21][12])} + {7'd0,(kernel[3][3] ~^ image[21][13])} + {7'd0,(kernel[3][4] ~^ image[21][14])} + {7'd0,(kernel[4][0] ~^ image[22][10])} + {7'd0,(kernel[4][1] ~^ image[22][11])} + {7'd0,(kernel[4][2] ~^ image[22][12])} + {7'd0,(kernel[4][3] ~^ image[22][13])} + {7'd0,(kernel[4][4] ~^ image[22][14])};
assign out_fmap[18][11][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[18][11])} + {7'd0,(kernel[0][1] ~^ image[18][12])} + {7'd0,(kernel[0][2] ~^ image[18][13])} + {7'd0,(kernel[0][3] ~^ image[18][14])} + {7'd0,(kernel[0][4] ~^ image[18][15])} + {7'd0,(kernel[1][0] ~^ image[19][11])} + {7'd0,(kernel[1][1] ~^ image[19][12])} + {7'd0,(kernel[1][2] ~^ image[19][13])} + {7'd0,(kernel[1][3] ~^ image[19][14])} + {7'd0,(kernel[1][4] ~^ image[19][15])} + {7'd0,(kernel[2][0] ~^ image[20][11])} + {7'd0,(kernel[2][1] ~^ image[20][12])} + {7'd0,(kernel[2][2] ~^ image[20][13])} + {7'd0,(kernel[2][3] ~^ image[20][14])} + {7'd0,(kernel[2][4] ~^ image[20][15])} + {7'd0,(kernel[3][0] ~^ image[21][11])} + {7'd0,(kernel[3][1] ~^ image[21][12])} + {7'd0,(kernel[3][2] ~^ image[21][13])} + {7'd0,(kernel[3][3] ~^ image[21][14])} + {7'd0,(kernel[3][4] ~^ image[21][15])} + {7'd0,(kernel[4][0] ~^ image[22][11])} + {7'd0,(kernel[4][1] ~^ image[22][12])} + {7'd0,(kernel[4][2] ~^ image[22][13])} + {7'd0,(kernel[4][3] ~^ image[22][14])} + {7'd0,(kernel[4][4] ~^ image[22][15])};
assign out_fmap[18][12][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[18][12])} + {7'd0,(kernel[0][1] ~^ image[18][13])} + {7'd0,(kernel[0][2] ~^ image[18][14])} + {7'd0,(kernel[0][3] ~^ image[18][15])} + {7'd0,(kernel[0][4] ~^ image[18][16])} + {7'd0,(kernel[1][0] ~^ image[19][12])} + {7'd0,(kernel[1][1] ~^ image[19][13])} + {7'd0,(kernel[1][2] ~^ image[19][14])} + {7'd0,(kernel[1][3] ~^ image[19][15])} + {7'd0,(kernel[1][4] ~^ image[19][16])} + {7'd0,(kernel[2][0] ~^ image[20][12])} + {7'd0,(kernel[2][1] ~^ image[20][13])} + {7'd0,(kernel[2][2] ~^ image[20][14])} + {7'd0,(kernel[2][3] ~^ image[20][15])} + {7'd0,(kernel[2][4] ~^ image[20][16])} + {7'd0,(kernel[3][0] ~^ image[21][12])} + {7'd0,(kernel[3][1] ~^ image[21][13])} + {7'd0,(kernel[3][2] ~^ image[21][14])} + {7'd0,(kernel[3][3] ~^ image[21][15])} + {7'd0,(kernel[3][4] ~^ image[21][16])} + {7'd0,(kernel[4][0] ~^ image[22][12])} + {7'd0,(kernel[4][1] ~^ image[22][13])} + {7'd0,(kernel[4][2] ~^ image[22][14])} + {7'd0,(kernel[4][3] ~^ image[22][15])} + {7'd0,(kernel[4][4] ~^ image[22][16])};
assign out_fmap[18][13][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[18][13])} + {7'd0,(kernel[0][1] ~^ image[18][14])} + {7'd0,(kernel[0][2] ~^ image[18][15])} + {7'd0,(kernel[0][3] ~^ image[18][16])} + {7'd0,(kernel[0][4] ~^ image[18][17])} + {7'd0,(kernel[1][0] ~^ image[19][13])} + {7'd0,(kernel[1][1] ~^ image[19][14])} + {7'd0,(kernel[1][2] ~^ image[19][15])} + {7'd0,(kernel[1][3] ~^ image[19][16])} + {7'd0,(kernel[1][4] ~^ image[19][17])} + {7'd0,(kernel[2][0] ~^ image[20][13])} + {7'd0,(kernel[2][1] ~^ image[20][14])} + {7'd0,(kernel[2][2] ~^ image[20][15])} + {7'd0,(kernel[2][3] ~^ image[20][16])} + {7'd0,(kernel[2][4] ~^ image[20][17])} + {7'd0,(kernel[3][0] ~^ image[21][13])} + {7'd0,(kernel[3][1] ~^ image[21][14])} + {7'd0,(kernel[3][2] ~^ image[21][15])} + {7'd0,(kernel[3][3] ~^ image[21][16])} + {7'd0,(kernel[3][4] ~^ image[21][17])} + {7'd0,(kernel[4][0] ~^ image[22][13])} + {7'd0,(kernel[4][1] ~^ image[22][14])} + {7'd0,(kernel[4][2] ~^ image[22][15])} + {7'd0,(kernel[4][3] ~^ image[22][16])} + {7'd0,(kernel[4][4] ~^ image[22][17])};
assign out_fmap[18][14][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[18][14])} + {7'd0,(kernel[0][1] ~^ image[18][15])} + {7'd0,(kernel[0][2] ~^ image[18][16])} + {7'd0,(kernel[0][3] ~^ image[18][17])} + {7'd0,(kernel[0][4] ~^ image[18][18])} + {7'd0,(kernel[1][0] ~^ image[19][14])} + {7'd0,(kernel[1][1] ~^ image[19][15])} + {7'd0,(kernel[1][2] ~^ image[19][16])} + {7'd0,(kernel[1][3] ~^ image[19][17])} + {7'd0,(kernel[1][4] ~^ image[19][18])} + {7'd0,(kernel[2][0] ~^ image[20][14])} + {7'd0,(kernel[2][1] ~^ image[20][15])} + {7'd0,(kernel[2][2] ~^ image[20][16])} + {7'd0,(kernel[2][3] ~^ image[20][17])} + {7'd0,(kernel[2][4] ~^ image[20][18])} + {7'd0,(kernel[3][0] ~^ image[21][14])} + {7'd0,(kernel[3][1] ~^ image[21][15])} + {7'd0,(kernel[3][2] ~^ image[21][16])} + {7'd0,(kernel[3][3] ~^ image[21][17])} + {7'd0,(kernel[3][4] ~^ image[21][18])} + {7'd0,(kernel[4][0] ~^ image[22][14])} + {7'd0,(kernel[4][1] ~^ image[22][15])} + {7'd0,(kernel[4][2] ~^ image[22][16])} + {7'd0,(kernel[4][3] ~^ image[22][17])} + {7'd0,(kernel[4][4] ~^ image[22][18])};
assign out_fmap[18][15][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[18][15])} + {7'd0,(kernel[0][1] ~^ image[18][16])} + {7'd0,(kernel[0][2] ~^ image[18][17])} + {7'd0,(kernel[0][3] ~^ image[18][18])} + {7'd0,(kernel[0][4] ~^ image[18][19])} + {7'd0,(kernel[1][0] ~^ image[19][15])} + {7'd0,(kernel[1][1] ~^ image[19][16])} + {7'd0,(kernel[1][2] ~^ image[19][17])} + {7'd0,(kernel[1][3] ~^ image[19][18])} + {7'd0,(kernel[1][4] ~^ image[19][19])} + {7'd0,(kernel[2][0] ~^ image[20][15])} + {7'd0,(kernel[2][1] ~^ image[20][16])} + {7'd0,(kernel[2][2] ~^ image[20][17])} + {7'd0,(kernel[2][3] ~^ image[20][18])} + {7'd0,(kernel[2][4] ~^ image[20][19])} + {7'd0,(kernel[3][0] ~^ image[21][15])} + {7'd0,(kernel[3][1] ~^ image[21][16])} + {7'd0,(kernel[3][2] ~^ image[21][17])} + {7'd0,(kernel[3][3] ~^ image[21][18])} + {7'd0,(kernel[3][4] ~^ image[21][19])} + {7'd0,(kernel[4][0] ~^ image[22][15])} + {7'd0,(kernel[4][1] ~^ image[22][16])} + {7'd0,(kernel[4][2] ~^ image[22][17])} + {7'd0,(kernel[4][3] ~^ image[22][18])} + {7'd0,(kernel[4][4] ~^ image[22][19])};
assign out_fmap[18][16][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[18][16])} + {7'd0,(kernel[0][1] ~^ image[18][17])} + {7'd0,(kernel[0][2] ~^ image[18][18])} + {7'd0,(kernel[0][3] ~^ image[18][19])} + {7'd0,(kernel[0][4] ~^ image[18][20])} + {7'd0,(kernel[1][0] ~^ image[19][16])} + {7'd0,(kernel[1][1] ~^ image[19][17])} + {7'd0,(kernel[1][2] ~^ image[19][18])} + {7'd0,(kernel[1][3] ~^ image[19][19])} + {7'd0,(kernel[1][4] ~^ image[19][20])} + {7'd0,(kernel[2][0] ~^ image[20][16])} + {7'd0,(kernel[2][1] ~^ image[20][17])} + {7'd0,(kernel[2][2] ~^ image[20][18])} + {7'd0,(kernel[2][3] ~^ image[20][19])} + {7'd0,(kernel[2][4] ~^ image[20][20])} + {7'd0,(kernel[3][0] ~^ image[21][16])} + {7'd0,(kernel[3][1] ~^ image[21][17])} + {7'd0,(kernel[3][2] ~^ image[21][18])} + {7'd0,(kernel[3][3] ~^ image[21][19])} + {7'd0,(kernel[3][4] ~^ image[21][20])} + {7'd0,(kernel[4][0] ~^ image[22][16])} + {7'd0,(kernel[4][1] ~^ image[22][17])} + {7'd0,(kernel[4][2] ~^ image[22][18])} + {7'd0,(kernel[4][3] ~^ image[22][19])} + {7'd0,(kernel[4][4] ~^ image[22][20])};
assign out_fmap[18][17][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[18][17])} + {7'd0,(kernel[0][1] ~^ image[18][18])} + {7'd0,(kernel[0][2] ~^ image[18][19])} + {7'd0,(kernel[0][3] ~^ image[18][20])} + {7'd0,(kernel[0][4] ~^ image[18][21])} + {7'd0,(kernel[1][0] ~^ image[19][17])} + {7'd0,(kernel[1][1] ~^ image[19][18])} + {7'd0,(kernel[1][2] ~^ image[19][19])} + {7'd0,(kernel[1][3] ~^ image[19][20])} + {7'd0,(kernel[1][4] ~^ image[19][21])} + {7'd0,(kernel[2][0] ~^ image[20][17])} + {7'd0,(kernel[2][1] ~^ image[20][18])} + {7'd0,(kernel[2][2] ~^ image[20][19])} + {7'd0,(kernel[2][3] ~^ image[20][20])} + {7'd0,(kernel[2][4] ~^ image[20][21])} + {7'd0,(kernel[3][0] ~^ image[21][17])} + {7'd0,(kernel[3][1] ~^ image[21][18])} + {7'd0,(kernel[3][2] ~^ image[21][19])} + {7'd0,(kernel[3][3] ~^ image[21][20])} + {7'd0,(kernel[3][4] ~^ image[21][21])} + {7'd0,(kernel[4][0] ~^ image[22][17])} + {7'd0,(kernel[4][1] ~^ image[22][18])} + {7'd0,(kernel[4][2] ~^ image[22][19])} + {7'd0,(kernel[4][3] ~^ image[22][20])} + {7'd0,(kernel[4][4] ~^ image[22][21])};
assign out_fmap[18][18][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[18][18])} + {7'd0,(kernel[0][1] ~^ image[18][19])} + {7'd0,(kernel[0][2] ~^ image[18][20])} + {7'd0,(kernel[0][3] ~^ image[18][21])} + {7'd0,(kernel[0][4] ~^ image[18][22])} + {7'd0,(kernel[1][0] ~^ image[19][18])} + {7'd0,(kernel[1][1] ~^ image[19][19])} + {7'd0,(kernel[1][2] ~^ image[19][20])} + {7'd0,(kernel[1][3] ~^ image[19][21])} + {7'd0,(kernel[1][4] ~^ image[19][22])} + {7'd0,(kernel[2][0] ~^ image[20][18])} + {7'd0,(kernel[2][1] ~^ image[20][19])} + {7'd0,(kernel[2][2] ~^ image[20][20])} + {7'd0,(kernel[2][3] ~^ image[20][21])} + {7'd0,(kernel[2][4] ~^ image[20][22])} + {7'd0,(kernel[3][0] ~^ image[21][18])} + {7'd0,(kernel[3][1] ~^ image[21][19])} + {7'd0,(kernel[3][2] ~^ image[21][20])} + {7'd0,(kernel[3][3] ~^ image[21][21])} + {7'd0,(kernel[3][4] ~^ image[21][22])} + {7'd0,(kernel[4][0] ~^ image[22][18])} + {7'd0,(kernel[4][1] ~^ image[22][19])} + {7'd0,(kernel[4][2] ~^ image[22][20])} + {7'd0,(kernel[4][3] ~^ image[22][21])} + {7'd0,(kernel[4][4] ~^ image[22][22])};
assign out_fmap[18][19][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[18][19])} + {7'd0,(kernel[0][1] ~^ image[18][20])} + {7'd0,(kernel[0][2] ~^ image[18][21])} + {7'd0,(kernel[0][3] ~^ image[18][22])} + {7'd0,(kernel[0][4] ~^ image[18][23])} + {7'd0,(kernel[1][0] ~^ image[19][19])} + {7'd0,(kernel[1][1] ~^ image[19][20])} + {7'd0,(kernel[1][2] ~^ image[19][21])} + {7'd0,(kernel[1][3] ~^ image[19][22])} + {7'd0,(kernel[1][4] ~^ image[19][23])} + {7'd0,(kernel[2][0] ~^ image[20][19])} + {7'd0,(kernel[2][1] ~^ image[20][20])} + {7'd0,(kernel[2][2] ~^ image[20][21])} + {7'd0,(kernel[2][3] ~^ image[20][22])} + {7'd0,(kernel[2][4] ~^ image[20][23])} + {7'd0,(kernel[3][0] ~^ image[21][19])} + {7'd0,(kernel[3][1] ~^ image[21][20])} + {7'd0,(kernel[3][2] ~^ image[21][21])} + {7'd0,(kernel[3][3] ~^ image[21][22])} + {7'd0,(kernel[3][4] ~^ image[21][23])} + {7'd0,(kernel[4][0] ~^ image[22][19])} + {7'd0,(kernel[4][1] ~^ image[22][20])} + {7'd0,(kernel[4][2] ~^ image[22][21])} + {7'd0,(kernel[4][3] ~^ image[22][22])} + {7'd0,(kernel[4][4] ~^ image[22][23])};
assign out_fmap[18][20][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[18][20])} + {7'd0,(kernel[0][1] ~^ image[18][21])} + {7'd0,(kernel[0][2] ~^ image[18][22])} + {7'd0,(kernel[0][3] ~^ image[18][23])} + {7'd0,(kernel[0][4] ~^ image[18][24])} + {7'd0,(kernel[1][0] ~^ image[19][20])} + {7'd0,(kernel[1][1] ~^ image[19][21])} + {7'd0,(kernel[1][2] ~^ image[19][22])} + {7'd0,(kernel[1][3] ~^ image[19][23])} + {7'd0,(kernel[1][4] ~^ image[19][24])} + {7'd0,(kernel[2][0] ~^ image[20][20])} + {7'd0,(kernel[2][1] ~^ image[20][21])} + {7'd0,(kernel[2][2] ~^ image[20][22])} + {7'd0,(kernel[2][3] ~^ image[20][23])} + {7'd0,(kernel[2][4] ~^ image[20][24])} + {7'd0,(kernel[3][0] ~^ image[21][20])} + {7'd0,(kernel[3][1] ~^ image[21][21])} + {7'd0,(kernel[3][2] ~^ image[21][22])} + {7'd0,(kernel[3][3] ~^ image[21][23])} + {7'd0,(kernel[3][4] ~^ image[21][24])} + {7'd0,(kernel[4][0] ~^ image[22][20])} + {7'd0,(kernel[4][1] ~^ image[22][21])} + {7'd0,(kernel[4][2] ~^ image[22][22])} + {7'd0,(kernel[4][3] ~^ image[22][23])} + {7'd0,(kernel[4][4] ~^ image[22][24])};
assign out_fmap[18][21][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[18][21])} + {7'd0,(kernel[0][1] ~^ image[18][22])} + {7'd0,(kernel[0][2] ~^ image[18][23])} + {7'd0,(kernel[0][3] ~^ image[18][24])} + {7'd0,(kernel[0][4] ~^ image[18][25])} + {7'd0,(kernel[1][0] ~^ image[19][21])} + {7'd0,(kernel[1][1] ~^ image[19][22])} + {7'd0,(kernel[1][2] ~^ image[19][23])} + {7'd0,(kernel[1][3] ~^ image[19][24])} + {7'd0,(kernel[1][4] ~^ image[19][25])} + {7'd0,(kernel[2][0] ~^ image[20][21])} + {7'd0,(kernel[2][1] ~^ image[20][22])} + {7'd0,(kernel[2][2] ~^ image[20][23])} + {7'd0,(kernel[2][3] ~^ image[20][24])} + {7'd0,(kernel[2][4] ~^ image[20][25])} + {7'd0,(kernel[3][0] ~^ image[21][21])} + {7'd0,(kernel[3][1] ~^ image[21][22])} + {7'd0,(kernel[3][2] ~^ image[21][23])} + {7'd0,(kernel[3][3] ~^ image[21][24])} + {7'd0,(kernel[3][4] ~^ image[21][25])} + {7'd0,(kernel[4][0] ~^ image[22][21])} + {7'd0,(kernel[4][1] ~^ image[22][22])} + {7'd0,(kernel[4][2] ~^ image[22][23])} + {7'd0,(kernel[4][3] ~^ image[22][24])} + {7'd0,(kernel[4][4] ~^ image[22][25])};
assign out_fmap[18][22][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[18][22])} + {7'd0,(kernel[0][1] ~^ image[18][23])} + {7'd0,(kernel[0][2] ~^ image[18][24])} + {7'd0,(kernel[0][3] ~^ image[18][25])} + {7'd0,(kernel[0][4] ~^ image[18][26])} + {7'd0,(kernel[1][0] ~^ image[19][22])} + {7'd0,(kernel[1][1] ~^ image[19][23])} + {7'd0,(kernel[1][2] ~^ image[19][24])} + {7'd0,(kernel[1][3] ~^ image[19][25])} + {7'd0,(kernel[1][4] ~^ image[19][26])} + {7'd0,(kernel[2][0] ~^ image[20][22])} + {7'd0,(kernel[2][1] ~^ image[20][23])} + {7'd0,(kernel[2][2] ~^ image[20][24])} + {7'd0,(kernel[2][3] ~^ image[20][25])} + {7'd0,(kernel[2][4] ~^ image[20][26])} + {7'd0,(kernel[3][0] ~^ image[21][22])} + {7'd0,(kernel[3][1] ~^ image[21][23])} + {7'd0,(kernel[3][2] ~^ image[21][24])} + {7'd0,(kernel[3][3] ~^ image[21][25])} + {7'd0,(kernel[3][4] ~^ image[21][26])} + {7'd0,(kernel[4][0] ~^ image[22][22])} + {7'd0,(kernel[4][1] ~^ image[22][23])} + {7'd0,(kernel[4][2] ~^ image[22][24])} + {7'd0,(kernel[4][3] ~^ image[22][25])} + {7'd0,(kernel[4][4] ~^ image[22][26])};
assign out_fmap[18][23][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[18][23])} + {7'd0,(kernel[0][1] ~^ image[18][24])} + {7'd0,(kernel[0][2] ~^ image[18][25])} + {7'd0,(kernel[0][3] ~^ image[18][26])} + {7'd0,(kernel[0][4] ~^ image[18][27])} + {7'd0,(kernel[1][0] ~^ image[19][23])} + {7'd0,(kernel[1][1] ~^ image[19][24])} + {7'd0,(kernel[1][2] ~^ image[19][25])} + {7'd0,(kernel[1][3] ~^ image[19][26])} + {7'd0,(kernel[1][4] ~^ image[19][27])} + {7'd0,(kernel[2][0] ~^ image[20][23])} + {7'd0,(kernel[2][1] ~^ image[20][24])} + {7'd0,(kernel[2][2] ~^ image[20][25])} + {7'd0,(kernel[2][3] ~^ image[20][26])} + {7'd0,(kernel[2][4] ~^ image[20][27])} + {7'd0,(kernel[3][0] ~^ image[21][23])} + {7'd0,(kernel[3][1] ~^ image[21][24])} + {7'd0,(kernel[3][2] ~^ image[21][25])} + {7'd0,(kernel[3][3] ~^ image[21][26])} + {7'd0,(kernel[3][4] ~^ image[21][27])} + {7'd0,(kernel[4][0] ~^ image[22][23])} + {7'd0,(kernel[4][1] ~^ image[22][24])} + {7'd0,(kernel[4][2] ~^ image[22][25])} + {7'd0,(kernel[4][3] ~^ image[22][26])} + {7'd0,(kernel[4][4] ~^ image[22][27])};
assign out_fmap[19][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[19][0])} + {7'd0,(kernel[0][1] ~^ image[19][1])} + {7'd0,(kernel[0][2] ~^ image[19][2])} + {7'd0,(kernel[0][3] ~^ image[19][3])} + {7'd0,(kernel[0][4] ~^ image[19][4])} + {7'd0,(kernel[1][0] ~^ image[20][0])} + {7'd0,(kernel[1][1] ~^ image[20][1])} + {7'd0,(kernel[1][2] ~^ image[20][2])} + {7'd0,(kernel[1][3] ~^ image[20][3])} + {7'd0,(kernel[1][4] ~^ image[20][4])} + {7'd0,(kernel[2][0] ~^ image[21][0])} + {7'd0,(kernel[2][1] ~^ image[21][1])} + {7'd0,(kernel[2][2] ~^ image[21][2])} + {7'd0,(kernel[2][3] ~^ image[21][3])} + {7'd0,(kernel[2][4] ~^ image[21][4])} + {7'd0,(kernel[3][0] ~^ image[22][0])} + {7'd0,(kernel[3][1] ~^ image[22][1])} + {7'd0,(kernel[3][2] ~^ image[22][2])} + {7'd0,(kernel[3][3] ~^ image[22][3])} + {7'd0,(kernel[3][4] ~^ image[22][4])} + {7'd0,(kernel[4][0] ~^ image[23][0])} + {7'd0,(kernel[4][1] ~^ image[23][1])} + {7'd0,(kernel[4][2] ~^ image[23][2])} + {7'd0,(kernel[4][3] ~^ image[23][3])} + {7'd0,(kernel[4][4] ~^ image[23][4])};
assign out_fmap[19][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[19][1])} + {7'd0,(kernel[0][1] ~^ image[19][2])} + {7'd0,(kernel[0][2] ~^ image[19][3])} + {7'd0,(kernel[0][3] ~^ image[19][4])} + {7'd0,(kernel[0][4] ~^ image[19][5])} + {7'd0,(kernel[1][0] ~^ image[20][1])} + {7'd0,(kernel[1][1] ~^ image[20][2])} + {7'd0,(kernel[1][2] ~^ image[20][3])} + {7'd0,(kernel[1][3] ~^ image[20][4])} + {7'd0,(kernel[1][4] ~^ image[20][5])} + {7'd0,(kernel[2][0] ~^ image[21][1])} + {7'd0,(kernel[2][1] ~^ image[21][2])} + {7'd0,(kernel[2][2] ~^ image[21][3])} + {7'd0,(kernel[2][3] ~^ image[21][4])} + {7'd0,(kernel[2][4] ~^ image[21][5])} + {7'd0,(kernel[3][0] ~^ image[22][1])} + {7'd0,(kernel[3][1] ~^ image[22][2])} + {7'd0,(kernel[3][2] ~^ image[22][3])} + {7'd0,(kernel[3][3] ~^ image[22][4])} + {7'd0,(kernel[3][4] ~^ image[22][5])} + {7'd0,(kernel[4][0] ~^ image[23][1])} + {7'd0,(kernel[4][1] ~^ image[23][2])} + {7'd0,(kernel[4][2] ~^ image[23][3])} + {7'd0,(kernel[4][3] ~^ image[23][4])} + {7'd0,(kernel[4][4] ~^ image[23][5])};
assign out_fmap[19][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[19][2])} + {7'd0,(kernel[0][1] ~^ image[19][3])} + {7'd0,(kernel[0][2] ~^ image[19][4])} + {7'd0,(kernel[0][3] ~^ image[19][5])} + {7'd0,(kernel[0][4] ~^ image[19][6])} + {7'd0,(kernel[1][0] ~^ image[20][2])} + {7'd0,(kernel[1][1] ~^ image[20][3])} + {7'd0,(kernel[1][2] ~^ image[20][4])} + {7'd0,(kernel[1][3] ~^ image[20][5])} + {7'd0,(kernel[1][4] ~^ image[20][6])} + {7'd0,(kernel[2][0] ~^ image[21][2])} + {7'd0,(kernel[2][1] ~^ image[21][3])} + {7'd0,(kernel[2][2] ~^ image[21][4])} + {7'd0,(kernel[2][3] ~^ image[21][5])} + {7'd0,(kernel[2][4] ~^ image[21][6])} + {7'd0,(kernel[3][0] ~^ image[22][2])} + {7'd0,(kernel[3][1] ~^ image[22][3])} + {7'd0,(kernel[3][2] ~^ image[22][4])} + {7'd0,(kernel[3][3] ~^ image[22][5])} + {7'd0,(kernel[3][4] ~^ image[22][6])} + {7'd0,(kernel[4][0] ~^ image[23][2])} + {7'd0,(kernel[4][1] ~^ image[23][3])} + {7'd0,(kernel[4][2] ~^ image[23][4])} + {7'd0,(kernel[4][3] ~^ image[23][5])} + {7'd0,(kernel[4][4] ~^ image[23][6])};
assign out_fmap[19][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[19][3])} + {7'd0,(kernel[0][1] ~^ image[19][4])} + {7'd0,(kernel[0][2] ~^ image[19][5])} + {7'd0,(kernel[0][3] ~^ image[19][6])} + {7'd0,(kernel[0][4] ~^ image[19][7])} + {7'd0,(kernel[1][0] ~^ image[20][3])} + {7'd0,(kernel[1][1] ~^ image[20][4])} + {7'd0,(kernel[1][2] ~^ image[20][5])} + {7'd0,(kernel[1][3] ~^ image[20][6])} + {7'd0,(kernel[1][4] ~^ image[20][7])} + {7'd0,(kernel[2][0] ~^ image[21][3])} + {7'd0,(kernel[2][1] ~^ image[21][4])} + {7'd0,(kernel[2][2] ~^ image[21][5])} + {7'd0,(kernel[2][3] ~^ image[21][6])} + {7'd0,(kernel[2][4] ~^ image[21][7])} + {7'd0,(kernel[3][0] ~^ image[22][3])} + {7'd0,(kernel[3][1] ~^ image[22][4])} + {7'd0,(kernel[3][2] ~^ image[22][5])} + {7'd0,(kernel[3][3] ~^ image[22][6])} + {7'd0,(kernel[3][4] ~^ image[22][7])} + {7'd0,(kernel[4][0] ~^ image[23][3])} + {7'd0,(kernel[4][1] ~^ image[23][4])} + {7'd0,(kernel[4][2] ~^ image[23][5])} + {7'd0,(kernel[4][3] ~^ image[23][6])} + {7'd0,(kernel[4][4] ~^ image[23][7])};
assign out_fmap[19][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[19][4])} + {7'd0,(kernel[0][1] ~^ image[19][5])} + {7'd0,(kernel[0][2] ~^ image[19][6])} + {7'd0,(kernel[0][3] ~^ image[19][7])} + {7'd0,(kernel[0][4] ~^ image[19][8])} + {7'd0,(kernel[1][0] ~^ image[20][4])} + {7'd0,(kernel[1][1] ~^ image[20][5])} + {7'd0,(kernel[1][2] ~^ image[20][6])} + {7'd0,(kernel[1][3] ~^ image[20][7])} + {7'd0,(kernel[1][4] ~^ image[20][8])} + {7'd0,(kernel[2][0] ~^ image[21][4])} + {7'd0,(kernel[2][1] ~^ image[21][5])} + {7'd0,(kernel[2][2] ~^ image[21][6])} + {7'd0,(kernel[2][3] ~^ image[21][7])} + {7'd0,(kernel[2][4] ~^ image[21][8])} + {7'd0,(kernel[3][0] ~^ image[22][4])} + {7'd0,(kernel[3][1] ~^ image[22][5])} + {7'd0,(kernel[3][2] ~^ image[22][6])} + {7'd0,(kernel[3][3] ~^ image[22][7])} + {7'd0,(kernel[3][4] ~^ image[22][8])} + {7'd0,(kernel[4][0] ~^ image[23][4])} + {7'd0,(kernel[4][1] ~^ image[23][5])} + {7'd0,(kernel[4][2] ~^ image[23][6])} + {7'd0,(kernel[4][3] ~^ image[23][7])} + {7'd0,(kernel[4][4] ~^ image[23][8])};
assign out_fmap[19][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[19][5])} + {7'd0,(kernel[0][1] ~^ image[19][6])} + {7'd0,(kernel[0][2] ~^ image[19][7])} + {7'd0,(kernel[0][3] ~^ image[19][8])} + {7'd0,(kernel[0][4] ~^ image[19][9])} + {7'd0,(kernel[1][0] ~^ image[20][5])} + {7'd0,(kernel[1][1] ~^ image[20][6])} + {7'd0,(kernel[1][2] ~^ image[20][7])} + {7'd0,(kernel[1][3] ~^ image[20][8])} + {7'd0,(kernel[1][4] ~^ image[20][9])} + {7'd0,(kernel[2][0] ~^ image[21][5])} + {7'd0,(kernel[2][1] ~^ image[21][6])} + {7'd0,(kernel[2][2] ~^ image[21][7])} + {7'd0,(kernel[2][3] ~^ image[21][8])} + {7'd0,(kernel[2][4] ~^ image[21][9])} + {7'd0,(kernel[3][0] ~^ image[22][5])} + {7'd0,(kernel[3][1] ~^ image[22][6])} + {7'd0,(kernel[3][2] ~^ image[22][7])} + {7'd0,(kernel[3][3] ~^ image[22][8])} + {7'd0,(kernel[3][4] ~^ image[22][9])} + {7'd0,(kernel[4][0] ~^ image[23][5])} + {7'd0,(kernel[4][1] ~^ image[23][6])} + {7'd0,(kernel[4][2] ~^ image[23][7])} + {7'd0,(kernel[4][3] ~^ image[23][8])} + {7'd0,(kernel[4][4] ~^ image[23][9])};
assign out_fmap[19][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[19][6])} + {7'd0,(kernel[0][1] ~^ image[19][7])} + {7'd0,(kernel[0][2] ~^ image[19][8])} + {7'd0,(kernel[0][3] ~^ image[19][9])} + {7'd0,(kernel[0][4] ~^ image[19][10])} + {7'd0,(kernel[1][0] ~^ image[20][6])} + {7'd0,(kernel[1][1] ~^ image[20][7])} + {7'd0,(kernel[1][2] ~^ image[20][8])} + {7'd0,(kernel[1][3] ~^ image[20][9])} + {7'd0,(kernel[1][4] ~^ image[20][10])} + {7'd0,(kernel[2][0] ~^ image[21][6])} + {7'd0,(kernel[2][1] ~^ image[21][7])} + {7'd0,(kernel[2][2] ~^ image[21][8])} + {7'd0,(kernel[2][3] ~^ image[21][9])} + {7'd0,(kernel[2][4] ~^ image[21][10])} + {7'd0,(kernel[3][0] ~^ image[22][6])} + {7'd0,(kernel[3][1] ~^ image[22][7])} + {7'd0,(kernel[3][2] ~^ image[22][8])} + {7'd0,(kernel[3][3] ~^ image[22][9])} + {7'd0,(kernel[3][4] ~^ image[22][10])} + {7'd0,(kernel[4][0] ~^ image[23][6])} + {7'd0,(kernel[4][1] ~^ image[23][7])} + {7'd0,(kernel[4][2] ~^ image[23][8])} + {7'd0,(kernel[4][3] ~^ image[23][9])} + {7'd0,(kernel[4][4] ~^ image[23][10])};
assign out_fmap[19][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[19][7])} + {7'd0,(kernel[0][1] ~^ image[19][8])} + {7'd0,(kernel[0][2] ~^ image[19][9])} + {7'd0,(kernel[0][3] ~^ image[19][10])} + {7'd0,(kernel[0][4] ~^ image[19][11])} + {7'd0,(kernel[1][0] ~^ image[20][7])} + {7'd0,(kernel[1][1] ~^ image[20][8])} + {7'd0,(kernel[1][2] ~^ image[20][9])} + {7'd0,(kernel[1][3] ~^ image[20][10])} + {7'd0,(kernel[1][4] ~^ image[20][11])} + {7'd0,(kernel[2][0] ~^ image[21][7])} + {7'd0,(kernel[2][1] ~^ image[21][8])} + {7'd0,(kernel[2][2] ~^ image[21][9])} + {7'd0,(kernel[2][3] ~^ image[21][10])} + {7'd0,(kernel[2][4] ~^ image[21][11])} + {7'd0,(kernel[3][0] ~^ image[22][7])} + {7'd0,(kernel[3][1] ~^ image[22][8])} + {7'd0,(kernel[3][2] ~^ image[22][9])} + {7'd0,(kernel[3][3] ~^ image[22][10])} + {7'd0,(kernel[3][4] ~^ image[22][11])} + {7'd0,(kernel[4][0] ~^ image[23][7])} + {7'd0,(kernel[4][1] ~^ image[23][8])} + {7'd0,(kernel[4][2] ~^ image[23][9])} + {7'd0,(kernel[4][3] ~^ image[23][10])} + {7'd0,(kernel[4][4] ~^ image[23][11])};
assign out_fmap[19][8][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[19][8])} + {7'd0,(kernel[0][1] ~^ image[19][9])} + {7'd0,(kernel[0][2] ~^ image[19][10])} + {7'd0,(kernel[0][3] ~^ image[19][11])} + {7'd0,(kernel[0][4] ~^ image[19][12])} + {7'd0,(kernel[1][0] ~^ image[20][8])} + {7'd0,(kernel[1][1] ~^ image[20][9])} + {7'd0,(kernel[1][2] ~^ image[20][10])} + {7'd0,(kernel[1][3] ~^ image[20][11])} + {7'd0,(kernel[1][4] ~^ image[20][12])} + {7'd0,(kernel[2][0] ~^ image[21][8])} + {7'd0,(kernel[2][1] ~^ image[21][9])} + {7'd0,(kernel[2][2] ~^ image[21][10])} + {7'd0,(kernel[2][3] ~^ image[21][11])} + {7'd0,(kernel[2][4] ~^ image[21][12])} + {7'd0,(kernel[3][0] ~^ image[22][8])} + {7'd0,(kernel[3][1] ~^ image[22][9])} + {7'd0,(kernel[3][2] ~^ image[22][10])} + {7'd0,(kernel[3][3] ~^ image[22][11])} + {7'd0,(kernel[3][4] ~^ image[22][12])} + {7'd0,(kernel[4][0] ~^ image[23][8])} + {7'd0,(kernel[4][1] ~^ image[23][9])} + {7'd0,(kernel[4][2] ~^ image[23][10])} + {7'd0,(kernel[4][3] ~^ image[23][11])} + {7'd0,(kernel[4][4] ~^ image[23][12])};
assign out_fmap[19][9][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[19][9])} + {7'd0,(kernel[0][1] ~^ image[19][10])} + {7'd0,(kernel[0][2] ~^ image[19][11])} + {7'd0,(kernel[0][3] ~^ image[19][12])} + {7'd0,(kernel[0][4] ~^ image[19][13])} + {7'd0,(kernel[1][0] ~^ image[20][9])} + {7'd0,(kernel[1][1] ~^ image[20][10])} + {7'd0,(kernel[1][2] ~^ image[20][11])} + {7'd0,(kernel[1][3] ~^ image[20][12])} + {7'd0,(kernel[1][4] ~^ image[20][13])} + {7'd0,(kernel[2][0] ~^ image[21][9])} + {7'd0,(kernel[2][1] ~^ image[21][10])} + {7'd0,(kernel[2][2] ~^ image[21][11])} + {7'd0,(kernel[2][3] ~^ image[21][12])} + {7'd0,(kernel[2][4] ~^ image[21][13])} + {7'd0,(kernel[3][0] ~^ image[22][9])} + {7'd0,(kernel[3][1] ~^ image[22][10])} + {7'd0,(kernel[3][2] ~^ image[22][11])} + {7'd0,(kernel[3][3] ~^ image[22][12])} + {7'd0,(kernel[3][4] ~^ image[22][13])} + {7'd0,(kernel[4][0] ~^ image[23][9])} + {7'd0,(kernel[4][1] ~^ image[23][10])} + {7'd0,(kernel[4][2] ~^ image[23][11])} + {7'd0,(kernel[4][3] ~^ image[23][12])} + {7'd0,(kernel[4][4] ~^ image[23][13])};
assign out_fmap[19][10][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[19][10])} + {7'd0,(kernel[0][1] ~^ image[19][11])} + {7'd0,(kernel[0][2] ~^ image[19][12])} + {7'd0,(kernel[0][3] ~^ image[19][13])} + {7'd0,(kernel[0][4] ~^ image[19][14])} + {7'd0,(kernel[1][0] ~^ image[20][10])} + {7'd0,(kernel[1][1] ~^ image[20][11])} + {7'd0,(kernel[1][2] ~^ image[20][12])} + {7'd0,(kernel[1][3] ~^ image[20][13])} + {7'd0,(kernel[1][4] ~^ image[20][14])} + {7'd0,(kernel[2][0] ~^ image[21][10])} + {7'd0,(kernel[2][1] ~^ image[21][11])} + {7'd0,(kernel[2][2] ~^ image[21][12])} + {7'd0,(kernel[2][3] ~^ image[21][13])} + {7'd0,(kernel[2][4] ~^ image[21][14])} + {7'd0,(kernel[3][0] ~^ image[22][10])} + {7'd0,(kernel[3][1] ~^ image[22][11])} + {7'd0,(kernel[3][2] ~^ image[22][12])} + {7'd0,(kernel[3][3] ~^ image[22][13])} + {7'd0,(kernel[3][4] ~^ image[22][14])} + {7'd0,(kernel[4][0] ~^ image[23][10])} + {7'd0,(kernel[4][1] ~^ image[23][11])} + {7'd0,(kernel[4][2] ~^ image[23][12])} + {7'd0,(kernel[4][3] ~^ image[23][13])} + {7'd0,(kernel[4][4] ~^ image[23][14])};
assign out_fmap[19][11][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[19][11])} + {7'd0,(kernel[0][1] ~^ image[19][12])} + {7'd0,(kernel[0][2] ~^ image[19][13])} + {7'd0,(kernel[0][3] ~^ image[19][14])} + {7'd0,(kernel[0][4] ~^ image[19][15])} + {7'd0,(kernel[1][0] ~^ image[20][11])} + {7'd0,(kernel[1][1] ~^ image[20][12])} + {7'd0,(kernel[1][2] ~^ image[20][13])} + {7'd0,(kernel[1][3] ~^ image[20][14])} + {7'd0,(kernel[1][4] ~^ image[20][15])} + {7'd0,(kernel[2][0] ~^ image[21][11])} + {7'd0,(kernel[2][1] ~^ image[21][12])} + {7'd0,(kernel[2][2] ~^ image[21][13])} + {7'd0,(kernel[2][3] ~^ image[21][14])} + {7'd0,(kernel[2][4] ~^ image[21][15])} + {7'd0,(kernel[3][0] ~^ image[22][11])} + {7'd0,(kernel[3][1] ~^ image[22][12])} + {7'd0,(kernel[3][2] ~^ image[22][13])} + {7'd0,(kernel[3][3] ~^ image[22][14])} + {7'd0,(kernel[3][4] ~^ image[22][15])} + {7'd0,(kernel[4][0] ~^ image[23][11])} + {7'd0,(kernel[4][1] ~^ image[23][12])} + {7'd0,(kernel[4][2] ~^ image[23][13])} + {7'd0,(kernel[4][3] ~^ image[23][14])} + {7'd0,(kernel[4][4] ~^ image[23][15])};
assign out_fmap[19][12][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[19][12])} + {7'd0,(kernel[0][1] ~^ image[19][13])} + {7'd0,(kernel[0][2] ~^ image[19][14])} + {7'd0,(kernel[0][3] ~^ image[19][15])} + {7'd0,(kernel[0][4] ~^ image[19][16])} + {7'd0,(kernel[1][0] ~^ image[20][12])} + {7'd0,(kernel[1][1] ~^ image[20][13])} + {7'd0,(kernel[1][2] ~^ image[20][14])} + {7'd0,(kernel[1][3] ~^ image[20][15])} + {7'd0,(kernel[1][4] ~^ image[20][16])} + {7'd0,(kernel[2][0] ~^ image[21][12])} + {7'd0,(kernel[2][1] ~^ image[21][13])} + {7'd0,(kernel[2][2] ~^ image[21][14])} + {7'd0,(kernel[2][3] ~^ image[21][15])} + {7'd0,(kernel[2][4] ~^ image[21][16])} + {7'd0,(kernel[3][0] ~^ image[22][12])} + {7'd0,(kernel[3][1] ~^ image[22][13])} + {7'd0,(kernel[3][2] ~^ image[22][14])} + {7'd0,(kernel[3][3] ~^ image[22][15])} + {7'd0,(kernel[3][4] ~^ image[22][16])} + {7'd0,(kernel[4][0] ~^ image[23][12])} + {7'd0,(kernel[4][1] ~^ image[23][13])} + {7'd0,(kernel[4][2] ~^ image[23][14])} + {7'd0,(kernel[4][3] ~^ image[23][15])} + {7'd0,(kernel[4][4] ~^ image[23][16])};
assign out_fmap[19][13][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[19][13])} + {7'd0,(kernel[0][1] ~^ image[19][14])} + {7'd0,(kernel[0][2] ~^ image[19][15])} + {7'd0,(kernel[0][3] ~^ image[19][16])} + {7'd0,(kernel[0][4] ~^ image[19][17])} + {7'd0,(kernel[1][0] ~^ image[20][13])} + {7'd0,(kernel[1][1] ~^ image[20][14])} + {7'd0,(kernel[1][2] ~^ image[20][15])} + {7'd0,(kernel[1][3] ~^ image[20][16])} + {7'd0,(kernel[1][4] ~^ image[20][17])} + {7'd0,(kernel[2][0] ~^ image[21][13])} + {7'd0,(kernel[2][1] ~^ image[21][14])} + {7'd0,(kernel[2][2] ~^ image[21][15])} + {7'd0,(kernel[2][3] ~^ image[21][16])} + {7'd0,(kernel[2][4] ~^ image[21][17])} + {7'd0,(kernel[3][0] ~^ image[22][13])} + {7'd0,(kernel[3][1] ~^ image[22][14])} + {7'd0,(kernel[3][2] ~^ image[22][15])} + {7'd0,(kernel[3][3] ~^ image[22][16])} + {7'd0,(kernel[3][4] ~^ image[22][17])} + {7'd0,(kernel[4][0] ~^ image[23][13])} + {7'd0,(kernel[4][1] ~^ image[23][14])} + {7'd0,(kernel[4][2] ~^ image[23][15])} + {7'd0,(kernel[4][3] ~^ image[23][16])} + {7'd0,(kernel[4][4] ~^ image[23][17])};
assign out_fmap[19][14][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[19][14])} + {7'd0,(kernel[0][1] ~^ image[19][15])} + {7'd0,(kernel[0][2] ~^ image[19][16])} + {7'd0,(kernel[0][3] ~^ image[19][17])} + {7'd0,(kernel[0][4] ~^ image[19][18])} + {7'd0,(kernel[1][0] ~^ image[20][14])} + {7'd0,(kernel[1][1] ~^ image[20][15])} + {7'd0,(kernel[1][2] ~^ image[20][16])} + {7'd0,(kernel[1][3] ~^ image[20][17])} + {7'd0,(kernel[1][4] ~^ image[20][18])} + {7'd0,(kernel[2][0] ~^ image[21][14])} + {7'd0,(kernel[2][1] ~^ image[21][15])} + {7'd0,(kernel[2][2] ~^ image[21][16])} + {7'd0,(kernel[2][3] ~^ image[21][17])} + {7'd0,(kernel[2][4] ~^ image[21][18])} + {7'd0,(kernel[3][0] ~^ image[22][14])} + {7'd0,(kernel[3][1] ~^ image[22][15])} + {7'd0,(kernel[3][2] ~^ image[22][16])} + {7'd0,(kernel[3][3] ~^ image[22][17])} + {7'd0,(kernel[3][4] ~^ image[22][18])} + {7'd0,(kernel[4][0] ~^ image[23][14])} + {7'd0,(kernel[4][1] ~^ image[23][15])} + {7'd0,(kernel[4][2] ~^ image[23][16])} + {7'd0,(kernel[4][3] ~^ image[23][17])} + {7'd0,(kernel[4][4] ~^ image[23][18])};
assign out_fmap[19][15][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[19][15])} + {7'd0,(kernel[0][1] ~^ image[19][16])} + {7'd0,(kernel[0][2] ~^ image[19][17])} + {7'd0,(kernel[0][3] ~^ image[19][18])} + {7'd0,(kernel[0][4] ~^ image[19][19])} + {7'd0,(kernel[1][0] ~^ image[20][15])} + {7'd0,(kernel[1][1] ~^ image[20][16])} + {7'd0,(kernel[1][2] ~^ image[20][17])} + {7'd0,(kernel[1][3] ~^ image[20][18])} + {7'd0,(kernel[1][4] ~^ image[20][19])} + {7'd0,(kernel[2][0] ~^ image[21][15])} + {7'd0,(kernel[2][1] ~^ image[21][16])} + {7'd0,(kernel[2][2] ~^ image[21][17])} + {7'd0,(kernel[2][3] ~^ image[21][18])} + {7'd0,(kernel[2][4] ~^ image[21][19])} + {7'd0,(kernel[3][0] ~^ image[22][15])} + {7'd0,(kernel[3][1] ~^ image[22][16])} + {7'd0,(kernel[3][2] ~^ image[22][17])} + {7'd0,(kernel[3][3] ~^ image[22][18])} + {7'd0,(kernel[3][4] ~^ image[22][19])} + {7'd0,(kernel[4][0] ~^ image[23][15])} + {7'd0,(kernel[4][1] ~^ image[23][16])} + {7'd0,(kernel[4][2] ~^ image[23][17])} + {7'd0,(kernel[4][3] ~^ image[23][18])} + {7'd0,(kernel[4][4] ~^ image[23][19])};
assign out_fmap[19][16][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[19][16])} + {7'd0,(kernel[0][1] ~^ image[19][17])} + {7'd0,(kernel[0][2] ~^ image[19][18])} + {7'd0,(kernel[0][3] ~^ image[19][19])} + {7'd0,(kernel[0][4] ~^ image[19][20])} + {7'd0,(kernel[1][0] ~^ image[20][16])} + {7'd0,(kernel[1][1] ~^ image[20][17])} + {7'd0,(kernel[1][2] ~^ image[20][18])} + {7'd0,(kernel[1][3] ~^ image[20][19])} + {7'd0,(kernel[1][4] ~^ image[20][20])} + {7'd0,(kernel[2][0] ~^ image[21][16])} + {7'd0,(kernel[2][1] ~^ image[21][17])} + {7'd0,(kernel[2][2] ~^ image[21][18])} + {7'd0,(kernel[2][3] ~^ image[21][19])} + {7'd0,(kernel[2][4] ~^ image[21][20])} + {7'd0,(kernel[3][0] ~^ image[22][16])} + {7'd0,(kernel[3][1] ~^ image[22][17])} + {7'd0,(kernel[3][2] ~^ image[22][18])} + {7'd0,(kernel[3][3] ~^ image[22][19])} + {7'd0,(kernel[3][4] ~^ image[22][20])} + {7'd0,(kernel[4][0] ~^ image[23][16])} + {7'd0,(kernel[4][1] ~^ image[23][17])} + {7'd0,(kernel[4][2] ~^ image[23][18])} + {7'd0,(kernel[4][3] ~^ image[23][19])} + {7'd0,(kernel[4][4] ~^ image[23][20])};
assign out_fmap[19][17][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[19][17])} + {7'd0,(kernel[0][1] ~^ image[19][18])} + {7'd0,(kernel[0][2] ~^ image[19][19])} + {7'd0,(kernel[0][3] ~^ image[19][20])} + {7'd0,(kernel[0][4] ~^ image[19][21])} + {7'd0,(kernel[1][0] ~^ image[20][17])} + {7'd0,(kernel[1][1] ~^ image[20][18])} + {7'd0,(kernel[1][2] ~^ image[20][19])} + {7'd0,(kernel[1][3] ~^ image[20][20])} + {7'd0,(kernel[1][4] ~^ image[20][21])} + {7'd0,(kernel[2][0] ~^ image[21][17])} + {7'd0,(kernel[2][1] ~^ image[21][18])} + {7'd0,(kernel[2][2] ~^ image[21][19])} + {7'd0,(kernel[2][3] ~^ image[21][20])} + {7'd0,(kernel[2][4] ~^ image[21][21])} + {7'd0,(kernel[3][0] ~^ image[22][17])} + {7'd0,(kernel[3][1] ~^ image[22][18])} + {7'd0,(kernel[3][2] ~^ image[22][19])} + {7'd0,(kernel[3][3] ~^ image[22][20])} + {7'd0,(kernel[3][4] ~^ image[22][21])} + {7'd0,(kernel[4][0] ~^ image[23][17])} + {7'd0,(kernel[4][1] ~^ image[23][18])} + {7'd0,(kernel[4][2] ~^ image[23][19])} + {7'd0,(kernel[4][3] ~^ image[23][20])} + {7'd0,(kernel[4][4] ~^ image[23][21])};
assign out_fmap[19][18][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[19][18])} + {7'd0,(kernel[0][1] ~^ image[19][19])} + {7'd0,(kernel[0][2] ~^ image[19][20])} + {7'd0,(kernel[0][3] ~^ image[19][21])} + {7'd0,(kernel[0][4] ~^ image[19][22])} + {7'd0,(kernel[1][0] ~^ image[20][18])} + {7'd0,(kernel[1][1] ~^ image[20][19])} + {7'd0,(kernel[1][2] ~^ image[20][20])} + {7'd0,(kernel[1][3] ~^ image[20][21])} + {7'd0,(kernel[1][4] ~^ image[20][22])} + {7'd0,(kernel[2][0] ~^ image[21][18])} + {7'd0,(kernel[2][1] ~^ image[21][19])} + {7'd0,(kernel[2][2] ~^ image[21][20])} + {7'd0,(kernel[2][3] ~^ image[21][21])} + {7'd0,(kernel[2][4] ~^ image[21][22])} + {7'd0,(kernel[3][0] ~^ image[22][18])} + {7'd0,(kernel[3][1] ~^ image[22][19])} + {7'd0,(kernel[3][2] ~^ image[22][20])} + {7'd0,(kernel[3][3] ~^ image[22][21])} + {7'd0,(kernel[3][4] ~^ image[22][22])} + {7'd0,(kernel[4][0] ~^ image[23][18])} + {7'd0,(kernel[4][1] ~^ image[23][19])} + {7'd0,(kernel[4][2] ~^ image[23][20])} + {7'd0,(kernel[4][3] ~^ image[23][21])} + {7'd0,(kernel[4][4] ~^ image[23][22])};
assign out_fmap[19][19][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[19][19])} + {7'd0,(kernel[0][1] ~^ image[19][20])} + {7'd0,(kernel[0][2] ~^ image[19][21])} + {7'd0,(kernel[0][3] ~^ image[19][22])} + {7'd0,(kernel[0][4] ~^ image[19][23])} + {7'd0,(kernel[1][0] ~^ image[20][19])} + {7'd0,(kernel[1][1] ~^ image[20][20])} + {7'd0,(kernel[1][2] ~^ image[20][21])} + {7'd0,(kernel[1][3] ~^ image[20][22])} + {7'd0,(kernel[1][4] ~^ image[20][23])} + {7'd0,(kernel[2][0] ~^ image[21][19])} + {7'd0,(kernel[2][1] ~^ image[21][20])} + {7'd0,(kernel[2][2] ~^ image[21][21])} + {7'd0,(kernel[2][3] ~^ image[21][22])} + {7'd0,(kernel[2][4] ~^ image[21][23])} + {7'd0,(kernel[3][0] ~^ image[22][19])} + {7'd0,(kernel[3][1] ~^ image[22][20])} + {7'd0,(kernel[3][2] ~^ image[22][21])} + {7'd0,(kernel[3][3] ~^ image[22][22])} + {7'd0,(kernel[3][4] ~^ image[22][23])} + {7'd0,(kernel[4][0] ~^ image[23][19])} + {7'd0,(kernel[4][1] ~^ image[23][20])} + {7'd0,(kernel[4][2] ~^ image[23][21])} + {7'd0,(kernel[4][3] ~^ image[23][22])} + {7'd0,(kernel[4][4] ~^ image[23][23])};
assign out_fmap[19][20][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[19][20])} + {7'd0,(kernel[0][1] ~^ image[19][21])} + {7'd0,(kernel[0][2] ~^ image[19][22])} + {7'd0,(kernel[0][3] ~^ image[19][23])} + {7'd0,(kernel[0][4] ~^ image[19][24])} + {7'd0,(kernel[1][0] ~^ image[20][20])} + {7'd0,(kernel[1][1] ~^ image[20][21])} + {7'd0,(kernel[1][2] ~^ image[20][22])} + {7'd0,(kernel[1][3] ~^ image[20][23])} + {7'd0,(kernel[1][4] ~^ image[20][24])} + {7'd0,(kernel[2][0] ~^ image[21][20])} + {7'd0,(kernel[2][1] ~^ image[21][21])} + {7'd0,(kernel[2][2] ~^ image[21][22])} + {7'd0,(kernel[2][3] ~^ image[21][23])} + {7'd0,(kernel[2][4] ~^ image[21][24])} + {7'd0,(kernel[3][0] ~^ image[22][20])} + {7'd0,(kernel[3][1] ~^ image[22][21])} + {7'd0,(kernel[3][2] ~^ image[22][22])} + {7'd0,(kernel[3][3] ~^ image[22][23])} + {7'd0,(kernel[3][4] ~^ image[22][24])} + {7'd0,(kernel[4][0] ~^ image[23][20])} + {7'd0,(kernel[4][1] ~^ image[23][21])} + {7'd0,(kernel[4][2] ~^ image[23][22])} + {7'd0,(kernel[4][3] ~^ image[23][23])} + {7'd0,(kernel[4][4] ~^ image[23][24])};
assign out_fmap[19][21][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[19][21])} + {7'd0,(kernel[0][1] ~^ image[19][22])} + {7'd0,(kernel[0][2] ~^ image[19][23])} + {7'd0,(kernel[0][3] ~^ image[19][24])} + {7'd0,(kernel[0][4] ~^ image[19][25])} + {7'd0,(kernel[1][0] ~^ image[20][21])} + {7'd0,(kernel[1][1] ~^ image[20][22])} + {7'd0,(kernel[1][2] ~^ image[20][23])} + {7'd0,(kernel[1][3] ~^ image[20][24])} + {7'd0,(kernel[1][4] ~^ image[20][25])} + {7'd0,(kernel[2][0] ~^ image[21][21])} + {7'd0,(kernel[2][1] ~^ image[21][22])} + {7'd0,(kernel[2][2] ~^ image[21][23])} + {7'd0,(kernel[2][3] ~^ image[21][24])} + {7'd0,(kernel[2][4] ~^ image[21][25])} + {7'd0,(kernel[3][0] ~^ image[22][21])} + {7'd0,(kernel[3][1] ~^ image[22][22])} + {7'd0,(kernel[3][2] ~^ image[22][23])} + {7'd0,(kernel[3][3] ~^ image[22][24])} + {7'd0,(kernel[3][4] ~^ image[22][25])} + {7'd0,(kernel[4][0] ~^ image[23][21])} + {7'd0,(kernel[4][1] ~^ image[23][22])} + {7'd0,(kernel[4][2] ~^ image[23][23])} + {7'd0,(kernel[4][3] ~^ image[23][24])} + {7'd0,(kernel[4][4] ~^ image[23][25])};
assign out_fmap[19][22][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[19][22])} + {7'd0,(kernel[0][1] ~^ image[19][23])} + {7'd0,(kernel[0][2] ~^ image[19][24])} + {7'd0,(kernel[0][3] ~^ image[19][25])} + {7'd0,(kernel[0][4] ~^ image[19][26])} + {7'd0,(kernel[1][0] ~^ image[20][22])} + {7'd0,(kernel[1][1] ~^ image[20][23])} + {7'd0,(kernel[1][2] ~^ image[20][24])} + {7'd0,(kernel[1][3] ~^ image[20][25])} + {7'd0,(kernel[1][4] ~^ image[20][26])} + {7'd0,(kernel[2][0] ~^ image[21][22])} + {7'd0,(kernel[2][1] ~^ image[21][23])} + {7'd0,(kernel[2][2] ~^ image[21][24])} + {7'd0,(kernel[2][3] ~^ image[21][25])} + {7'd0,(kernel[2][4] ~^ image[21][26])} + {7'd0,(kernel[3][0] ~^ image[22][22])} + {7'd0,(kernel[3][1] ~^ image[22][23])} + {7'd0,(kernel[3][2] ~^ image[22][24])} + {7'd0,(kernel[3][3] ~^ image[22][25])} + {7'd0,(kernel[3][4] ~^ image[22][26])} + {7'd0,(kernel[4][0] ~^ image[23][22])} + {7'd0,(kernel[4][1] ~^ image[23][23])} + {7'd0,(kernel[4][2] ~^ image[23][24])} + {7'd0,(kernel[4][3] ~^ image[23][25])} + {7'd0,(kernel[4][4] ~^ image[23][26])};
assign out_fmap[19][23][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[19][23])} + {7'd0,(kernel[0][1] ~^ image[19][24])} + {7'd0,(kernel[0][2] ~^ image[19][25])} + {7'd0,(kernel[0][3] ~^ image[19][26])} + {7'd0,(kernel[0][4] ~^ image[19][27])} + {7'd0,(kernel[1][0] ~^ image[20][23])} + {7'd0,(kernel[1][1] ~^ image[20][24])} + {7'd0,(kernel[1][2] ~^ image[20][25])} + {7'd0,(kernel[1][3] ~^ image[20][26])} + {7'd0,(kernel[1][4] ~^ image[20][27])} + {7'd0,(kernel[2][0] ~^ image[21][23])} + {7'd0,(kernel[2][1] ~^ image[21][24])} + {7'd0,(kernel[2][2] ~^ image[21][25])} + {7'd0,(kernel[2][3] ~^ image[21][26])} + {7'd0,(kernel[2][4] ~^ image[21][27])} + {7'd0,(kernel[3][0] ~^ image[22][23])} + {7'd0,(kernel[3][1] ~^ image[22][24])} + {7'd0,(kernel[3][2] ~^ image[22][25])} + {7'd0,(kernel[3][3] ~^ image[22][26])} + {7'd0,(kernel[3][4] ~^ image[22][27])} + {7'd0,(kernel[4][0] ~^ image[23][23])} + {7'd0,(kernel[4][1] ~^ image[23][24])} + {7'd0,(kernel[4][2] ~^ image[23][25])} + {7'd0,(kernel[4][3] ~^ image[23][26])} + {7'd0,(kernel[4][4] ~^ image[23][27])};
assign out_fmap[20][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[20][0])} + {7'd0,(kernel[0][1] ~^ image[20][1])} + {7'd0,(kernel[0][2] ~^ image[20][2])} + {7'd0,(kernel[0][3] ~^ image[20][3])} + {7'd0,(kernel[0][4] ~^ image[20][4])} + {7'd0,(kernel[1][0] ~^ image[21][0])} + {7'd0,(kernel[1][1] ~^ image[21][1])} + {7'd0,(kernel[1][2] ~^ image[21][2])} + {7'd0,(kernel[1][3] ~^ image[21][3])} + {7'd0,(kernel[1][4] ~^ image[21][4])} + {7'd0,(kernel[2][0] ~^ image[22][0])} + {7'd0,(kernel[2][1] ~^ image[22][1])} + {7'd0,(kernel[2][2] ~^ image[22][2])} + {7'd0,(kernel[2][3] ~^ image[22][3])} + {7'd0,(kernel[2][4] ~^ image[22][4])} + {7'd0,(kernel[3][0] ~^ image[23][0])} + {7'd0,(kernel[3][1] ~^ image[23][1])} + {7'd0,(kernel[3][2] ~^ image[23][2])} + {7'd0,(kernel[3][3] ~^ image[23][3])} + {7'd0,(kernel[3][4] ~^ image[23][4])} + {7'd0,(kernel[4][0] ~^ image[24][0])} + {7'd0,(kernel[4][1] ~^ image[24][1])} + {7'd0,(kernel[4][2] ~^ image[24][2])} + {7'd0,(kernel[4][3] ~^ image[24][3])} + {7'd0,(kernel[4][4] ~^ image[24][4])};
assign out_fmap[20][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[20][1])} + {7'd0,(kernel[0][1] ~^ image[20][2])} + {7'd0,(kernel[0][2] ~^ image[20][3])} + {7'd0,(kernel[0][3] ~^ image[20][4])} + {7'd0,(kernel[0][4] ~^ image[20][5])} + {7'd0,(kernel[1][0] ~^ image[21][1])} + {7'd0,(kernel[1][1] ~^ image[21][2])} + {7'd0,(kernel[1][2] ~^ image[21][3])} + {7'd0,(kernel[1][3] ~^ image[21][4])} + {7'd0,(kernel[1][4] ~^ image[21][5])} + {7'd0,(kernel[2][0] ~^ image[22][1])} + {7'd0,(kernel[2][1] ~^ image[22][2])} + {7'd0,(kernel[2][2] ~^ image[22][3])} + {7'd0,(kernel[2][3] ~^ image[22][4])} + {7'd0,(kernel[2][4] ~^ image[22][5])} + {7'd0,(kernel[3][0] ~^ image[23][1])} + {7'd0,(kernel[3][1] ~^ image[23][2])} + {7'd0,(kernel[3][2] ~^ image[23][3])} + {7'd0,(kernel[3][3] ~^ image[23][4])} + {7'd0,(kernel[3][4] ~^ image[23][5])} + {7'd0,(kernel[4][0] ~^ image[24][1])} + {7'd0,(kernel[4][1] ~^ image[24][2])} + {7'd0,(kernel[4][2] ~^ image[24][3])} + {7'd0,(kernel[4][3] ~^ image[24][4])} + {7'd0,(kernel[4][4] ~^ image[24][5])};
assign out_fmap[20][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[20][2])} + {7'd0,(kernel[0][1] ~^ image[20][3])} + {7'd0,(kernel[0][2] ~^ image[20][4])} + {7'd0,(kernel[0][3] ~^ image[20][5])} + {7'd0,(kernel[0][4] ~^ image[20][6])} + {7'd0,(kernel[1][0] ~^ image[21][2])} + {7'd0,(kernel[1][1] ~^ image[21][3])} + {7'd0,(kernel[1][2] ~^ image[21][4])} + {7'd0,(kernel[1][3] ~^ image[21][5])} + {7'd0,(kernel[1][4] ~^ image[21][6])} + {7'd0,(kernel[2][0] ~^ image[22][2])} + {7'd0,(kernel[2][1] ~^ image[22][3])} + {7'd0,(kernel[2][2] ~^ image[22][4])} + {7'd0,(kernel[2][3] ~^ image[22][5])} + {7'd0,(kernel[2][4] ~^ image[22][6])} + {7'd0,(kernel[3][0] ~^ image[23][2])} + {7'd0,(kernel[3][1] ~^ image[23][3])} + {7'd0,(kernel[3][2] ~^ image[23][4])} + {7'd0,(kernel[3][3] ~^ image[23][5])} + {7'd0,(kernel[3][4] ~^ image[23][6])} + {7'd0,(kernel[4][0] ~^ image[24][2])} + {7'd0,(kernel[4][1] ~^ image[24][3])} + {7'd0,(kernel[4][2] ~^ image[24][4])} + {7'd0,(kernel[4][3] ~^ image[24][5])} + {7'd0,(kernel[4][4] ~^ image[24][6])};
assign out_fmap[20][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[20][3])} + {7'd0,(kernel[0][1] ~^ image[20][4])} + {7'd0,(kernel[0][2] ~^ image[20][5])} + {7'd0,(kernel[0][3] ~^ image[20][6])} + {7'd0,(kernel[0][4] ~^ image[20][7])} + {7'd0,(kernel[1][0] ~^ image[21][3])} + {7'd0,(kernel[1][1] ~^ image[21][4])} + {7'd0,(kernel[1][2] ~^ image[21][5])} + {7'd0,(kernel[1][3] ~^ image[21][6])} + {7'd0,(kernel[1][4] ~^ image[21][7])} + {7'd0,(kernel[2][0] ~^ image[22][3])} + {7'd0,(kernel[2][1] ~^ image[22][4])} + {7'd0,(kernel[2][2] ~^ image[22][5])} + {7'd0,(kernel[2][3] ~^ image[22][6])} + {7'd0,(kernel[2][4] ~^ image[22][7])} + {7'd0,(kernel[3][0] ~^ image[23][3])} + {7'd0,(kernel[3][1] ~^ image[23][4])} + {7'd0,(kernel[3][2] ~^ image[23][5])} + {7'd0,(kernel[3][3] ~^ image[23][6])} + {7'd0,(kernel[3][4] ~^ image[23][7])} + {7'd0,(kernel[4][0] ~^ image[24][3])} + {7'd0,(kernel[4][1] ~^ image[24][4])} + {7'd0,(kernel[4][2] ~^ image[24][5])} + {7'd0,(kernel[4][3] ~^ image[24][6])} + {7'd0,(kernel[4][4] ~^ image[24][7])};
assign out_fmap[20][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[20][4])} + {7'd0,(kernel[0][1] ~^ image[20][5])} + {7'd0,(kernel[0][2] ~^ image[20][6])} + {7'd0,(kernel[0][3] ~^ image[20][7])} + {7'd0,(kernel[0][4] ~^ image[20][8])} + {7'd0,(kernel[1][0] ~^ image[21][4])} + {7'd0,(kernel[1][1] ~^ image[21][5])} + {7'd0,(kernel[1][2] ~^ image[21][6])} + {7'd0,(kernel[1][3] ~^ image[21][7])} + {7'd0,(kernel[1][4] ~^ image[21][8])} + {7'd0,(kernel[2][0] ~^ image[22][4])} + {7'd0,(kernel[2][1] ~^ image[22][5])} + {7'd0,(kernel[2][2] ~^ image[22][6])} + {7'd0,(kernel[2][3] ~^ image[22][7])} + {7'd0,(kernel[2][4] ~^ image[22][8])} + {7'd0,(kernel[3][0] ~^ image[23][4])} + {7'd0,(kernel[3][1] ~^ image[23][5])} + {7'd0,(kernel[3][2] ~^ image[23][6])} + {7'd0,(kernel[3][3] ~^ image[23][7])} + {7'd0,(kernel[3][4] ~^ image[23][8])} + {7'd0,(kernel[4][0] ~^ image[24][4])} + {7'd0,(kernel[4][1] ~^ image[24][5])} + {7'd0,(kernel[4][2] ~^ image[24][6])} + {7'd0,(kernel[4][3] ~^ image[24][7])} + {7'd0,(kernel[4][4] ~^ image[24][8])};
assign out_fmap[20][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[20][5])} + {7'd0,(kernel[0][1] ~^ image[20][6])} + {7'd0,(kernel[0][2] ~^ image[20][7])} + {7'd0,(kernel[0][3] ~^ image[20][8])} + {7'd0,(kernel[0][4] ~^ image[20][9])} + {7'd0,(kernel[1][0] ~^ image[21][5])} + {7'd0,(kernel[1][1] ~^ image[21][6])} + {7'd0,(kernel[1][2] ~^ image[21][7])} + {7'd0,(kernel[1][3] ~^ image[21][8])} + {7'd0,(kernel[1][4] ~^ image[21][9])} + {7'd0,(kernel[2][0] ~^ image[22][5])} + {7'd0,(kernel[2][1] ~^ image[22][6])} + {7'd0,(kernel[2][2] ~^ image[22][7])} + {7'd0,(kernel[2][3] ~^ image[22][8])} + {7'd0,(kernel[2][4] ~^ image[22][9])} + {7'd0,(kernel[3][0] ~^ image[23][5])} + {7'd0,(kernel[3][1] ~^ image[23][6])} + {7'd0,(kernel[3][2] ~^ image[23][7])} + {7'd0,(kernel[3][3] ~^ image[23][8])} + {7'd0,(kernel[3][4] ~^ image[23][9])} + {7'd0,(kernel[4][0] ~^ image[24][5])} + {7'd0,(kernel[4][1] ~^ image[24][6])} + {7'd0,(kernel[4][2] ~^ image[24][7])} + {7'd0,(kernel[4][3] ~^ image[24][8])} + {7'd0,(kernel[4][4] ~^ image[24][9])};
assign out_fmap[20][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[20][6])} + {7'd0,(kernel[0][1] ~^ image[20][7])} + {7'd0,(kernel[0][2] ~^ image[20][8])} + {7'd0,(kernel[0][3] ~^ image[20][9])} + {7'd0,(kernel[0][4] ~^ image[20][10])} + {7'd0,(kernel[1][0] ~^ image[21][6])} + {7'd0,(kernel[1][1] ~^ image[21][7])} + {7'd0,(kernel[1][2] ~^ image[21][8])} + {7'd0,(kernel[1][3] ~^ image[21][9])} + {7'd0,(kernel[1][4] ~^ image[21][10])} + {7'd0,(kernel[2][0] ~^ image[22][6])} + {7'd0,(kernel[2][1] ~^ image[22][7])} + {7'd0,(kernel[2][2] ~^ image[22][8])} + {7'd0,(kernel[2][3] ~^ image[22][9])} + {7'd0,(kernel[2][4] ~^ image[22][10])} + {7'd0,(kernel[3][0] ~^ image[23][6])} + {7'd0,(kernel[3][1] ~^ image[23][7])} + {7'd0,(kernel[3][2] ~^ image[23][8])} + {7'd0,(kernel[3][3] ~^ image[23][9])} + {7'd0,(kernel[3][4] ~^ image[23][10])} + {7'd0,(kernel[4][0] ~^ image[24][6])} + {7'd0,(kernel[4][1] ~^ image[24][7])} + {7'd0,(kernel[4][2] ~^ image[24][8])} + {7'd0,(kernel[4][3] ~^ image[24][9])} + {7'd0,(kernel[4][4] ~^ image[24][10])};
assign out_fmap[20][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[20][7])} + {7'd0,(kernel[0][1] ~^ image[20][8])} + {7'd0,(kernel[0][2] ~^ image[20][9])} + {7'd0,(kernel[0][3] ~^ image[20][10])} + {7'd0,(kernel[0][4] ~^ image[20][11])} + {7'd0,(kernel[1][0] ~^ image[21][7])} + {7'd0,(kernel[1][1] ~^ image[21][8])} + {7'd0,(kernel[1][2] ~^ image[21][9])} + {7'd0,(kernel[1][3] ~^ image[21][10])} + {7'd0,(kernel[1][4] ~^ image[21][11])} + {7'd0,(kernel[2][0] ~^ image[22][7])} + {7'd0,(kernel[2][1] ~^ image[22][8])} + {7'd0,(kernel[2][2] ~^ image[22][9])} + {7'd0,(kernel[2][3] ~^ image[22][10])} + {7'd0,(kernel[2][4] ~^ image[22][11])} + {7'd0,(kernel[3][0] ~^ image[23][7])} + {7'd0,(kernel[3][1] ~^ image[23][8])} + {7'd0,(kernel[3][2] ~^ image[23][9])} + {7'd0,(kernel[3][3] ~^ image[23][10])} + {7'd0,(kernel[3][4] ~^ image[23][11])} + {7'd0,(kernel[4][0] ~^ image[24][7])} + {7'd0,(kernel[4][1] ~^ image[24][8])} + {7'd0,(kernel[4][2] ~^ image[24][9])} + {7'd0,(kernel[4][3] ~^ image[24][10])} + {7'd0,(kernel[4][4] ~^ image[24][11])};
assign out_fmap[20][8][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[20][8])} + {7'd0,(kernel[0][1] ~^ image[20][9])} + {7'd0,(kernel[0][2] ~^ image[20][10])} + {7'd0,(kernel[0][3] ~^ image[20][11])} + {7'd0,(kernel[0][4] ~^ image[20][12])} + {7'd0,(kernel[1][0] ~^ image[21][8])} + {7'd0,(kernel[1][1] ~^ image[21][9])} + {7'd0,(kernel[1][2] ~^ image[21][10])} + {7'd0,(kernel[1][3] ~^ image[21][11])} + {7'd0,(kernel[1][4] ~^ image[21][12])} + {7'd0,(kernel[2][0] ~^ image[22][8])} + {7'd0,(kernel[2][1] ~^ image[22][9])} + {7'd0,(kernel[2][2] ~^ image[22][10])} + {7'd0,(kernel[2][3] ~^ image[22][11])} + {7'd0,(kernel[2][4] ~^ image[22][12])} + {7'd0,(kernel[3][0] ~^ image[23][8])} + {7'd0,(kernel[3][1] ~^ image[23][9])} + {7'd0,(kernel[3][2] ~^ image[23][10])} + {7'd0,(kernel[3][3] ~^ image[23][11])} + {7'd0,(kernel[3][4] ~^ image[23][12])} + {7'd0,(kernel[4][0] ~^ image[24][8])} + {7'd0,(kernel[4][1] ~^ image[24][9])} + {7'd0,(kernel[4][2] ~^ image[24][10])} + {7'd0,(kernel[4][3] ~^ image[24][11])} + {7'd0,(kernel[4][4] ~^ image[24][12])};
assign out_fmap[20][9][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[20][9])} + {7'd0,(kernel[0][1] ~^ image[20][10])} + {7'd0,(kernel[0][2] ~^ image[20][11])} + {7'd0,(kernel[0][3] ~^ image[20][12])} + {7'd0,(kernel[0][4] ~^ image[20][13])} + {7'd0,(kernel[1][0] ~^ image[21][9])} + {7'd0,(kernel[1][1] ~^ image[21][10])} + {7'd0,(kernel[1][2] ~^ image[21][11])} + {7'd0,(kernel[1][3] ~^ image[21][12])} + {7'd0,(kernel[1][4] ~^ image[21][13])} + {7'd0,(kernel[2][0] ~^ image[22][9])} + {7'd0,(kernel[2][1] ~^ image[22][10])} + {7'd0,(kernel[2][2] ~^ image[22][11])} + {7'd0,(kernel[2][3] ~^ image[22][12])} + {7'd0,(kernel[2][4] ~^ image[22][13])} + {7'd0,(kernel[3][0] ~^ image[23][9])} + {7'd0,(kernel[3][1] ~^ image[23][10])} + {7'd0,(kernel[3][2] ~^ image[23][11])} + {7'd0,(kernel[3][3] ~^ image[23][12])} + {7'd0,(kernel[3][4] ~^ image[23][13])} + {7'd0,(kernel[4][0] ~^ image[24][9])} + {7'd0,(kernel[4][1] ~^ image[24][10])} + {7'd0,(kernel[4][2] ~^ image[24][11])} + {7'd0,(kernel[4][3] ~^ image[24][12])} + {7'd0,(kernel[4][4] ~^ image[24][13])};
assign out_fmap[20][10][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[20][10])} + {7'd0,(kernel[0][1] ~^ image[20][11])} + {7'd0,(kernel[0][2] ~^ image[20][12])} + {7'd0,(kernel[0][3] ~^ image[20][13])} + {7'd0,(kernel[0][4] ~^ image[20][14])} + {7'd0,(kernel[1][0] ~^ image[21][10])} + {7'd0,(kernel[1][1] ~^ image[21][11])} + {7'd0,(kernel[1][2] ~^ image[21][12])} + {7'd0,(kernel[1][3] ~^ image[21][13])} + {7'd0,(kernel[1][4] ~^ image[21][14])} + {7'd0,(kernel[2][0] ~^ image[22][10])} + {7'd0,(kernel[2][1] ~^ image[22][11])} + {7'd0,(kernel[2][2] ~^ image[22][12])} + {7'd0,(kernel[2][3] ~^ image[22][13])} + {7'd0,(kernel[2][4] ~^ image[22][14])} + {7'd0,(kernel[3][0] ~^ image[23][10])} + {7'd0,(kernel[3][1] ~^ image[23][11])} + {7'd0,(kernel[3][2] ~^ image[23][12])} + {7'd0,(kernel[3][3] ~^ image[23][13])} + {7'd0,(kernel[3][4] ~^ image[23][14])} + {7'd0,(kernel[4][0] ~^ image[24][10])} + {7'd0,(kernel[4][1] ~^ image[24][11])} + {7'd0,(kernel[4][2] ~^ image[24][12])} + {7'd0,(kernel[4][3] ~^ image[24][13])} + {7'd0,(kernel[4][4] ~^ image[24][14])};
assign out_fmap[20][11][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[20][11])} + {7'd0,(kernel[0][1] ~^ image[20][12])} + {7'd0,(kernel[0][2] ~^ image[20][13])} + {7'd0,(kernel[0][3] ~^ image[20][14])} + {7'd0,(kernel[0][4] ~^ image[20][15])} + {7'd0,(kernel[1][0] ~^ image[21][11])} + {7'd0,(kernel[1][1] ~^ image[21][12])} + {7'd0,(kernel[1][2] ~^ image[21][13])} + {7'd0,(kernel[1][3] ~^ image[21][14])} + {7'd0,(kernel[1][4] ~^ image[21][15])} + {7'd0,(kernel[2][0] ~^ image[22][11])} + {7'd0,(kernel[2][1] ~^ image[22][12])} + {7'd0,(kernel[2][2] ~^ image[22][13])} + {7'd0,(kernel[2][3] ~^ image[22][14])} + {7'd0,(kernel[2][4] ~^ image[22][15])} + {7'd0,(kernel[3][0] ~^ image[23][11])} + {7'd0,(kernel[3][1] ~^ image[23][12])} + {7'd0,(kernel[3][2] ~^ image[23][13])} + {7'd0,(kernel[3][3] ~^ image[23][14])} + {7'd0,(kernel[3][4] ~^ image[23][15])} + {7'd0,(kernel[4][0] ~^ image[24][11])} + {7'd0,(kernel[4][1] ~^ image[24][12])} + {7'd0,(kernel[4][2] ~^ image[24][13])} + {7'd0,(kernel[4][3] ~^ image[24][14])} + {7'd0,(kernel[4][4] ~^ image[24][15])};
assign out_fmap[20][12][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[20][12])} + {7'd0,(kernel[0][1] ~^ image[20][13])} + {7'd0,(kernel[0][2] ~^ image[20][14])} + {7'd0,(kernel[0][3] ~^ image[20][15])} + {7'd0,(kernel[0][4] ~^ image[20][16])} + {7'd0,(kernel[1][0] ~^ image[21][12])} + {7'd0,(kernel[1][1] ~^ image[21][13])} + {7'd0,(kernel[1][2] ~^ image[21][14])} + {7'd0,(kernel[1][3] ~^ image[21][15])} + {7'd0,(kernel[1][4] ~^ image[21][16])} + {7'd0,(kernel[2][0] ~^ image[22][12])} + {7'd0,(kernel[2][1] ~^ image[22][13])} + {7'd0,(kernel[2][2] ~^ image[22][14])} + {7'd0,(kernel[2][3] ~^ image[22][15])} + {7'd0,(kernel[2][4] ~^ image[22][16])} + {7'd0,(kernel[3][0] ~^ image[23][12])} + {7'd0,(kernel[3][1] ~^ image[23][13])} + {7'd0,(kernel[3][2] ~^ image[23][14])} + {7'd0,(kernel[3][3] ~^ image[23][15])} + {7'd0,(kernel[3][4] ~^ image[23][16])} + {7'd0,(kernel[4][0] ~^ image[24][12])} + {7'd0,(kernel[4][1] ~^ image[24][13])} + {7'd0,(kernel[4][2] ~^ image[24][14])} + {7'd0,(kernel[4][3] ~^ image[24][15])} + {7'd0,(kernel[4][4] ~^ image[24][16])};
assign out_fmap[20][13][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[20][13])} + {7'd0,(kernel[0][1] ~^ image[20][14])} + {7'd0,(kernel[0][2] ~^ image[20][15])} + {7'd0,(kernel[0][3] ~^ image[20][16])} + {7'd0,(kernel[0][4] ~^ image[20][17])} + {7'd0,(kernel[1][0] ~^ image[21][13])} + {7'd0,(kernel[1][1] ~^ image[21][14])} + {7'd0,(kernel[1][2] ~^ image[21][15])} + {7'd0,(kernel[1][3] ~^ image[21][16])} + {7'd0,(kernel[1][4] ~^ image[21][17])} + {7'd0,(kernel[2][0] ~^ image[22][13])} + {7'd0,(kernel[2][1] ~^ image[22][14])} + {7'd0,(kernel[2][2] ~^ image[22][15])} + {7'd0,(kernel[2][3] ~^ image[22][16])} + {7'd0,(kernel[2][4] ~^ image[22][17])} + {7'd0,(kernel[3][0] ~^ image[23][13])} + {7'd0,(kernel[3][1] ~^ image[23][14])} + {7'd0,(kernel[3][2] ~^ image[23][15])} + {7'd0,(kernel[3][3] ~^ image[23][16])} + {7'd0,(kernel[3][4] ~^ image[23][17])} + {7'd0,(kernel[4][0] ~^ image[24][13])} + {7'd0,(kernel[4][1] ~^ image[24][14])} + {7'd0,(kernel[4][2] ~^ image[24][15])} + {7'd0,(kernel[4][3] ~^ image[24][16])} + {7'd0,(kernel[4][4] ~^ image[24][17])};
assign out_fmap[20][14][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[20][14])} + {7'd0,(kernel[0][1] ~^ image[20][15])} + {7'd0,(kernel[0][2] ~^ image[20][16])} + {7'd0,(kernel[0][3] ~^ image[20][17])} + {7'd0,(kernel[0][4] ~^ image[20][18])} + {7'd0,(kernel[1][0] ~^ image[21][14])} + {7'd0,(kernel[1][1] ~^ image[21][15])} + {7'd0,(kernel[1][2] ~^ image[21][16])} + {7'd0,(kernel[1][3] ~^ image[21][17])} + {7'd0,(kernel[1][4] ~^ image[21][18])} + {7'd0,(kernel[2][0] ~^ image[22][14])} + {7'd0,(kernel[2][1] ~^ image[22][15])} + {7'd0,(kernel[2][2] ~^ image[22][16])} + {7'd0,(kernel[2][3] ~^ image[22][17])} + {7'd0,(kernel[2][4] ~^ image[22][18])} + {7'd0,(kernel[3][0] ~^ image[23][14])} + {7'd0,(kernel[3][1] ~^ image[23][15])} + {7'd0,(kernel[3][2] ~^ image[23][16])} + {7'd0,(kernel[3][3] ~^ image[23][17])} + {7'd0,(kernel[3][4] ~^ image[23][18])} + {7'd0,(kernel[4][0] ~^ image[24][14])} + {7'd0,(kernel[4][1] ~^ image[24][15])} + {7'd0,(kernel[4][2] ~^ image[24][16])} + {7'd0,(kernel[4][3] ~^ image[24][17])} + {7'd0,(kernel[4][4] ~^ image[24][18])};
assign out_fmap[20][15][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[20][15])} + {7'd0,(kernel[0][1] ~^ image[20][16])} + {7'd0,(kernel[0][2] ~^ image[20][17])} + {7'd0,(kernel[0][3] ~^ image[20][18])} + {7'd0,(kernel[0][4] ~^ image[20][19])} + {7'd0,(kernel[1][0] ~^ image[21][15])} + {7'd0,(kernel[1][1] ~^ image[21][16])} + {7'd0,(kernel[1][2] ~^ image[21][17])} + {7'd0,(kernel[1][3] ~^ image[21][18])} + {7'd0,(kernel[1][4] ~^ image[21][19])} + {7'd0,(kernel[2][0] ~^ image[22][15])} + {7'd0,(kernel[2][1] ~^ image[22][16])} + {7'd0,(kernel[2][2] ~^ image[22][17])} + {7'd0,(kernel[2][3] ~^ image[22][18])} + {7'd0,(kernel[2][4] ~^ image[22][19])} + {7'd0,(kernel[3][0] ~^ image[23][15])} + {7'd0,(kernel[3][1] ~^ image[23][16])} + {7'd0,(kernel[3][2] ~^ image[23][17])} + {7'd0,(kernel[3][3] ~^ image[23][18])} + {7'd0,(kernel[3][4] ~^ image[23][19])} + {7'd0,(kernel[4][0] ~^ image[24][15])} + {7'd0,(kernel[4][1] ~^ image[24][16])} + {7'd0,(kernel[4][2] ~^ image[24][17])} + {7'd0,(kernel[4][3] ~^ image[24][18])} + {7'd0,(kernel[4][4] ~^ image[24][19])};
assign out_fmap[20][16][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[20][16])} + {7'd0,(kernel[0][1] ~^ image[20][17])} + {7'd0,(kernel[0][2] ~^ image[20][18])} + {7'd0,(kernel[0][3] ~^ image[20][19])} + {7'd0,(kernel[0][4] ~^ image[20][20])} + {7'd0,(kernel[1][0] ~^ image[21][16])} + {7'd0,(kernel[1][1] ~^ image[21][17])} + {7'd0,(kernel[1][2] ~^ image[21][18])} + {7'd0,(kernel[1][3] ~^ image[21][19])} + {7'd0,(kernel[1][4] ~^ image[21][20])} + {7'd0,(kernel[2][0] ~^ image[22][16])} + {7'd0,(kernel[2][1] ~^ image[22][17])} + {7'd0,(kernel[2][2] ~^ image[22][18])} + {7'd0,(kernel[2][3] ~^ image[22][19])} + {7'd0,(kernel[2][4] ~^ image[22][20])} + {7'd0,(kernel[3][0] ~^ image[23][16])} + {7'd0,(kernel[3][1] ~^ image[23][17])} + {7'd0,(kernel[3][2] ~^ image[23][18])} + {7'd0,(kernel[3][3] ~^ image[23][19])} + {7'd0,(kernel[3][4] ~^ image[23][20])} + {7'd0,(kernel[4][0] ~^ image[24][16])} + {7'd0,(kernel[4][1] ~^ image[24][17])} + {7'd0,(kernel[4][2] ~^ image[24][18])} + {7'd0,(kernel[4][3] ~^ image[24][19])} + {7'd0,(kernel[4][4] ~^ image[24][20])};
assign out_fmap[20][17][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[20][17])} + {7'd0,(kernel[0][1] ~^ image[20][18])} + {7'd0,(kernel[0][2] ~^ image[20][19])} + {7'd0,(kernel[0][3] ~^ image[20][20])} + {7'd0,(kernel[0][4] ~^ image[20][21])} + {7'd0,(kernel[1][0] ~^ image[21][17])} + {7'd0,(kernel[1][1] ~^ image[21][18])} + {7'd0,(kernel[1][2] ~^ image[21][19])} + {7'd0,(kernel[1][3] ~^ image[21][20])} + {7'd0,(kernel[1][4] ~^ image[21][21])} + {7'd0,(kernel[2][0] ~^ image[22][17])} + {7'd0,(kernel[2][1] ~^ image[22][18])} + {7'd0,(kernel[2][2] ~^ image[22][19])} + {7'd0,(kernel[2][3] ~^ image[22][20])} + {7'd0,(kernel[2][4] ~^ image[22][21])} + {7'd0,(kernel[3][0] ~^ image[23][17])} + {7'd0,(kernel[3][1] ~^ image[23][18])} + {7'd0,(kernel[3][2] ~^ image[23][19])} + {7'd0,(kernel[3][3] ~^ image[23][20])} + {7'd0,(kernel[3][4] ~^ image[23][21])} + {7'd0,(kernel[4][0] ~^ image[24][17])} + {7'd0,(kernel[4][1] ~^ image[24][18])} + {7'd0,(kernel[4][2] ~^ image[24][19])} + {7'd0,(kernel[4][3] ~^ image[24][20])} + {7'd0,(kernel[4][4] ~^ image[24][21])};
assign out_fmap[20][18][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[20][18])} + {7'd0,(kernel[0][1] ~^ image[20][19])} + {7'd0,(kernel[0][2] ~^ image[20][20])} + {7'd0,(kernel[0][3] ~^ image[20][21])} + {7'd0,(kernel[0][4] ~^ image[20][22])} + {7'd0,(kernel[1][0] ~^ image[21][18])} + {7'd0,(kernel[1][1] ~^ image[21][19])} + {7'd0,(kernel[1][2] ~^ image[21][20])} + {7'd0,(kernel[1][3] ~^ image[21][21])} + {7'd0,(kernel[1][4] ~^ image[21][22])} + {7'd0,(kernel[2][0] ~^ image[22][18])} + {7'd0,(kernel[2][1] ~^ image[22][19])} + {7'd0,(kernel[2][2] ~^ image[22][20])} + {7'd0,(kernel[2][3] ~^ image[22][21])} + {7'd0,(kernel[2][4] ~^ image[22][22])} + {7'd0,(kernel[3][0] ~^ image[23][18])} + {7'd0,(kernel[3][1] ~^ image[23][19])} + {7'd0,(kernel[3][2] ~^ image[23][20])} + {7'd0,(kernel[3][3] ~^ image[23][21])} + {7'd0,(kernel[3][4] ~^ image[23][22])} + {7'd0,(kernel[4][0] ~^ image[24][18])} + {7'd0,(kernel[4][1] ~^ image[24][19])} + {7'd0,(kernel[4][2] ~^ image[24][20])} + {7'd0,(kernel[4][3] ~^ image[24][21])} + {7'd0,(kernel[4][4] ~^ image[24][22])};
assign out_fmap[20][19][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[20][19])} + {7'd0,(kernel[0][1] ~^ image[20][20])} + {7'd0,(kernel[0][2] ~^ image[20][21])} + {7'd0,(kernel[0][3] ~^ image[20][22])} + {7'd0,(kernel[0][4] ~^ image[20][23])} + {7'd0,(kernel[1][0] ~^ image[21][19])} + {7'd0,(kernel[1][1] ~^ image[21][20])} + {7'd0,(kernel[1][2] ~^ image[21][21])} + {7'd0,(kernel[1][3] ~^ image[21][22])} + {7'd0,(kernel[1][4] ~^ image[21][23])} + {7'd0,(kernel[2][0] ~^ image[22][19])} + {7'd0,(kernel[2][1] ~^ image[22][20])} + {7'd0,(kernel[2][2] ~^ image[22][21])} + {7'd0,(kernel[2][3] ~^ image[22][22])} + {7'd0,(kernel[2][4] ~^ image[22][23])} + {7'd0,(kernel[3][0] ~^ image[23][19])} + {7'd0,(kernel[3][1] ~^ image[23][20])} + {7'd0,(kernel[3][2] ~^ image[23][21])} + {7'd0,(kernel[3][3] ~^ image[23][22])} + {7'd0,(kernel[3][4] ~^ image[23][23])} + {7'd0,(kernel[4][0] ~^ image[24][19])} + {7'd0,(kernel[4][1] ~^ image[24][20])} + {7'd0,(kernel[4][2] ~^ image[24][21])} + {7'd0,(kernel[4][3] ~^ image[24][22])} + {7'd0,(kernel[4][4] ~^ image[24][23])};
assign out_fmap[20][20][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[20][20])} + {7'd0,(kernel[0][1] ~^ image[20][21])} + {7'd0,(kernel[0][2] ~^ image[20][22])} + {7'd0,(kernel[0][3] ~^ image[20][23])} + {7'd0,(kernel[0][4] ~^ image[20][24])} + {7'd0,(kernel[1][0] ~^ image[21][20])} + {7'd0,(kernel[1][1] ~^ image[21][21])} + {7'd0,(kernel[1][2] ~^ image[21][22])} + {7'd0,(kernel[1][3] ~^ image[21][23])} + {7'd0,(kernel[1][4] ~^ image[21][24])} + {7'd0,(kernel[2][0] ~^ image[22][20])} + {7'd0,(kernel[2][1] ~^ image[22][21])} + {7'd0,(kernel[2][2] ~^ image[22][22])} + {7'd0,(kernel[2][3] ~^ image[22][23])} + {7'd0,(kernel[2][4] ~^ image[22][24])} + {7'd0,(kernel[3][0] ~^ image[23][20])} + {7'd0,(kernel[3][1] ~^ image[23][21])} + {7'd0,(kernel[3][2] ~^ image[23][22])} + {7'd0,(kernel[3][3] ~^ image[23][23])} + {7'd0,(kernel[3][4] ~^ image[23][24])} + {7'd0,(kernel[4][0] ~^ image[24][20])} + {7'd0,(kernel[4][1] ~^ image[24][21])} + {7'd0,(kernel[4][2] ~^ image[24][22])} + {7'd0,(kernel[4][3] ~^ image[24][23])} + {7'd0,(kernel[4][4] ~^ image[24][24])};
assign out_fmap[20][21][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[20][21])} + {7'd0,(kernel[0][1] ~^ image[20][22])} + {7'd0,(kernel[0][2] ~^ image[20][23])} + {7'd0,(kernel[0][3] ~^ image[20][24])} + {7'd0,(kernel[0][4] ~^ image[20][25])} + {7'd0,(kernel[1][0] ~^ image[21][21])} + {7'd0,(kernel[1][1] ~^ image[21][22])} + {7'd0,(kernel[1][2] ~^ image[21][23])} + {7'd0,(kernel[1][3] ~^ image[21][24])} + {7'd0,(kernel[1][4] ~^ image[21][25])} + {7'd0,(kernel[2][0] ~^ image[22][21])} + {7'd0,(kernel[2][1] ~^ image[22][22])} + {7'd0,(kernel[2][2] ~^ image[22][23])} + {7'd0,(kernel[2][3] ~^ image[22][24])} + {7'd0,(kernel[2][4] ~^ image[22][25])} + {7'd0,(kernel[3][0] ~^ image[23][21])} + {7'd0,(kernel[3][1] ~^ image[23][22])} + {7'd0,(kernel[3][2] ~^ image[23][23])} + {7'd0,(kernel[3][3] ~^ image[23][24])} + {7'd0,(kernel[3][4] ~^ image[23][25])} + {7'd0,(kernel[4][0] ~^ image[24][21])} + {7'd0,(kernel[4][1] ~^ image[24][22])} + {7'd0,(kernel[4][2] ~^ image[24][23])} + {7'd0,(kernel[4][3] ~^ image[24][24])} + {7'd0,(kernel[4][4] ~^ image[24][25])};
assign out_fmap[20][22][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[20][22])} + {7'd0,(kernel[0][1] ~^ image[20][23])} + {7'd0,(kernel[0][2] ~^ image[20][24])} + {7'd0,(kernel[0][3] ~^ image[20][25])} + {7'd0,(kernel[0][4] ~^ image[20][26])} + {7'd0,(kernel[1][0] ~^ image[21][22])} + {7'd0,(kernel[1][1] ~^ image[21][23])} + {7'd0,(kernel[1][2] ~^ image[21][24])} + {7'd0,(kernel[1][3] ~^ image[21][25])} + {7'd0,(kernel[1][4] ~^ image[21][26])} + {7'd0,(kernel[2][0] ~^ image[22][22])} + {7'd0,(kernel[2][1] ~^ image[22][23])} + {7'd0,(kernel[2][2] ~^ image[22][24])} + {7'd0,(kernel[2][3] ~^ image[22][25])} + {7'd0,(kernel[2][4] ~^ image[22][26])} + {7'd0,(kernel[3][0] ~^ image[23][22])} + {7'd0,(kernel[3][1] ~^ image[23][23])} + {7'd0,(kernel[3][2] ~^ image[23][24])} + {7'd0,(kernel[3][3] ~^ image[23][25])} + {7'd0,(kernel[3][4] ~^ image[23][26])} + {7'd0,(kernel[4][0] ~^ image[24][22])} + {7'd0,(kernel[4][1] ~^ image[24][23])} + {7'd0,(kernel[4][2] ~^ image[24][24])} + {7'd0,(kernel[4][3] ~^ image[24][25])} + {7'd0,(kernel[4][4] ~^ image[24][26])};
assign out_fmap[20][23][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[20][23])} + {7'd0,(kernel[0][1] ~^ image[20][24])} + {7'd0,(kernel[0][2] ~^ image[20][25])} + {7'd0,(kernel[0][3] ~^ image[20][26])} + {7'd0,(kernel[0][4] ~^ image[20][27])} + {7'd0,(kernel[1][0] ~^ image[21][23])} + {7'd0,(kernel[1][1] ~^ image[21][24])} + {7'd0,(kernel[1][2] ~^ image[21][25])} + {7'd0,(kernel[1][3] ~^ image[21][26])} + {7'd0,(kernel[1][4] ~^ image[21][27])} + {7'd0,(kernel[2][0] ~^ image[22][23])} + {7'd0,(kernel[2][1] ~^ image[22][24])} + {7'd0,(kernel[2][2] ~^ image[22][25])} + {7'd0,(kernel[2][3] ~^ image[22][26])} + {7'd0,(kernel[2][4] ~^ image[22][27])} + {7'd0,(kernel[3][0] ~^ image[23][23])} + {7'd0,(kernel[3][1] ~^ image[23][24])} + {7'd0,(kernel[3][2] ~^ image[23][25])} + {7'd0,(kernel[3][3] ~^ image[23][26])} + {7'd0,(kernel[3][4] ~^ image[23][27])} + {7'd0,(kernel[4][0] ~^ image[24][23])} + {7'd0,(kernel[4][1] ~^ image[24][24])} + {7'd0,(kernel[4][2] ~^ image[24][25])} + {7'd0,(kernel[4][3] ~^ image[24][26])} + {7'd0,(kernel[4][4] ~^ image[24][27])};
assign out_fmap[21][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[21][0])} + {7'd0,(kernel[0][1] ~^ image[21][1])} + {7'd0,(kernel[0][2] ~^ image[21][2])} + {7'd0,(kernel[0][3] ~^ image[21][3])} + {7'd0,(kernel[0][4] ~^ image[21][4])} + {7'd0,(kernel[1][0] ~^ image[22][0])} + {7'd0,(kernel[1][1] ~^ image[22][1])} + {7'd0,(kernel[1][2] ~^ image[22][2])} + {7'd0,(kernel[1][3] ~^ image[22][3])} + {7'd0,(kernel[1][4] ~^ image[22][4])} + {7'd0,(kernel[2][0] ~^ image[23][0])} + {7'd0,(kernel[2][1] ~^ image[23][1])} + {7'd0,(kernel[2][2] ~^ image[23][2])} + {7'd0,(kernel[2][3] ~^ image[23][3])} + {7'd0,(kernel[2][4] ~^ image[23][4])} + {7'd0,(kernel[3][0] ~^ image[24][0])} + {7'd0,(kernel[3][1] ~^ image[24][1])} + {7'd0,(kernel[3][2] ~^ image[24][2])} + {7'd0,(kernel[3][3] ~^ image[24][3])} + {7'd0,(kernel[3][4] ~^ image[24][4])} + {7'd0,(kernel[4][0] ~^ image[25][0])} + {7'd0,(kernel[4][1] ~^ image[25][1])} + {7'd0,(kernel[4][2] ~^ image[25][2])} + {7'd0,(kernel[4][3] ~^ image[25][3])} + {7'd0,(kernel[4][4] ~^ image[25][4])};
assign out_fmap[21][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[21][1])} + {7'd0,(kernel[0][1] ~^ image[21][2])} + {7'd0,(kernel[0][2] ~^ image[21][3])} + {7'd0,(kernel[0][3] ~^ image[21][4])} + {7'd0,(kernel[0][4] ~^ image[21][5])} + {7'd0,(kernel[1][0] ~^ image[22][1])} + {7'd0,(kernel[1][1] ~^ image[22][2])} + {7'd0,(kernel[1][2] ~^ image[22][3])} + {7'd0,(kernel[1][3] ~^ image[22][4])} + {7'd0,(kernel[1][4] ~^ image[22][5])} + {7'd0,(kernel[2][0] ~^ image[23][1])} + {7'd0,(kernel[2][1] ~^ image[23][2])} + {7'd0,(kernel[2][2] ~^ image[23][3])} + {7'd0,(kernel[2][3] ~^ image[23][4])} + {7'd0,(kernel[2][4] ~^ image[23][5])} + {7'd0,(kernel[3][0] ~^ image[24][1])} + {7'd0,(kernel[3][1] ~^ image[24][2])} + {7'd0,(kernel[3][2] ~^ image[24][3])} + {7'd0,(kernel[3][3] ~^ image[24][4])} + {7'd0,(kernel[3][4] ~^ image[24][5])} + {7'd0,(kernel[4][0] ~^ image[25][1])} + {7'd0,(kernel[4][1] ~^ image[25][2])} + {7'd0,(kernel[4][2] ~^ image[25][3])} + {7'd0,(kernel[4][3] ~^ image[25][4])} + {7'd0,(kernel[4][4] ~^ image[25][5])};
assign out_fmap[21][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[21][2])} + {7'd0,(kernel[0][1] ~^ image[21][3])} + {7'd0,(kernel[0][2] ~^ image[21][4])} + {7'd0,(kernel[0][3] ~^ image[21][5])} + {7'd0,(kernel[0][4] ~^ image[21][6])} + {7'd0,(kernel[1][0] ~^ image[22][2])} + {7'd0,(kernel[1][1] ~^ image[22][3])} + {7'd0,(kernel[1][2] ~^ image[22][4])} + {7'd0,(kernel[1][3] ~^ image[22][5])} + {7'd0,(kernel[1][4] ~^ image[22][6])} + {7'd0,(kernel[2][0] ~^ image[23][2])} + {7'd0,(kernel[2][1] ~^ image[23][3])} + {7'd0,(kernel[2][2] ~^ image[23][4])} + {7'd0,(kernel[2][3] ~^ image[23][5])} + {7'd0,(kernel[2][4] ~^ image[23][6])} + {7'd0,(kernel[3][0] ~^ image[24][2])} + {7'd0,(kernel[3][1] ~^ image[24][3])} + {7'd0,(kernel[3][2] ~^ image[24][4])} + {7'd0,(kernel[3][3] ~^ image[24][5])} + {7'd0,(kernel[3][4] ~^ image[24][6])} + {7'd0,(kernel[4][0] ~^ image[25][2])} + {7'd0,(kernel[4][1] ~^ image[25][3])} + {7'd0,(kernel[4][2] ~^ image[25][4])} + {7'd0,(kernel[4][3] ~^ image[25][5])} + {7'd0,(kernel[4][4] ~^ image[25][6])};
assign out_fmap[21][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[21][3])} + {7'd0,(kernel[0][1] ~^ image[21][4])} + {7'd0,(kernel[0][2] ~^ image[21][5])} + {7'd0,(kernel[0][3] ~^ image[21][6])} + {7'd0,(kernel[0][4] ~^ image[21][7])} + {7'd0,(kernel[1][0] ~^ image[22][3])} + {7'd0,(kernel[1][1] ~^ image[22][4])} + {7'd0,(kernel[1][2] ~^ image[22][5])} + {7'd0,(kernel[1][3] ~^ image[22][6])} + {7'd0,(kernel[1][4] ~^ image[22][7])} + {7'd0,(kernel[2][0] ~^ image[23][3])} + {7'd0,(kernel[2][1] ~^ image[23][4])} + {7'd0,(kernel[2][2] ~^ image[23][5])} + {7'd0,(kernel[2][3] ~^ image[23][6])} + {7'd0,(kernel[2][4] ~^ image[23][7])} + {7'd0,(kernel[3][0] ~^ image[24][3])} + {7'd0,(kernel[3][1] ~^ image[24][4])} + {7'd0,(kernel[3][2] ~^ image[24][5])} + {7'd0,(kernel[3][3] ~^ image[24][6])} + {7'd0,(kernel[3][4] ~^ image[24][7])} + {7'd0,(kernel[4][0] ~^ image[25][3])} + {7'd0,(kernel[4][1] ~^ image[25][4])} + {7'd0,(kernel[4][2] ~^ image[25][5])} + {7'd0,(kernel[4][3] ~^ image[25][6])} + {7'd0,(kernel[4][4] ~^ image[25][7])};
assign out_fmap[21][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[21][4])} + {7'd0,(kernel[0][1] ~^ image[21][5])} + {7'd0,(kernel[0][2] ~^ image[21][6])} + {7'd0,(kernel[0][3] ~^ image[21][7])} + {7'd0,(kernel[0][4] ~^ image[21][8])} + {7'd0,(kernel[1][0] ~^ image[22][4])} + {7'd0,(kernel[1][1] ~^ image[22][5])} + {7'd0,(kernel[1][2] ~^ image[22][6])} + {7'd0,(kernel[1][3] ~^ image[22][7])} + {7'd0,(kernel[1][4] ~^ image[22][8])} + {7'd0,(kernel[2][0] ~^ image[23][4])} + {7'd0,(kernel[2][1] ~^ image[23][5])} + {7'd0,(kernel[2][2] ~^ image[23][6])} + {7'd0,(kernel[2][3] ~^ image[23][7])} + {7'd0,(kernel[2][4] ~^ image[23][8])} + {7'd0,(kernel[3][0] ~^ image[24][4])} + {7'd0,(kernel[3][1] ~^ image[24][5])} + {7'd0,(kernel[3][2] ~^ image[24][6])} + {7'd0,(kernel[3][3] ~^ image[24][7])} + {7'd0,(kernel[3][4] ~^ image[24][8])} + {7'd0,(kernel[4][0] ~^ image[25][4])} + {7'd0,(kernel[4][1] ~^ image[25][5])} + {7'd0,(kernel[4][2] ~^ image[25][6])} + {7'd0,(kernel[4][3] ~^ image[25][7])} + {7'd0,(kernel[4][4] ~^ image[25][8])};
assign out_fmap[21][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[21][5])} + {7'd0,(kernel[0][1] ~^ image[21][6])} + {7'd0,(kernel[0][2] ~^ image[21][7])} + {7'd0,(kernel[0][3] ~^ image[21][8])} + {7'd0,(kernel[0][4] ~^ image[21][9])} + {7'd0,(kernel[1][0] ~^ image[22][5])} + {7'd0,(kernel[1][1] ~^ image[22][6])} + {7'd0,(kernel[1][2] ~^ image[22][7])} + {7'd0,(kernel[1][3] ~^ image[22][8])} + {7'd0,(kernel[1][4] ~^ image[22][9])} + {7'd0,(kernel[2][0] ~^ image[23][5])} + {7'd0,(kernel[2][1] ~^ image[23][6])} + {7'd0,(kernel[2][2] ~^ image[23][7])} + {7'd0,(kernel[2][3] ~^ image[23][8])} + {7'd0,(kernel[2][4] ~^ image[23][9])} + {7'd0,(kernel[3][0] ~^ image[24][5])} + {7'd0,(kernel[3][1] ~^ image[24][6])} + {7'd0,(kernel[3][2] ~^ image[24][7])} + {7'd0,(kernel[3][3] ~^ image[24][8])} + {7'd0,(kernel[3][4] ~^ image[24][9])} + {7'd0,(kernel[4][0] ~^ image[25][5])} + {7'd0,(kernel[4][1] ~^ image[25][6])} + {7'd0,(kernel[4][2] ~^ image[25][7])} + {7'd0,(kernel[4][3] ~^ image[25][8])} + {7'd0,(kernel[4][4] ~^ image[25][9])};
assign out_fmap[21][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[21][6])} + {7'd0,(kernel[0][1] ~^ image[21][7])} + {7'd0,(kernel[0][2] ~^ image[21][8])} + {7'd0,(kernel[0][3] ~^ image[21][9])} + {7'd0,(kernel[0][4] ~^ image[21][10])} + {7'd0,(kernel[1][0] ~^ image[22][6])} + {7'd0,(kernel[1][1] ~^ image[22][7])} + {7'd0,(kernel[1][2] ~^ image[22][8])} + {7'd0,(kernel[1][3] ~^ image[22][9])} + {7'd0,(kernel[1][4] ~^ image[22][10])} + {7'd0,(kernel[2][0] ~^ image[23][6])} + {7'd0,(kernel[2][1] ~^ image[23][7])} + {7'd0,(kernel[2][2] ~^ image[23][8])} + {7'd0,(kernel[2][3] ~^ image[23][9])} + {7'd0,(kernel[2][4] ~^ image[23][10])} + {7'd0,(kernel[3][0] ~^ image[24][6])} + {7'd0,(kernel[3][1] ~^ image[24][7])} + {7'd0,(kernel[3][2] ~^ image[24][8])} + {7'd0,(kernel[3][3] ~^ image[24][9])} + {7'd0,(kernel[3][4] ~^ image[24][10])} + {7'd0,(kernel[4][0] ~^ image[25][6])} + {7'd0,(kernel[4][1] ~^ image[25][7])} + {7'd0,(kernel[4][2] ~^ image[25][8])} + {7'd0,(kernel[4][3] ~^ image[25][9])} + {7'd0,(kernel[4][4] ~^ image[25][10])};
assign out_fmap[21][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[21][7])} + {7'd0,(kernel[0][1] ~^ image[21][8])} + {7'd0,(kernel[0][2] ~^ image[21][9])} + {7'd0,(kernel[0][3] ~^ image[21][10])} + {7'd0,(kernel[0][4] ~^ image[21][11])} + {7'd0,(kernel[1][0] ~^ image[22][7])} + {7'd0,(kernel[1][1] ~^ image[22][8])} + {7'd0,(kernel[1][2] ~^ image[22][9])} + {7'd0,(kernel[1][3] ~^ image[22][10])} + {7'd0,(kernel[1][4] ~^ image[22][11])} + {7'd0,(kernel[2][0] ~^ image[23][7])} + {7'd0,(kernel[2][1] ~^ image[23][8])} + {7'd0,(kernel[2][2] ~^ image[23][9])} + {7'd0,(kernel[2][3] ~^ image[23][10])} + {7'd0,(kernel[2][4] ~^ image[23][11])} + {7'd0,(kernel[3][0] ~^ image[24][7])} + {7'd0,(kernel[3][1] ~^ image[24][8])} + {7'd0,(kernel[3][2] ~^ image[24][9])} + {7'd0,(kernel[3][3] ~^ image[24][10])} + {7'd0,(kernel[3][4] ~^ image[24][11])} + {7'd0,(kernel[4][0] ~^ image[25][7])} + {7'd0,(kernel[4][1] ~^ image[25][8])} + {7'd0,(kernel[4][2] ~^ image[25][9])} + {7'd0,(kernel[4][3] ~^ image[25][10])} + {7'd0,(kernel[4][4] ~^ image[25][11])};
assign out_fmap[21][8][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[21][8])} + {7'd0,(kernel[0][1] ~^ image[21][9])} + {7'd0,(kernel[0][2] ~^ image[21][10])} + {7'd0,(kernel[0][3] ~^ image[21][11])} + {7'd0,(kernel[0][4] ~^ image[21][12])} + {7'd0,(kernel[1][0] ~^ image[22][8])} + {7'd0,(kernel[1][1] ~^ image[22][9])} + {7'd0,(kernel[1][2] ~^ image[22][10])} + {7'd0,(kernel[1][3] ~^ image[22][11])} + {7'd0,(kernel[1][4] ~^ image[22][12])} + {7'd0,(kernel[2][0] ~^ image[23][8])} + {7'd0,(kernel[2][1] ~^ image[23][9])} + {7'd0,(kernel[2][2] ~^ image[23][10])} + {7'd0,(kernel[2][3] ~^ image[23][11])} + {7'd0,(kernel[2][4] ~^ image[23][12])} + {7'd0,(kernel[3][0] ~^ image[24][8])} + {7'd0,(kernel[3][1] ~^ image[24][9])} + {7'd0,(kernel[3][2] ~^ image[24][10])} + {7'd0,(kernel[3][3] ~^ image[24][11])} + {7'd0,(kernel[3][4] ~^ image[24][12])} + {7'd0,(kernel[4][0] ~^ image[25][8])} + {7'd0,(kernel[4][1] ~^ image[25][9])} + {7'd0,(kernel[4][2] ~^ image[25][10])} + {7'd0,(kernel[4][3] ~^ image[25][11])} + {7'd0,(kernel[4][4] ~^ image[25][12])};
assign out_fmap[21][9][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[21][9])} + {7'd0,(kernel[0][1] ~^ image[21][10])} + {7'd0,(kernel[0][2] ~^ image[21][11])} + {7'd0,(kernel[0][3] ~^ image[21][12])} + {7'd0,(kernel[0][4] ~^ image[21][13])} + {7'd0,(kernel[1][0] ~^ image[22][9])} + {7'd0,(kernel[1][1] ~^ image[22][10])} + {7'd0,(kernel[1][2] ~^ image[22][11])} + {7'd0,(kernel[1][3] ~^ image[22][12])} + {7'd0,(kernel[1][4] ~^ image[22][13])} + {7'd0,(kernel[2][0] ~^ image[23][9])} + {7'd0,(kernel[2][1] ~^ image[23][10])} + {7'd0,(kernel[2][2] ~^ image[23][11])} + {7'd0,(kernel[2][3] ~^ image[23][12])} + {7'd0,(kernel[2][4] ~^ image[23][13])} + {7'd0,(kernel[3][0] ~^ image[24][9])} + {7'd0,(kernel[3][1] ~^ image[24][10])} + {7'd0,(kernel[3][2] ~^ image[24][11])} + {7'd0,(kernel[3][3] ~^ image[24][12])} + {7'd0,(kernel[3][4] ~^ image[24][13])} + {7'd0,(kernel[4][0] ~^ image[25][9])} + {7'd0,(kernel[4][1] ~^ image[25][10])} + {7'd0,(kernel[4][2] ~^ image[25][11])} + {7'd0,(kernel[4][3] ~^ image[25][12])} + {7'd0,(kernel[4][4] ~^ image[25][13])};
assign out_fmap[21][10][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[21][10])} + {7'd0,(kernel[0][1] ~^ image[21][11])} + {7'd0,(kernel[0][2] ~^ image[21][12])} + {7'd0,(kernel[0][3] ~^ image[21][13])} + {7'd0,(kernel[0][4] ~^ image[21][14])} + {7'd0,(kernel[1][0] ~^ image[22][10])} + {7'd0,(kernel[1][1] ~^ image[22][11])} + {7'd0,(kernel[1][2] ~^ image[22][12])} + {7'd0,(kernel[1][3] ~^ image[22][13])} + {7'd0,(kernel[1][4] ~^ image[22][14])} + {7'd0,(kernel[2][0] ~^ image[23][10])} + {7'd0,(kernel[2][1] ~^ image[23][11])} + {7'd0,(kernel[2][2] ~^ image[23][12])} + {7'd0,(kernel[2][3] ~^ image[23][13])} + {7'd0,(kernel[2][4] ~^ image[23][14])} + {7'd0,(kernel[3][0] ~^ image[24][10])} + {7'd0,(kernel[3][1] ~^ image[24][11])} + {7'd0,(kernel[3][2] ~^ image[24][12])} + {7'd0,(kernel[3][3] ~^ image[24][13])} + {7'd0,(kernel[3][4] ~^ image[24][14])} + {7'd0,(kernel[4][0] ~^ image[25][10])} + {7'd0,(kernel[4][1] ~^ image[25][11])} + {7'd0,(kernel[4][2] ~^ image[25][12])} + {7'd0,(kernel[4][3] ~^ image[25][13])} + {7'd0,(kernel[4][4] ~^ image[25][14])};
assign out_fmap[21][11][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[21][11])} + {7'd0,(kernel[0][1] ~^ image[21][12])} + {7'd0,(kernel[0][2] ~^ image[21][13])} + {7'd0,(kernel[0][3] ~^ image[21][14])} + {7'd0,(kernel[0][4] ~^ image[21][15])} + {7'd0,(kernel[1][0] ~^ image[22][11])} + {7'd0,(kernel[1][1] ~^ image[22][12])} + {7'd0,(kernel[1][2] ~^ image[22][13])} + {7'd0,(kernel[1][3] ~^ image[22][14])} + {7'd0,(kernel[1][4] ~^ image[22][15])} + {7'd0,(kernel[2][0] ~^ image[23][11])} + {7'd0,(kernel[2][1] ~^ image[23][12])} + {7'd0,(kernel[2][2] ~^ image[23][13])} + {7'd0,(kernel[2][3] ~^ image[23][14])} + {7'd0,(kernel[2][4] ~^ image[23][15])} + {7'd0,(kernel[3][0] ~^ image[24][11])} + {7'd0,(kernel[3][1] ~^ image[24][12])} + {7'd0,(kernel[3][2] ~^ image[24][13])} + {7'd0,(kernel[3][3] ~^ image[24][14])} + {7'd0,(kernel[3][4] ~^ image[24][15])} + {7'd0,(kernel[4][0] ~^ image[25][11])} + {7'd0,(kernel[4][1] ~^ image[25][12])} + {7'd0,(kernel[4][2] ~^ image[25][13])} + {7'd0,(kernel[4][3] ~^ image[25][14])} + {7'd0,(kernel[4][4] ~^ image[25][15])};
assign out_fmap[21][12][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[21][12])} + {7'd0,(kernel[0][1] ~^ image[21][13])} + {7'd0,(kernel[0][2] ~^ image[21][14])} + {7'd0,(kernel[0][3] ~^ image[21][15])} + {7'd0,(kernel[0][4] ~^ image[21][16])} + {7'd0,(kernel[1][0] ~^ image[22][12])} + {7'd0,(kernel[1][1] ~^ image[22][13])} + {7'd0,(kernel[1][2] ~^ image[22][14])} + {7'd0,(kernel[1][3] ~^ image[22][15])} + {7'd0,(kernel[1][4] ~^ image[22][16])} + {7'd0,(kernel[2][0] ~^ image[23][12])} + {7'd0,(kernel[2][1] ~^ image[23][13])} + {7'd0,(kernel[2][2] ~^ image[23][14])} + {7'd0,(kernel[2][3] ~^ image[23][15])} + {7'd0,(kernel[2][4] ~^ image[23][16])} + {7'd0,(kernel[3][0] ~^ image[24][12])} + {7'd0,(kernel[3][1] ~^ image[24][13])} + {7'd0,(kernel[3][2] ~^ image[24][14])} + {7'd0,(kernel[3][3] ~^ image[24][15])} + {7'd0,(kernel[3][4] ~^ image[24][16])} + {7'd0,(kernel[4][0] ~^ image[25][12])} + {7'd0,(kernel[4][1] ~^ image[25][13])} + {7'd0,(kernel[4][2] ~^ image[25][14])} + {7'd0,(kernel[4][3] ~^ image[25][15])} + {7'd0,(kernel[4][4] ~^ image[25][16])};
assign out_fmap[21][13][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[21][13])} + {7'd0,(kernel[0][1] ~^ image[21][14])} + {7'd0,(kernel[0][2] ~^ image[21][15])} + {7'd0,(kernel[0][3] ~^ image[21][16])} + {7'd0,(kernel[0][4] ~^ image[21][17])} + {7'd0,(kernel[1][0] ~^ image[22][13])} + {7'd0,(kernel[1][1] ~^ image[22][14])} + {7'd0,(kernel[1][2] ~^ image[22][15])} + {7'd0,(kernel[1][3] ~^ image[22][16])} + {7'd0,(kernel[1][4] ~^ image[22][17])} + {7'd0,(kernel[2][0] ~^ image[23][13])} + {7'd0,(kernel[2][1] ~^ image[23][14])} + {7'd0,(kernel[2][2] ~^ image[23][15])} + {7'd0,(kernel[2][3] ~^ image[23][16])} + {7'd0,(kernel[2][4] ~^ image[23][17])} + {7'd0,(kernel[3][0] ~^ image[24][13])} + {7'd0,(kernel[3][1] ~^ image[24][14])} + {7'd0,(kernel[3][2] ~^ image[24][15])} + {7'd0,(kernel[3][3] ~^ image[24][16])} + {7'd0,(kernel[3][4] ~^ image[24][17])} + {7'd0,(kernel[4][0] ~^ image[25][13])} + {7'd0,(kernel[4][1] ~^ image[25][14])} + {7'd0,(kernel[4][2] ~^ image[25][15])} + {7'd0,(kernel[4][3] ~^ image[25][16])} + {7'd0,(kernel[4][4] ~^ image[25][17])};
assign out_fmap[21][14][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[21][14])} + {7'd0,(kernel[0][1] ~^ image[21][15])} + {7'd0,(kernel[0][2] ~^ image[21][16])} + {7'd0,(kernel[0][3] ~^ image[21][17])} + {7'd0,(kernel[0][4] ~^ image[21][18])} + {7'd0,(kernel[1][0] ~^ image[22][14])} + {7'd0,(kernel[1][1] ~^ image[22][15])} + {7'd0,(kernel[1][2] ~^ image[22][16])} + {7'd0,(kernel[1][3] ~^ image[22][17])} + {7'd0,(kernel[1][4] ~^ image[22][18])} + {7'd0,(kernel[2][0] ~^ image[23][14])} + {7'd0,(kernel[2][1] ~^ image[23][15])} + {7'd0,(kernel[2][2] ~^ image[23][16])} + {7'd0,(kernel[2][3] ~^ image[23][17])} + {7'd0,(kernel[2][4] ~^ image[23][18])} + {7'd0,(kernel[3][0] ~^ image[24][14])} + {7'd0,(kernel[3][1] ~^ image[24][15])} + {7'd0,(kernel[3][2] ~^ image[24][16])} + {7'd0,(kernel[3][3] ~^ image[24][17])} + {7'd0,(kernel[3][4] ~^ image[24][18])} + {7'd0,(kernel[4][0] ~^ image[25][14])} + {7'd0,(kernel[4][1] ~^ image[25][15])} + {7'd0,(kernel[4][2] ~^ image[25][16])} + {7'd0,(kernel[4][3] ~^ image[25][17])} + {7'd0,(kernel[4][4] ~^ image[25][18])};
assign out_fmap[21][15][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[21][15])} + {7'd0,(kernel[0][1] ~^ image[21][16])} + {7'd0,(kernel[0][2] ~^ image[21][17])} + {7'd0,(kernel[0][3] ~^ image[21][18])} + {7'd0,(kernel[0][4] ~^ image[21][19])} + {7'd0,(kernel[1][0] ~^ image[22][15])} + {7'd0,(kernel[1][1] ~^ image[22][16])} + {7'd0,(kernel[1][2] ~^ image[22][17])} + {7'd0,(kernel[1][3] ~^ image[22][18])} + {7'd0,(kernel[1][4] ~^ image[22][19])} + {7'd0,(kernel[2][0] ~^ image[23][15])} + {7'd0,(kernel[2][1] ~^ image[23][16])} + {7'd0,(kernel[2][2] ~^ image[23][17])} + {7'd0,(kernel[2][3] ~^ image[23][18])} + {7'd0,(kernel[2][4] ~^ image[23][19])} + {7'd0,(kernel[3][0] ~^ image[24][15])} + {7'd0,(kernel[3][1] ~^ image[24][16])} + {7'd0,(kernel[3][2] ~^ image[24][17])} + {7'd0,(kernel[3][3] ~^ image[24][18])} + {7'd0,(kernel[3][4] ~^ image[24][19])} + {7'd0,(kernel[4][0] ~^ image[25][15])} + {7'd0,(kernel[4][1] ~^ image[25][16])} + {7'd0,(kernel[4][2] ~^ image[25][17])} + {7'd0,(kernel[4][3] ~^ image[25][18])} + {7'd0,(kernel[4][4] ~^ image[25][19])};
assign out_fmap[21][16][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[21][16])} + {7'd0,(kernel[0][1] ~^ image[21][17])} + {7'd0,(kernel[0][2] ~^ image[21][18])} + {7'd0,(kernel[0][3] ~^ image[21][19])} + {7'd0,(kernel[0][4] ~^ image[21][20])} + {7'd0,(kernel[1][0] ~^ image[22][16])} + {7'd0,(kernel[1][1] ~^ image[22][17])} + {7'd0,(kernel[1][2] ~^ image[22][18])} + {7'd0,(kernel[1][3] ~^ image[22][19])} + {7'd0,(kernel[1][4] ~^ image[22][20])} + {7'd0,(kernel[2][0] ~^ image[23][16])} + {7'd0,(kernel[2][1] ~^ image[23][17])} + {7'd0,(kernel[2][2] ~^ image[23][18])} + {7'd0,(kernel[2][3] ~^ image[23][19])} + {7'd0,(kernel[2][4] ~^ image[23][20])} + {7'd0,(kernel[3][0] ~^ image[24][16])} + {7'd0,(kernel[3][1] ~^ image[24][17])} + {7'd0,(kernel[3][2] ~^ image[24][18])} + {7'd0,(kernel[3][3] ~^ image[24][19])} + {7'd0,(kernel[3][4] ~^ image[24][20])} + {7'd0,(kernel[4][0] ~^ image[25][16])} + {7'd0,(kernel[4][1] ~^ image[25][17])} + {7'd0,(kernel[4][2] ~^ image[25][18])} + {7'd0,(kernel[4][3] ~^ image[25][19])} + {7'd0,(kernel[4][4] ~^ image[25][20])};
assign out_fmap[21][17][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[21][17])} + {7'd0,(kernel[0][1] ~^ image[21][18])} + {7'd0,(kernel[0][2] ~^ image[21][19])} + {7'd0,(kernel[0][3] ~^ image[21][20])} + {7'd0,(kernel[0][4] ~^ image[21][21])} + {7'd0,(kernel[1][0] ~^ image[22][17])} + {7'd0,(kernel[1][1] ~^ image[22][18])} + {7'd0,(kernel[1][2] ~^ image[22][19])} + {7'd0,(kernel[1][3] ~^ image[22][20])} + {7'd0,(kernel[1][4] ~^ image[22][21])} + {7'd0,(kernel[2][0] ~^ image[23][17])} + {7'd0,(kernel[2][1] ~^ image[23][18])} + {7'd0,(kernel[2][2] ~^ image[23][19])} + {7'd0,(kernel[2][3] ~^ image[23][20])} + {7'd0,(kernel[2][4] ~^ image[23][21])} + {7'd0,(kernel[3][0] ~^ image[24][17])} + {7'd0,(kernel[3][1] ~^ image[24][18])} + {7'd0,(kernel[3][2] ~^ image[24][19])} + {7'd0,(kernel[3][3] ~^ image[24][20])} + {7'd0,(kernel[3][4] ~^ image[24][21])} + {7'd0,(kernel[4][0] ~^ image[25][17])} + {7'd0,(kernel[4][1] ~^ image[25][18])} + {7'd0,(kernel[4][2] ~^ image[25][19])} + {7'd0,(kernel[4][3] ~^ image[25][20])} + {7'd0,(kernel[4][4] ~^ image[25][21])};
assign out_fmap[21][18][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[21][18])} + {7'd0,(kernel[0][1] ~^ image[21][19])} + {7'd0,(kernel[0][2] ~^ image[21][20])} + {7'd0,(kernel[0][3] ~^ image[21][21])} + {7'd0,(kernel[0][4] ~^ image[21][22])} + {7'd0,(kernel[1][0] ~^ image[22][18])} + {7'd0,(kernel[1][1] ~^ image[22][19])} + {7'd0,(kernel[1][2] ~^ image[22][20])} + {7'd0,(kernel[1][3] ~^ image[22][21])} + {7'd0,(kernel[1][4] ~^ image[22][22])} + {7'd0,(kernel[2][0] ~^ image[23][18])} + {7'd0,(kernel[2][1] ~^ image[23][19])} + {7'd0,(kernel[2][2] ~^ image[23][20])} + {7'd0,(kernel[2][3] ~^ image[23][21])} + {7'd0,(kernel[2][4] ~^ image[23][22])} + {7'd0,(kernel[3][0] ~^ image[24][18])} + {7'd0,(kernel[3][1] ~^ image[24][19])} + {7'd0,(kernel[3][2] ~^ image[24][20])} + {7'd0,(kernel[3][3] ~^ image[24][21])} + {7'd0,(kernel[3][4] ~^ image[24][22])} + {7'd0,(kernel[4][0] ~^ image[25][18])} + {7'd0,(kernel[4][1] ~^ image[25][19])} + {7'd0,(kernel[4][2] ~^ image[25][20])} + {7'd0,(kernel[4][3] ~^ image[25][21])} + {7'd0,(kernel[4][4] ~^ image[25][22])};
assign out_fmap[21][19][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[21][19])} + {7'd0,(kernel[0][1] ~^ image[21][20])} + {7'd0,(kernel[0][2] ~^ image[21][21])} + {7'd0,(kernel[0][3] ~^ image[21][22])} + {7'd0,(kernel[0][4] ~^ image[21][23])} + {7'd0,(kernel[1][0] ~^ image[22][19])} + {7'd0,(kernel[1][1] ~^ image[22][20])} + {7'd0,(kernel[1][2] ~^ image[22][21])} + {7'd0,(kernel[1][3] ~^ image[22][22])} + {7'd0,(kernel[1][4] ~^ image[22][23])} + {7'd0,(kernel[2][0] ~^ image[23][19])} + {7'd0,(kernel[2][1] ~^ image[23][20])} + {7'd0,(kernel[2][2] ~^ image[23][21])} + {7'd0,(kernel[2][3] ~^ image[23][22])} + {7'd0,(kernel[2][4] ~^ image[23][23])} + {7'd0,(kernel[3][0] ~^ image[24][19])} + {7'd0,(kernel[3][1] ~^ image[24][20])} + {7'd0,(kernel[3][2] ~^ image[24][21])} + {7'd0,(kernel[3][3] ~^ image[24][22])} + {7'd0,(kernel[3][4] ~^ image[24][23])} + {7'd0,(kernel[4][0] ~^ image[25][19])} + {7'd0,(kernel[4][1] ~^ image[25][20])} + {7'd0,(kernel[4][2] ~^ image[25][21])} + {7'd0,(kernel[4][3] ~^ image[25][22])} + {7'd0,(kernel[4][4] ~^ image[25][23])};
assign out_fmap[21][20][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[21][20])} + {7'd0,(kernel[0][1] ~^ image[21][21])} + {7'd0,(kernel[0][2] ~^ image[21][22])} + {7'd0,(kernel[0][3] ~^ image[21][23])} + {7'd0,(kernel[0][4] ~^ image[21][24])} + {7'd0,(kernel[1][0] ~^ image[22][20])} + {7'd0,(kernel[1][1] ~^ image[22][21])} + {7'd0,(kernel[1][2] ~^ image[22][22])} + {7'd0,(kernel[1][3] ~^ image[22][23])} + {7'd0,(kernel[1][4] ~^ image[22][24])} + {7'd0,(kernel[2][0] ~^ image[23][20])} + {7'd0,(kernel[2][1] ~^ image[23][21])} + {7'd0,(kernel[2][2] ~^ image[23][22])} + {7'd0,(kernel[2][3] ~^ image[23][23])} + {7'd0,(kernel[2][4] ~^ image[23][24])} + {7'd0,(kernel[3][0] ~^ image[24][20])} + {7'd0,(kernel[3][1] ~^ image[24][21])} + {7'd0,(kernel[3][2] ~^ image[24][22])} + {7'd0,(kernel[3][3] ~^ image[24][23])} + {7'd0,(kernel[3][4] ~^ image[24][24])} + {7'd0,(kernel[4][0] ~^ image[25][20])} + {7'd0,(kernel[4][1] ~^ image[25][21])} + {7'd0,(kernel[4][2] ~^ image[25][22])} + {7'd0,(kernel[4][3] ~^ image[25][23])} + {7'd0,(kernel[4][4] ~^ image[25][24])};
assign out_fmap[21][21][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[21][21])} + {7'd0,(kernel[0][1] ~^ image[21][22])} + {7'd0,(kernel[0][2] ~^ image[21][23])} + {7'd0,(kernel[0][3] ~^ image[21][24])} + {7'd0,(kernel[0][4] ~^ image[21][25])} + {7'd0,(kernel[1][0] ~^ image[22][21])} + {7'd0,(kernel[1][1] ~^ image[22][22])} + {7'd0,(kernel[1][2] ~^ image[22][23])} + {7'd0,(kernel[1][3] ~^ image[22][24])} + {7'd0,(kernel[1][4] ~^ image[22][25])} + {7'd0,(kernel[2][0] ~^ image[23][21])} + {7'd0,(kernel[2][1] ~^ image[23][22])} + {7'd0,(kernel[2][2] ~^ image[23][23])} + {7'd0,(kernel[2][3] ~^ image[23][24])} + {7'd0,(kernel[2][4] ~^ image[23][25])} + {7'd0,(kernel[3][0] ~^ image[24][21])} + {7'd0,(kernel[3][1] ~^ image[24][22])} + {7'd0,(kernel[3][2] ~^ image[24][23])} + {7'd0,(kernel[3][3] ~^ image[24][24])} + {7'd0,(kernel[3][4] ~^ image[24][25])} + {7'd0,(kernel[4][0] ~^ image[25][21])} + {7'd0,(kernel[4][1] ~^ image[25][22])} + {7'd0,(kernel[4][2] ~^ image[25][23])} + {7'd0,(kernel[4][3] ~^ image[25][24])} + {7'd0,(kernel[4][4] ~^ image[25][25])};
assign out_fmap[21][22][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[21][22])} + {7'd0,(kernel[0][1] ~^ image[21][23])} + {7'd0,(kernel[0][2] ~^ image[21][24])} + {7'd0,(kernel[0][3] ~^ image[21][25])} + {7'd0,(kernel[0][4] ~^ image[21][26])} + {7'd0,(kernel[1][0] ~^ image[22][22])} + {7'd0,(kernel[1][1] ~^ image[22][23])} + {7'd0,(kernel[1][2] ~^ image[22][24])} + {7'd0,(kernel[1][3] ~^ image[22][25])} + {7'd0,(kernel[1][4] ~^ image[22][26])} + {7'd0,(kernel[2][0] ~^ image[23][22])} + {7'd0,(kernel[2][1] ~^ image[23][23])} + {7'd0,(kernel[2][2] ~^ image[23][24])} + {7'd0,(kernel[2][3] ~^ image[23][25])} + {7'd0,(kernel[2][4] ~^ image[23][26])} + {7'd0,(kernel[3][0] ~^ image[24][22])} + {7'd0,(kernel[3][1] ~^ image[24][23])} + {7'd0,(kernel[3][2] ~^ image[24][24])} + {7'd0,(kernel[3][3] ~^ image[24][25])} + {7'd0,(kernel[3][4] ~^ image[24][26])} + {7'd0,(kernel[4][0] ~^ image[25][22])} + {7'd0,(kernel[4][1] ~^ image[25][23])} + {7'd0,(kernel[4][2] ~^ image[25][24])} + {7'd0,(kernel[4][3] ~^ image[25][25])} + {7'd0,(kernel[4][4] ~^ image[25][26])};
assign out_fmap[21][23][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[21][23])} + {7'd0,(kernel[0][1] ~^ image[21][24])} + {7'd0,(kernel[0][2] ~^ image[21][25])} + {7'd0,(kernel[0][3] ~^ image[21][26])} + {7'd0,(kernel[0][4] ~^ image[21][27])} + {7'd0,(kernel[1][0] ~^ image[22][23])} + {7'd0,(kernel[1][1] ~^ image[22][24])} + {7'd0,(kernel[1][2] ~^ image[22][25])} + {7'd0,(kernel[1][3] ~^ image[22][26])} + {7'd0,(kernel[1][4] ~^ image[22][27])} + {7'd0,(kernel[2][0] ~^ image[23][23])} + {7'd0,(kernel[2][1] ~^ image[23][24])} + {7'd0,(kernel[2][2] ~^ image[23][25])} + {7'd0,(kernel[2][3] ~^ image[23][26])} + {7'd0,(kernel[2][4] ~^ image[23][27])} + {7'd0,(kernel[3][0] ~^ image[24][23])} + {7'd0,(kernel[3][1] ~^ image[24][24])} + {7'd0,(kernel[3][2] ~^ image[24][25])} + {7'd0,(kernel[3][3] ~^ image[24][26])} + {7'd0,(kernel[3][4] ~^ image[24][27])} + {7'd0,(kernel[4][0] ~^ image[25][23])} + {7'd0,(kernel[4][1] ~^ image[25][24])} + {7'd0,(kernel[4][2] ~^ image[25][25])} + {7'd0,(kernel[4][3] ~^ image[25][26])} + {7'd0,(kernel[4][4] ~^ image[25][27])};
assign out_fmap[22][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[22][0])} + {7'd0,(kernel[0][1] ~^ image[22][1])} + {7'd0,(kernel[0][2] ~^ image[22][2])} + {7'd0,(kernel[0][3] ~^ image[22][3])} + {7'd0,(kernel[0][4] ~^ image[22][4])} + {7'd0,(kernel[1][0] ~^ image[23][0])} + {7'd0,(kernel[1][1] ~^ image[23][1])} + {7'd0,(kernel[1][2] ~^ image[23][2])} + {7'd0,(kernel[1][3] ~^ image[23][3])} + {7'd0,(kernel[1][4] ~^ image[23][4])} + {7'd0,(kernel[2][0] ~^ image[24][0])} + {7'd0,(kernel[2][1] ~^ image[24][1])} + {7'd0,(kernel[2][2] ~^ image[24][2])} + {7'd0,(kernel[2][3] ~^ image[24][3])} + {7'd0,(kernel[2][4] ~^ image[24][4])} + {7'd0,(kernel[3][0] ~^ image[25][0])} + {7'd0,(kernel[3][1] ~^ image[25][1])} + {7'd0,(kernel[3][2] ~^ image[25][2])} + {7'd0,(kernel[3][3] ~^ image[25][3])} + {7'd0,(kernel[3][4] ~^ image[25][4])} + {7'd0,(kernel[4][0] ~^ image[26][0])} + {7'd0,(kernel[4][1] ~^ image[26][1])} + {7'd0,(kernel[4][2] ~^ image[26][2])} + {7'd0,(kernel[4][3] ~^ image[26][3])} + {7'd0,(kernel[4][4] ~^ image[26][4])};
assign out_fmap[22][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[22][1])} + {7'd0,(kernel[0][1] ~^ image[22][2])} + {7'd0,(kernel[0][2] ~^ image[22][3])} + {7'd0,(kernel[0][3] ~^ image[22][4])} + {7'd0,(kernel[0][4] ~^ image[22][5])} + {7'd0,(kernel[1][0] ~^ image[23][1])} + {7'd0,(kernel[1][1] ~^ image[23][2])} + {7'd0,(kernel[1][2] ~^ image[23][3])} + {7'd0,(kernel[1][3] ~^ image[23][4])} + {7'd0,(kernel[1][4] ~^ image[23][5])} + {7'd0,(kernel[2][0] ~^ image[24][1])} + {7'd0,(kernel[2][1] ~^ image[24][2])} + {7'd0,(kernel[2][2] ~^ image[24][3])} + {7'd0,(kernel[2][3] ~^ image[24][4])} + {7'd0,(kernel[2][4] ~^ image[24][5])} + {7'd0,(kernel[3][0] ~^ image[25][1])} + {7'd0,(kernel[3][1] ~^ image[25][2])} + {7'd0,(kernel[3][2] ~^ image[25][3])} + {7'd0,(kernel[3][3] ~^ image[25][4])} + {7'd0,(kernel[3][4] ~^ image[25][5])} + {7'd0,(kernel[4][0] ~^ image[26][1])} + {7'd0,(kernel[4][1] ~^ image[26][2])} + {7'd0,(kernel[4][2] ~^ image[26][3])} + {7'd0,(kernel[4][3] ~^ image[26][4])} + {7'd0,(kernel[4][4] ~^ image[26][5])};
assign out_fmap[22][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[22][2])} + {7'd0,(kernel[0][1] ~^ image[22][3])} + {7'd0,(kernel[0][2] ~^ image[22][4])} + {7'd0,(kernel[0][3] ~^ image[22][5])} + {7'd0,(kernel[0][4] ~^ image[22][6])} + {7'd0,(kernel[1][0] ~^ image[23][2])} + {7'd0,(kernel[1][1] ~^ image[23][3])} + {7'd0,(kernel[1][2] ~^ image[23][4])} + {7'd0,(kernel[1][3] ~^ image[23][5])} + {7'd0,(kernel[1][4] ~^ image[23][6])} + {7'd0,(kernel[2][0] ~^ image[24][2])} + {7'd0,(kernel[2][1] ~^ image[24][3])} + {7'd0,(kernel[2][2] ~^ image[24][4])} + {7'd0,(kernel[2][3] ~^ image[24][5])} + {7'd0,(kernel[2][4] ~^ image[24][6])} + {7'd0,(kernel[3][0] ~^ image[25][2])} + {7'd0,(kernel[3][1] ~^ image[25][3])} + {7'd0,(kernel[3][2] ~^ image[25][4])} + {7'd0,(kernel[3][3] ~^ image[25][5])} + {7'd0,(kernel[3][4] ~^ image[25][6])} + {7'd0,(kernel[4][0] ~^ image[26][2])} + {7'd0,(kernel[4][1] ~^ image[26][3])} + {7'd0,(kernel[4][2] ~^ image[26][4])} + {7'd0,(kernel[4][3] ~^ image[26][5])} + {7'd0,(kernel[4][4] ~^ image[26][6])};
assign out_fmap[22][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[22][3])} + {7'd0,(kernel[0][1] ~^ image[22][4])} + {7'd0,(kernel[0][2] ~^ image[22][5])} + {7'd0,(kernel[0][3] ~^ image[22][6])} + {7'd0,(kernel[0][4] ~^ image[22][7])} + {7'd0,(kernel[1][0] ~^ image[23][3])} + {7'd0,(kernel[1][1] ~^ image[23][4])} + {7'd0,(kernel[1][2] ~^ image[23][5])} + {7'd0,(kernel[1][3] ~^ image[23][6])} + {7'd0,(kernel[1][4] ~^ image[23][7])} + {7'd0,(kernel[2][0] ~^ image[24][3])} + {7'd0,(kernel[2][1] ~^ image[24][4])} + {7'd0,(kernel[2][2] ~^ image[24][5])} + {7'd0,(kernel[2][3] ~^ image[24][6])} + {7'd0,(kernel[2][4] ~^ image[24][7])} + {7'd0,(kernel[3][0] ~^ image[25][3])} + {7'd0,(kernel[3][1] ~^ image[25][4])} + {7'd0,(kernel[3][2] ~^ image[25][5])} + {7'd0,(kernel[3][3] ~^ image[25][6])} + {7'd0,(kernel[3][4] ~^ image[25][7])} + {7'd0,(kernel[4][0] ~^ image[26][3])} + {7'd0,(kernel[4][1] ~^ image[26][4])} + {7'd0,(kernel[4][2] ~^ image[26][5])} + {7'd0,(kernel[4][3] ~^ image[26][6])} + {7'd0,(kernel[4][4] ~^ image[26][7])};
assign out_fmap[22][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[22][4])} + {7'd0,(kernel[0][1] ~^ image[22][5])} + {7'd0,(kernel[0][2] ~^ image[22][6])} + {7'd0,(kernel[0][3] ~^ image[22][7])} + {7'd0,(kernel[0][4] ~^ image[22][8])} + {7'd0,(kernel[1][0] ~^ image[23][4])} + {7'd0,(kernel[1][1] ~^ image[23][5])} + {7'd0,(kernel[1][2] ~^ image[23][6])} + {7'd0,(kernel[1][3] ~^ image[23][7])} + {7'd0,(kernel[1][4] ~^ image[23][8])} + {7'd0,(kernel[2][0] ~^ image[24][4])} + {7'd0,(kernel[2][1] ~^ image[24][5])} + {7'd0,(kernel[2][2] ~^ image[24][6])} + {7'd0,(kernel[2][3] ~^ image[24][7])} + {7'd0,(kernel[2][4] ~^ image[24][8])} + {7'd0,(kernel[3][0] ~^ image[25][4])} + {7'd0,(kernel[3][1] ~^ image[25][5])} + {7'd0,(kernel[3][2] ~^ image[25][6])} + {7'd0,(kernel[3][3] ~^ image[25][7])} + {7'd0,(kernel[3][4] ~^ image[25][8])} + {7'd0,(kernel[4][0] ~^ image[26][4])} + {7'd0,(kernel[4][1] ~^ image[26][5])} + {7'd0,(kernel[4][2] ~^ image[26][6])} + {7'd0,(kernel[4][3] ~^ image[26][7])} + {7'd0,(kernel[4][4] ~^ image[26][8])};
assign out_fmap[22][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[22][5])} + {7'd0,(kernel[0][1] ~^ image[22][6])} + {7'd0,(kernel[0][2] ~^ image[22][7])} + {7'd0,(kernel[0][3] ~^ image[22][8])} + {7'd0,(kernel[0][4] ~^ image[22][9])} + {7'd0,(kernel[1][0] ~^ image[23][5])} + {7'd0,(kernel[1][1] ~^ image[23][6])} + {7'd0,(kernel[1][2] ~^ image[23][7])} + {7'd0,(kernel[1][3] ~^ image[23][8])} + {7'd0,(kernel[1][4] ~^ image[23][9])} + {7'd0,(kernel[2][0] ~^ image[24][5])} + {7'd0,(kernel[2][1] ~^ image[24][6])} + {7'd0,(kernel[2][2] ~^ image[24][7])} + {7'd0,(kernel[2][3] ~^ image[24][8])} + {7'd0,(kernel[2][4] ~^ image[24][9])} + {7'd0,(kernel[3][0] ~^ image[25][5])} + {7'd0,(kernel[3][1] ~^ image[25][6])} + {7'd0,(kernel[3][2] ~^ image[25][7])} + {7'd0,(kernel[3][3] ~^ image[25][8])} + {7'd0,(kernel[3][4] ~^ image[25][9])} + {7'd0,(kernel[4][0] ~^ image[26][5])} + {7'd0,(kernel[4][1] ~^ image[26][6])} + {7'd0,(kernel[4][2] ~^ image[26][7])} + {7'd0,(kernel[4][3] ~^ image[26][8])} + {7'd0,(kernel[4][4] ~^ image[26][9])};
assign out_fmap[22][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[22][6])} + {7'd0,(kernel[0][1] ~^ image[22][7])} + {7'd0,(kernel[0][2] ~^ image[22][8])} + {7'd0,(kernel[0][3] ~^ image[22][9])} + {7'd0,(kernel[0][4] ~^ image[22][10])} + {7'd0,(kernel[1][0] ~^ image[23][6])} + {7'd0,(kernel[1][1] ~^ image[23][7])} + {7'd0,(kernel[1][2] ~^ image[23][8])} + {7'd0,(kernel[1][3] ~^ image[23][9])} + {7'd0,(kernel[1][4] ~^ image[23][10])} + {7'd0,(kernel[2][0] ~^ image[24][6])} + {7'd0,(kernel[2][1] ~^ image[24][7])} + {7'd0,(kernel[2][2] ~^ image[24][8])} + {7'd0,(kernel[2][3] ~^ image[24][9])} + {7'd0,(kernel[2][4] ~^ image[24][10])} + {7'd0,(kernel[3][0] ~^ image[25][6])} + {7'd0,(kernel[3][1] ~^ image[25][7])} + {7'd0,(kernel[3][2] ~^ image[25][8])} + {7'd0,(kernel[3][3] ~^ image[25][9])} + {7'd0,(kernel[3][4] ~^ image[25][10])} + {7'd0,(kernel[4][0] ~^ image[26][6])} + {7'd0,(kernel[4][1] ~^ image[26][7])} + {7'd0,(kernel[4][2] ~^ image[26][8])} + {7'd0,(kernel[4][3] ~^ image[26][9])} + {7'd0,(kernel[4][4] ~^ image[26][10])};
assign out_fmap[22][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[22][7])} + {7'd0,(kernel[0][1] ~^ image[22][8])} + {7'd0,(kernel[0][2] ~^ image[22][9])} + {7'd0,(kernel[0][3] ~^ image[22][10])} + {7'd0,(kernel[0][4] ~^ image[22][11])} + {7'd0,(kernel[1][0] ~^ image[23][7])} + {7'd0,(kernel[1][1] ~^ image[23][8])} + {7'd0,(kernel[1][2] ~^ image[23][9])} + {7'd0,(kernel[1][3] ~^ image[23][10])} + {7'd0,(kernel[1][4] ~^ image[23][11])} + {7'd0,(kernel[2][0] ~^ image[24][7])} + {7'd0,(kernel[2][1] ~^ image[24][8])} + {7'd0,(kernel[2][2] ~^ image[24][9])} + {7'd0,(kernel[2][3] ~^ image[24][10])} + {7'd0,(kernel[2][4] ~^ image[24][11])} + {7'd0,(kernel[3][0] ~^ image[25][7])} + {7'd0,(kernel[3][1] ~^ image[25][8])} + {7'd0,(kernel[3][2] ~^ image[25][9])} + {7'd0,(kernel[3][3] ~^ image[25][10])} + {7'd0,(kernel[3][4] ~^ image[25][11])} + {7'd0,(kernel[4][0] ~^ image[26][7])} + {7'd0,(kernel[4][1] ~^ image[26][8])} + {7'd0,(kernel[4][2] ~^ image[26][9])} + {7'd0,(kernel[4][3] ~^ image[26][10])} + {7'd0,(kernel[4][4] ~^ image[26][11])};
assign out_fmap[22][8][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[22][8])} + {7'd0,(kernel[0][1] ~^ image[22][9])} + {7'd0,(kernel[0][2] ~^ image[22][10])} + {7'd0,(kernel[0][3] ~^ image[22][11])} + {7'd0,(kernel[0][4] ~^ image[22][12])} + {7'd0,(kernel[1][0] ~^ image[23][8])} + {7'd0,(kernel[1][1] ~^ image[23][9])} + {7'd0,(kernel[1][2] ~^ image[23][10])} + {7'd0,(kernel[1][3] ~^ image[23][11])} + {7'd0,(kernel[1][4] ~^ image[23][12])} + {7'd0,(kernel[2][0] ~^ image[24][8])} + {7'd0,(kernel[2][1] ~^ image[24][9])} + {7'd0,(kernel[2][2] ~^ image[24][10])} + {7'd0,(kernel[2][3] ~^ image[24][11])} + {7'd0,(kernel[2][4] ~^ image[24][12])} + {7'd0,(kernel[3][0] ~^ image[25][8])} + {7'd0,(kernel[3][1] ~^ image[25][9])} + {7'd0,(kernel[3][2] ~^ image[25][10])} + {7'd0,(kernel[3][3] ~^ image[25][11])} + {7'd0,(kernel[3][4] ~^ image[25][12])} + {7'd0,(kernel[4][0] ~^ image[26][8])} + {7'd0,(kernel[4][1] ~^ image[26][9])} + {7'd0,(kernel[4][2] ~^ image[26][10])} + {7'd0,(kernel[4][3] ~^ image[26][11])} + {7'd0,(kernel[4][4] ~^ image[26][12])};
assign out_fmap[22][9][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[22][9])} + {7'd0,(kernel[0][1] ~^ image[22][10])} + {7'd0,(kernel[0][2] ~^ image[22][11])} + {7'd0,(kernel[0][3] ~^ image[22][12])} + {7'd0,(kernel[0][4] ~^ image[22][13])} + {7'd0,(kernel[1][0] ~^ image[23][9])} + {7'd0,(kernel[1][1] ~^ image[23][10])} + {7'd0,(kernel[1][2] ~^ image[23][11])} + {7'd0,(kernel[1][3] ~^ image[23][12])} + {7'd0,(kernel[1][4] ~^ image[23][13])} + {7'd0,(kernel[2][0] ~^ image[24][9])} + {7'd0,(kernel[2][1] ~^ image[24][10])} + {7'd0,(kernel[2][2] ~^ image[24][11])} + {7'd0,(kernel[2][3] ~^ image[24][12])} + {7'd0,(kernel[2][4] ~^ image[24][13])} + {7'd0,(kernel[3][0] ~^ image[25][9])} + {7'd0,(kernel[3][1] ~^ image[25][10])} + {7'd0,(kernel[3][2] ~^ image[25][11])} + {7'd0,(kernel[3][3] ~^ image[25][12])} + {7'd0,(kernel[3][4] ~^ image[25][13])} + {7'd0,(kernel[4][0] ~^ image[26][9])} + {7'd0,(kernel[4][1] ~^ image[26][10])} + {7'd0,(kernel[4][2] ~^ image[26][11])} + {7'd0,(kernel[4][3] ~^ image[26][12])} + {7'd0,(kernel[4][4] ~^ image[26][13])};
assign out_fmap[22][10][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[22][10])} + {7'd0,(kernel[0][1] ~^ image[22][11])} + {7'd0,(kernel[0][2] ~^ image[22][12])} + {7'd0,(kernel[0][3] ~^ image[22][13])} + {7'd0,(kernel[0][4] ~^ image[22][14])} + {7'd0,(kernel[1][0] ~^ image[23][10])} + {7'd0,(kernel[1][1] ~^ image[23][11])} + {7'd0,(kernel[1][2] ~^ image[23][12])} + {7'd0,(kernel[1][3] ~^ image[23][13])} + {7'd0,(kernel[1][4] ~^ image[23][14])} + {7'd0,(kernel[2][0] ~^ image[24][10])} + {7'd0,(kernel[2][1] ~^ image[24][11])} + {7'd0,(kernel[2][2] ~^ image[24][12])} + {7'd0,(kernel[2][3] ~^ image[24][13])} + {7'd0,(kernel[2][4] ~^ image[24][14])} + {7'd0,(kernel[3][0] ~^ image[25][10])} + {7'd0,(kernel[3][1] ~^ image[25][11])} + {7'd0,(kernel[3][2] ~^ image[25][12])} + {7'd0,(kernel[3][3] ~^ image[25][13])} + {7'd0,(kernel[3][4] ~^ image[25][14])} + {7'd0,(kernel[4][0] ~^ image[26][10])} + {7'd0,(kernel[4][1] ~^ image[26][11])} + {7'd0,(kernel[4][2] ~^ image[26][12])} + {7'd0,(kernel[4][3] ~^ image[26][13])} + {7'd0,(kernel[4][4] ~^ image[26][14])};
assign out_fmap[22][11][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[22][11])} + {7'd0,(kernel[0][1] ~^ image[22][12])} + {7'd0,(kernel[0][2] ~^ image[22][13])} + {7'd0,(kernel[0][3] ~^ image[22][14])} + {7'd0,(kernel[0][4] ~^ image[22][15])} + {7'd0,(kernel[1][0] ~^ image[23][11])} + {7'd0,(kernel[1][1] ~^ image[23][12])} + {7'd0,(kernel[1][2] ~^ image[23][13])} + {7'd0,(kernel[1][3] ~^ image[23][14])} + {7'd0,(kernel[1][4] ~^ image[23][15])} + {7'd0,(kernel[2][0] ~^ image[24][11])} + {7'd0,(kernel[2][1] ~^ image[24][12])} + {7'd0,(kernel[2][2] ~^ image[24][13])} + {7'd0,(kernel[2][3] ~^ image[24][14])} + {7'd0,(kernel[2][4] ~^ image[24][15])} + {7'd0,(kernel[3][0] ~^ image[25][11])} + {7'd0,(kernel[3][1] ~^ image[25][12])} + {7'd0,(kernel[3][2] ~^ image[25][13])} + {7'd0,(kernel[3][3] ~^ image[25][14])} + {7'd0,(kernel[3][4] ~^ image[25][15])} + {7'd0,(kernel[4][0] ~^ image[26][11])} + {7'd0,(kernel[4][1] ~^ image[26][12])} + {7'd0,(kernel[4][2] ~^ image[26][13])} + {7'd0,(kernel[4][3] ~^ image[26][14])} + {7'd0,(kernel[4][4] ~^ image[26][15])};
assign out_fmap[22][12][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[22][12])} + {7'd0,(kernel[0][1] ~^ image[22][13])} + {7'd0,(kernel[0][2] ~^ image[22][14])} + {7'd0,(kernel[0][3] ~^ image[22][15])} + {7'd0,(kernel[0][4] ~^ image[22][16])} + {7'd0,(kernel[1][0] ~^ image[23][12])} + {7'd0,(kernel[1][1] ~^ image[23][13])} + {7'd0,(kernel[1][2] ~^ image[23][14])} + {7'd0,(kernel[1][3] ~^ image[23][15])} + {7'd0,(kernel[1][4] ~^ image[23][16])} + {7'd0,(kernel[2][0] ~^ image[24][12])} + {7'd0,(kernel[2][1] ~^ image[24][13])} + {7'd0,(kernel[2][2] ~^ image[24][14])} + {7'd0,(kernel[2][3] ~^ image[24][15])} + {7'd0,(kernel[2][4] ~^ image[24][16])} + {7'd0,(kernel[3][0] ~^ image[25][12])} + {7'd0,(kernel[3][1] ~^ image[25][13])} + {7'd0,(kernel[3][2] ~^ image[25][14])} + {7'd0,(kernel[3][3] ~^ image[25][15])} + {7'd0,(kernel[3][4] ~^ image[25][16])} + {7'd0,(kernel[4][0] ~^ image[26][12])} + {7'd0,(kernel[4][1] ~^ image[26][13])} + {7'd0,(kernel[4][2] ~^ image[26][14])} + {7'd0,(kernel[4][3] ~^ image[26][15])} + {7'd0,(kernel[4][4] ~^ image[26][16])};
assign out_fmap[22][13][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[22][13])} + {7'd0,(kernel[0][1] ~^ image[22][14])} + {7'd0,(kernel[0][2] ~^ image[22][15])} + {7'd0,(kernel[0][3] ~^ image[22][16])} + {7'd0,(kernel[0][4] ~^ image[22][17])} + {7'd0,(kernel[1][0] ~^ image[23][13])} + {7'd0,(kernel[1][1] ~^ image[23][14])} + {7'd0,(kernel[1][2] ~^ image[23][15])} + {7'd0,(kernel[1][3] ~^ image[23][16])} + {7'd0,(kernel[1][4] ~^ image[23][17])} + {7'd0,(kernel[2][0] ~^ image[24][13])} + {7'd0,(kernel[2][1] ~^ image[24][14])} + {7'd0,(kernel[2][2] ~^ image[24][15])} + {7'd0,(kernel[2][3] ~^ image[24][16])} + {7'd0,(kernel[2][4] ~^ image[24][17])} + {7'd0,(kernel[3][0] ~^ image[25][13])} + {7'd0,(kernel[3][1] ~^ image[25][14])} + {7'd0,(kernel[3][2] ~^ image[25][15])} + {7'd0,(kernel[3][3] ~^ image[25][16])} + {7'd0,(kernel[3][4] ~^ image[25][17])} + {7'd0,(kernel[4][0] ~^ image[26][13])} + {7'd0,(kernel[4][1] ~^ image[26][14])} + {7'd0,(kernel[4][2] ~^ image[26][15])} + {7'd0,(kernel[4][3] ~^ image[26][16])} + {7'd0,(kernel[4][4] ~^ image[26][17])};
assign out_fmap[22][14][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[22][14])} + {7'd0,(kernel[0][1] ~^ image[22][15])} + {7'd0,(kernel[0][2] ~^ image[22][16])} + {7'd0,(kernel[0][3] ~^ image[22][17])} + {7'd0,(kernel[0][4] ~^ image[22][18])} + {7'd0,(kernel[1][0] ~^ image[23][14])} + {7'd0,(kernel[1][1] ~^ image[23][15])} + {7'd0,(kernel[1][2] ~^ image[23][16])} + {7'd0,(kernel[1][3] ~^ image[23][17])} + {7'd0,(kernel[1][4] ~^ image[23][18])} + {7'd0,(kernel[2][0] ~^ image[24][14])} + {7'd0,(kernel[2][1] ~^ image[24][15])} + {7'd0,(kernel[2][2] ~^ image[24][16])} + {7'd0,(kernel[2][3] ~^ image[24][17])} + {7'd0,(kernel[2][4] ~^ image[24][18])} + {7'd0,(kernel[3][0] ~^ image[25][14])} + {7'd0,(kernel[3][1] ~^ image[25][15])} + {7'd0,(kernel[3][2] ~^ image[25][16])} + {7'd0,(kernel[3][3] ~^ image[25][17])} + {7'd0,(kernel[3][4] ~^ image[25][18])} + {7'd0,(kernel[4][0] ~^ image[26][14])} + {7'd0,(kernel[4][1] ~^ image[26][15])} + {7'd0,(kernel[4][2] ~^ image[26][16])} + {7'd0,(kernel[4][3] ~^ image[26][17])} + {7'd0,(kernel[4][4] ~^ image[26][18])};
assign out_fmap[22][15][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[22][15])} + {7'd0,(kernel[0][1] ~^ image[22][16])} + {7'd0,(kernel[0][2] ~^ image[22][17])} + {7'd0,(kernel[0][3] ~^ image[22][18])} + {7'd0,(kernel[0][4] ~^ image[22][19])} + {7'd0,(kernel[1][0] ~^ image[23][15])} + {7'd0,(kernel[1][1] ~^ image[23][16])} + {7'd0,(kernel[1][2] ~^ image[23][17])} + {7'd0,(kernel[1][3] ~^ image[23][18])} + {7'd0,(kernel[1][4] ~^ image[23][19])} + {7'd0,(kernel[2][0] ~^ image[24][15])} + {7'd0,(kernel[2][1] ~^ image[24][16])} + {7'd0,(kernel[2][2] ~^ image[24][17])} + {7'd0,(kernel[2][3] ~^ image[24][18])} + {7'd0,(kernel[2][4] ~^ image[24][19])} + {7'd0,(kernel[3][0] ~^ image[25][15])} + {7'd0,(kernel[3][1] ~^ image[25][16])} + {7'd0,(kernel[3][2] ~^ image[25][17])} + {7'd0,(kernel[3][3] ~^ image[25][18])} + {7'd0,(kernel[3][4] ~^ image[25][19])} + {7'd0,(kernel[4][0] ~^ image[26][15])} + {7'd0,(kernel[4][1] ~^ image[26][16])} + {7'd0,(kernel[4][2] ~^ image[26][17])} + {7'd0,(kernel[4][3] ~^ image[26][18])} + {7'd0,(kernel[4][4] ~^ image[26][19])};
assign out_fmap[22][16][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[22][16])} + {7'd0,(kernel[0][1] ~^ image[22][17])} + {7'd0,(kernel[0][2] ~^ image[22][18])} + {7'd0,(kernel[0][3] ~^ image[22][19])} + {7'd0,(kernel[0][4] ~^ image[22][20])} + {7'd0,(kernel[1][0] ~^ image[23][16])} + {7'd0,(kernel[1][1] ~^ image[23][17])} + {7'd0,(kernel[1][2] ~^ image[23][18])} + {7'd0,(kernel[1][3] ~^ image[23][19])} + {7'd0,(kernel[1][4] ~^ image[23][20])} + {7'd0,(kernel[2][0] ~^ image[24][16])} + {7'd0,(kernel[2][1] ~^ image[24][17])} + {7'd0,(kernel[2][2] ~^ image[24][18])} + {7'd0,(kernel[2][3] ~^ image[24][19])} + {7'd0,(kernel[2][4] ~^ image[24][20])} + {7'd0,(kernel[3][0] ~^ image[25][16])} + {7'd0,(kernel[3][1] ~^ image[25][17])} + {7'd0,(kernel[3][2] ~^ image[25][18])} + {7'd0,(kernel[3][3] ~^ image[25][19])} + {7'd0,(kernel[3][4] ~^ image[25][20])} + {7'd0,(kernel[4][0] ~^ image[26][16])} + {7'd0,(kernel[4][1] ~^ image[26][17])} + {7'd0,(kernel[4][2] ~^ image[26][18])} + {7'd0,(kernel[4][3] ~^ image[26][19])} + {7'd0,(kernel[4][4] ~^ image[26][20])};
assign out_fmap[22][17][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[22][17])} + {7'd0,(kernel[0][1] ~^ image[22][18])} + {7'd0,(kernel[0][2] ~^ image[22][19])} + {7'd0,(kernel[0][3] ~^ image[22][20])} + {7'd0,(kernel[0][4] ~^ image[22][21])} + {7'd0,(kernel[1][0] ~^ image[23][17])} + {7'd0,(kernel[1][1] ~^ image[23][18])} + {7'd0,(kernel[1][2] ~^ image[23][19])} + {7'd0,(kernel[1][3] ~^ image[23][20])} + {7'd0,(kernel[1][4] ~^ image[23][21])} + {7'd0,(kernel[2][0] ~^ image[24][17])} + {7'd0,(kernel[2][1] ~^ image[24][18])} + {7'd0,(kernel[2][2] ~^ image[24][19])} + {7'd0,(kernel[2][3] ~^ image[24][20])} + {7'd0,(kernel[2][4] ~^ image[24][21])} + {7'd0,(kernel[3][0] ~^ image[25][17])} + {7'd0,(kernel[3][1] ~^ image[25][18])} + {7'd0,(kernel[3][2] ~^ image[25][19])} + {7'd0,(kernel[3][3] ~^ image[25][20])} + {7'd0,(kernel[3][4] ~^ image[25][21])} + {7'd0,(kernel[4][0] ~^ image[26][17])} + {7'd0,(kernel[4][1] ~^ image[26][18])} + {7'd0,(kernel[4][2] ~^ image[26][19])} + {7'd0,(kernel[4][3] ~^ image[26][20])} + {7'd0,(kernel[4][4] ~^ image[26][21])};
assign out_fmap[22][18][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[22][18])} + {7'd0,(kernel[0][1] ~^ image[22][19])} + {7'd0,(kernel[0][2] ~^ image[22][20])} + {7'd0,(kernel[0][3] ~^ image[22][21])} + {7'd0,(kernel[0][4] ~^ image[22][22])} + {7'd0,(kernel[1][0] ~^ image[23][18])} + {7'd0,(kernel[1][1] ~^ image[23][19])} + {7'd0,(kernel[1][2] ~^ image[23][20])} + {7'd0,(kernel[1][3] ~^ image[23][21])} + {7'd0,(kernel[1][4] ~^ image[23][22])} + {7'd0,(kernel[2][0] ~^ image[24][18])} + {7'd0,(kernel[2][1] ~^ image[24][19])} + {7'd0,(kernel[2][2] ~^ image[24][20])} + {7'd0,(kernel[2][3] ~^ image[24][21])} + {7'd0,(kernel[2][4] ~^ image[24][22])} + {7'd0,(kernel[3][0] ~^ image[25][18])} + {7'd0,(kernel[3][1] ~^ image[25][19])} + {7'd0,(kernel[3][2] ~^ image[25][20])} + {7'd0,(kernel[3][3] ~^ image[25][21])} + {7'd0,(kernel[3][4] ~^ image[25][22])} + {7'd0,(kernel[4][0] ~^ image[26][18])} + {7'd0,(kernel[4][1] ~^ image[26][19])} + {7'd0,(kernel[4][2] ~^ image[26][20])} + {7'd0,(kernel[4][3] ~^ image[26][21])} + {7'd0,(kernel[4][4] ~^ image[26][22])};
assign out_fmap[22][19][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[22][19])} + {7'd0,(kernel[0][1] ~^ image[22][20])} + {7'd0,(kernel[0][2] ~^ image[22][21])} + {7'd0,(kernel[0][3] ~^ image[22][22])} + {7'd0,(kernel[0][4] ~^ image[22][23])} + {7'd0,(kernel[1][0] ~^ image[23][19])} + {7'd0,(kernel[1][1] ~^ image[23][20])} + {7'd0,(kernel[1][2] ~^ image[23][21])} + {7'd0,(kernel[1][3] ~^ image[23][22])} + {7'd0,(kernel[1][4] ~^ image[23][23])} + {7'd0,(kernel[2][0] ~^ image[24][19])} + {7'd0,(kernel[2][1] ~^ image[24][20])} + {7'd0,(kernel[2][2] ~^ image[24][21])} + {7'd0,(kernel[2][3] ~^ image[24][22])} + {7'd0,(kernel[2][4] ~^ image[24][23])} + {7'd0,(kernel[3][0] ~^ image[25][19])} + {7'd0,(kernel[3][1] ~^ image[25][20])} + {7'd0,(kernel[3][2] ~^ image[25][21])} + {7'd0,(kernel[3][3] ~^ image[25][22])} + {7'd0,(kernel[3][4] ~^ image[25][23])} + {7'd0,(kernel[4][0] ~^ image[26][19])} + {7'd0,(kernel[4][1] ~^ image[26][20])} + {7'd0,(kernel[4][2] ~^ image[26][21])} + {7'd0,(kernel[4][3] ~^ image[26][22])} + {7'd0,(kernel[4][4] ~^ image[26][23])};
assign out_fmap[22][20][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[22][20])} + {7'd0,(kernel[0][1] ~^ image[22][21])} + {7'd0,(kernel[0][2] ~^ image[22][22])} + {7'd0,(kernel[0][3] ~^ image[22][23])} + {7'd0,(kernel[0][4] ~^ image[22][24])} + {7'd0,(kernel[1][0] ~^ image[23][20])} + {7'd0,(kernel[1][1] ~^ image[23][21])} + {7'd0,(kernel[1][2] ~^ image[23][22])} + {7'd0,(kernel[1][3] ~^ image[23][23])} + {7'd0,(kernel[1][4] ~^ image[23][24])} + {7'd0,(kernel[2][0] ~^ image[24][20])} + {7'd0,(kernel[2][1] ~^ image[24][21])} + {7'd0,(kernel[2][2] ~^ image[24][22])} + {7'd0,(kernel[2][3] ~^ image[24][23])} + {7'd0,(kernel[2][4] ~^ image[24][24])} + {7'd0,(kernel[3][0] ~^ image[25][20])} + {7'd0,(kernel[3][1] ~^ image[25][21])} + {7'd0,(kernel[3][2] ~^ image[25][22])} + {7'd0,(kernel[3][3] ~^ image[25][23])} + {7'd0,(kernel[3][4] ~^ image[25][24])} + {7'd0,(kernel[4][0] ~^ image[26][20])} + {7'd0,(kernel[4][1] ~^ image[26][21])} + {7'd0,(kernel[4][2] ~^ image[26][22])} + {7'd0,(kernel[4][3] ~^ image[26][23])} + {7'd0,(kernel[4][4] ~^ image[26][24])};
assign out_fmap[22][21][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[22][21])} + {7'd0,(kernel[0][1] ~^ image[22][22])} + {7'd0,(kernel[0][2] ~^ image[22][23])} + {7'd0,(kernel[0][3] ~^ image[22][24])} + {7'd0,(kernel[0][4] ~^ image[22][25])} + {7'd0,(kernel[1][0] ~^ image[23][21])} + {7'd0,(kernel[1][1] ~^ image[23][22])} + {7'd0,(kernel[1][2] ~^ image[23][23])} + {7'd0,(kernel[1][3] ~^ image[23][24])} + {7'd0,(kernel[1][4] ~^ image[23][25])} + {7'd0,(kernel[2][0] ~^ image[24][21])} + {7'd0,(kernel[2][1] ~^ image[24][22])} + {7'd0,(kernel[2][2] ~^ image[24][23])} + {7'd0,(kernel[2][3] ~^ image[24][24])} + {7'd0,(kernel[2][4] ~^ image[24][25])} + {7'd0,(kernel[3][0] ~^ image[25][21])} + {7'd0,(kernel[3][1] ~^ image[25][22])} + {7'd0,(kernel[3][2] ~^ image[25][23])} + {7'd0,(kernel[3][3] ~^ image[25][24])} + {7'd0,(kernel[3][4] ~^ image[25][25])} + {7'd0,(kernel[4][0] ~^ image[26][21])} + {7'd0,(kernel[4][1] ~^ image[26][22])} + {7'd0,(kernel[4][2] ~^ image[26][23])} + {7'd0,(kernel[4][3] ~^ image[26][24])} + {7'd0,(kernel[4][4] ~^ image[26][25])};
assign out_fmap[22][22][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[22][22])} + {7'd0,(kernel[0][1] ~^ image[22][23])} + {7'd0,(kernel[0][2] ~^ image[22][24])} + {7'd0,(kernel[0][3] ~^ image[22][25])} + {7'd0,(kernel[0][4] ~^ image[22][26])} + {7'd0,(kernel[1][0] ~^ image[23][22])} + {7'd0,(kernel[1][1] ~^ image[23][23])} + {7'd0,(kernel[1][2] ~^ image[23][24])} + {7'd0,(kernel[1][3] ~^ image[23][25])} + {7'd0,(kernel[1][4] ~^ image[23][26])} + {7'd0,(kernel[2][0] ~^ image[24][22])} + {7'd0,(kernel[2][1] ~^ image[24][23])} + {7'd0,(kernel[2][2] ~^ image[24][24])} + {7'd0,(kernel[2][3] ~^ image[24][25])} + {7'd0,(kernel[2][4] ~^ image[24][26])} + {7'd0,(kernel[3][0] ~^ image[25][22])} + {7'd0,(kernel[3][1] ~^ image[25][23])} + {7'd0,(kernel[3][2] ~^ image[25][24])} + {7'd0,(kernel[3][3] ~^ image[25][25])} + {7'd0,(kernel[3][4] ~^ image[25][26])} + {7'd0,(kernel[4][0] ~^ image[26][22])} + {7'd0,(kernel[4][1] ~^ image[26][23])} + {7'd0,(kernel[4][2] ~^ image[26][24])} + {7'd0,(kernel[4][3] ~^ image[26][25])} + {7'd0,(kernel[4][4] ~^ image[26][26])};
assign out_fmap[22][23][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[22][23])} + {7'd0,(kernel[0][1] ~^ image[22][24])} + {7'd0,(kernel[0][2] ~^ image[22][25])} + {7'd0,(kernel[0][3] ~^ image[22][26])} + {7'd0,(kernel[0][4] ~^ image[22][27])} + {7'd0,(kernel[1][0] ~^ image[23][23])} + {7'd0,(kernel[1][1] ~^ image[23][24])} + {7'd0,(kernel[1][2] ~^ image[23][25])} + {7'd0,(kernel[1][3] ~^ image[23][26])} + {7'd0,(kernel[1][4] ~^ image[23][27])} + {7'd0,(kernel[2][0] ~^ image[24][23])} + {7'd0,(kernel[2][1] ~^ image[24][24])} + {7'd0,(kernel[2][2] ~^ image[24][25])} + {7'd0,(kernel[2][3] ~^ image[24][26])} + {7'd0,(kernel[2][4] ~^ image[24][27])} + {7'd0,(kernel[3][0] ~^ image[25][23])} + {7'd0,(kernel[3][1] ~^ image[25][24])} + {7'd0,(kernel[3][2] ~^ image[25][25])} + {7'd0,(kernel[3][3] ~^ image[25][26])} + {7'd0,(kernel[3][4] ~^ image[25][27])} + {7'd0,(kernel[4][0] ~^ image[26][23])} + {7'd0,(kernel[4][1] ~^ image[26][24])} + {7'd0,(kernel[4][2] ~^ image[26][25])} + {7'd0,(kernel[4][3] ~^ image[26][26])} + {7'd0,(kernel[4][4] ~^ image[26][27])};
assign out_fmap[23][0][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[23][0])} + {7'd0,(kernel[0][1] ~^ image[23][1])} + {7'd0,(kernel[0][2] ~^ image[23][2])} + {7'd0,(kernel[0][3] ~^ image[23][3])} + {7'd0,(kernel[0][4] ~^ image[23][4])} + {7'd0,(kernel[1][0] ~^ image[24][0])} + {7'd0,(kernel[1][1] ~^ image[24][1])} + {7'd0,(kernel[1][2] ~^ image[24][2])} + {7'd0,(kernel[1][3] ~^ image[24][3])} + {7'd0,(kernel[1][4] ~^ image[24][4])} + {7'd0,(kernel[2][0] ~^ image[25][0])} + {7'd0,(kernel[2][1] ~^ image[25][1])} + {7'd0,(kernel[2][2] ~^ image[25][2])} + {7'd0,(kernel[2][3] ~^ image[25][3])} + {7'd0,(kernel[2][4] ~^ image[25][4])} + {7'd0,(kernel[3][0] ~^ image[26][0])} + {7'd0,(kernel[3][1] ~^ image[26][1])} + {7'd0,(kernel[3][2] ~^ image[26][2])} + {7'd0,(kernel[3][3] ~^ image[26][3])} + {7'd0,(kernel[3][4] ~^ image[26][4])} + {7'd0,(kernel[4][0] ~^ image[27][0])} + {7'd0,(kernel[4][1] ~^ image[27][1])} + {7'd0,(kernel[4][2] ~^ image[27][2])} + {7'd0,(kernel[4][3] ~^ image[27][3])} + {7'd0,(kernel[4][4] ~^ image[27][4])};
assign out_fmap[23][1][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[23][1])} + {7'd0,(kernel[0][1] ~^ image[23][2])} + {7'd0,(kernel[0][2] ~^ image[23][3])} + {7'd0,(kernel[0][3] ~^ image[23][4])} + {7'd0,(kernel[0][4] ~^ image[23][5])} + {7'd0,(kernel[1][0] ~^ image[24][1])} + {7'd0,(kernel[1][1] ~^ image[24][2])} + {7'd0,(kernel[1][2] ~^ image[24][3])} + {7'd0,(kernel[1][3] ~^ image[24][4])} + {7'd0,(kernel[1][4] ~^ image[24][5])} + {7'd0,(kernel[2][0] ~^ image[25][1])} + {7'd0,(kernel[2][1] ~^ image[25][2])} + {7'd0,(kernel[2][2] ~^ image[25][3])} + {7'd0,(kernel[2][3] ~^ image[25][4])} + {7'd0,(kernel[2][4] ~^ image[25][5])} + {7'd0,(kernel[3][0] ~^ image[26][1])} + {7'd0,(kernel[3][1] ~^ image[26][2])} + {7'd0,(kernel[3][2] ~^ image[26][3])} + {7'd0,(kernel[3][3] ~^ image[26][4])} + {7'd0,(kernel[3][4] ~^ image[26][5])} + {7'd0,(kernel[4][0] ~^ image[27][1])} + {7'd0,(kernel[4][1] ~^ image[27][2])} + {7'd0,(kernel[4][2] ~^ image[27][3])} + {7'd0,(kernel[4][3] ~^ image[27][4])} + {7'd0,(kernel[4][4] ~^ image[27][5])};
assign out_fmap[23][2][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[23][2])} + {7'd0,(kernel[0][1] ~^ image[23][3])} + {7'd0,(kernel[0][2] ~^ image[23][4])} + {7'd0,(kernel[0][3] ~^ image[23][5])} + {7'd0,(kernel[0][4] ~^ image[23][6])} + {7'd0,(kernel[1][0] ~^ image[24][2])} + {7'd0,(kernel[1][1] ~^ image[24][3])} + {7'd0,(kernel[1][2] ~^ image[24][4])} + {7'd0,(kernel[1][3] ~^ image[24][5])} + {7'd0,(kernel[1][4] ~^ image[24][6])} + {7'd0,(kernel[2][0] ~^ image[25][2])} + {7'd0,(kernel[2][1] ~^ image[25][3])} + {7'd0,(kernel[2][2] ~^ image[25][4])} + {7'd0,(kernel[2][3] ~^ image[25][5])} + {7'd0,(kernel[2][4] ~^ image[25][6])} + {7'd0,(kernel[3][0] ~^ image[26][2])} + {7'd0,(kernel[3][1] ~^ image[26][3])} + {7'd0,(kernel[3][2] ~^ image[26][4])} + {7'd0,(kernel[3][3] ~^ image[26][5])} + {7'd0,(kernel[3][4] ~^ image[26][6])} + {7'd0,(kernel[4][0] ~^ image[27][2])} + {7'd0,(kernel[4][1] ~^ image[27][3])} + {7'd0,(kernel[4][2] ~^ image[27][4])} + {7'd0,(kernel[4][3] ~^ image[27][5])} + {7'd0,(kernel[4][4] ~^ image[27][6])};
assign out_fmap[23][3][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[23][3])} + {7'd0,(kernel[0][1] ~^ image[23][4])} + {7'd0,(kernel[0][2] ~^ image[23][5])} + {7'd0,(kernel[0][3] ~^ image[23][6])} + {7'd0,(kernel[0][4] ~^ image[23][7])} + {7'd0,(kernel[1][0] ~^ image[24][3])} + {7'd0,(kernel[1][1] ~^ image[24][4])} + {7'd0,(kernel[1][2] ~^ image[24][5])} + {7'd0,(kernel[1][3] ~^ image[24][6])} + {7'd0,(kernel[1][4] ~^ image[24][7])} + {7'd0,(kernel[2][0] ~^ image[25][3])} + {7'd0,(kernel[2][1] ~^ image[25][4])} + {7'd0,(kernel[2][2] ~^ image[25][5])} + {7'd0,(kernel[2][3] ~^ image[25][6])} + {7'd0,(kernel[2][4] ~^ image[25][7])} + {7'd0,(kernel[3][0] ~^ image[26][3])} + {7'd0,(kernel[3][1] ~^ image[26][4])} + {7'd0,(kernel[3][2] ~^ image[26][5])} + {7'd0,(kernel[3][3] ~^ image[26][6])} + {7'd0,(kernel[3][4] ~^ image[26][7])} + {7'd0,(kernel[4][0] ~^ image[27][3])} + {7'd0,(kernel[4][1] ~^ image[27][4])} + {7'd0,(kernel[4][2] ~^ image[27][5])} + {7'd0,(kernel[4][3] ~^ image[27][6])} + {7'd0,(kernel[4][4] ~^ image[27][7])};
assign out_fmap[23][4][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[23][4])} + {7'd0,(kernel[0][1] ~^ image[23][5])} + {7'd0,(kernel[0][2] ~^ image[23][6])} + {7'd0,(kernel[0][3] ~^ image[23][7])} + {7'd0,(kernel[0][4] ~^ image[23][8])} + {7'd0,(kernel[1][0] ~^ image[24][4])} + {7'd0,(kernel[1][1] ~^ image[24][5])} + {7'd0,(kernel[1][2] ~^ image[24][6])} + {7'd0,(kernel[1][3] ~^ image[24][7])} + {7'd0,(kernel[1][4] ~^ image[24][8])} + {7'd0,(kernel[2][0] ~^ image[25][4])} + {7'd0,(kernel[2][1] ~^ image[25][5])} + {7'd0,(kernel[2][2] ~^ image[25][6])} + {7'd0,(kernel[2][3] ~^ image[25][7])} + {7'd0,(kernel[2][4] ~^ image[25][8])} + {7'd0,(kernel[3][0] ~^ image[26][4])} + {7'd0,(kernel[3][1] ~^ image[26][5])} + {7'd0,(kernel[3][2] ~^ image[26][6])} + {7'd0,(kernel[3][3] ~^ image[26][7])} + {7'd0,(kernel[3][4] ~^ image[26][8])} + {7'd0,(kernel[4][0] ~^ image[27][4])} + {7'd0,(kernel[4][1] ~^ image[27][5])} + {7'd0,(kernel[4][2] ~^ image[27][6])} + {7'd0,(kernel[4][3] ~^ image[27][7])} + {7'd0,(kernel[4][4] ~^ image[27][8])};
assign out_fmap[23][5][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[23][5])} + {7'd0,(kernel[0][1] ~^ image[23][6])} + {7'd0,(kernel[0][2] ~^ image[23][7])} + {7'd0,(kernel[0][3] ~^ image[23][8])} + {7'd0,(kernel[0][4] ~^ image[23][9])} + {7'd0,(kernel[1][0] ~^ image[24][5])} + {7'd0,(kernel[1][1] ~^ image[24][6])} + {7'd0,(kernel[1][2] ~^ image[24][7])} + {7'd0,(kernel[1][3] ~^ image[24][8])} + {7'd0,(kernel[1][4] ~^ image[24][9])} + {7'd0,(kernel[2][0] ~^ image[25][5])} + {7'd0,(kernel[2][1] ~^ image[25][6])} + {7'd0,(kernel[2][2] ~^ image[25][7])} + {7'd0,(kernel[2][3] ~^ image[25][8])} + {7'd0,(kernel[2][4] ~^ image[25][9])} + {7'd0,(kernel[3][0] ~^ image[26][5])} + {7'd0,(kernel[3][1] ~^ image[26][6])} + {7'd0,(kernel[3][2] ~^ image[26][7])} + {7'd0,(kernel[3][3] ~^ image[26][8])} + {7'd0,(kernel[3][4] ~^ image[26][9])} + {7'd0,(kernel[4][0] ~^ image[27][5])} + {7'd0,(kernel[4][1] ~^ image[27][6])} + {7'd0,(kernel[4][2] ~^ image[27][7])} + {7'd0,(kernel[4][3] ~^ image[27][8])} + {7'd0,(kernel[4][4] ~^ image[27][9])};
assign out_fmap[23][6][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[23][6])} + {7'd0,(kernel[0][1] ~^ image[23][7])} + {7'd0,(kernel[0][2] ~^ image[23][8])} + {7'd0,(kernel[0][3] ~^ image[23][9])} + {7'd0,(kernel[0][4] ~^ image[23][10])} + {7'd0,(kernel[1][0] ~^ image[24][6])} + {7'd0,(kernel[1][1] ~^ image[24][7])} + {7'd0,(kernel[1][2] ~^ image[24][8])} + {7'd0,(kernel[1][3] ~^ image[24][9])} + {7'd0,(kernel[1][4] ~^ image[24][10])} + {7'd0,(kernel[2][0] ~^ image[25][6])} + {7'd0,(kernel[2][1] ~^ image[25][7])} + {7'd0,(kernel[2][2] ~^ image[25][8])} + {7'd0,(kernel[2][3] ~^ image[25][9])} + {7'd0,(kernel[2][4] ~^ image[25][10])} + {7'd0,(kernel[3][0] ~^ image[26][6])} + {7'd0,(kernel[3][1] ~^ image[26][7])} + {7'd0,(kernel[3][2] ~^ image[26][8])} + {7'd0,(kernel[3][3] ~^ image[26][9])} + {7'd0,(kernel[3][4] ~^ image[26][10])} + {7'd0,(kernel[4][0] ~^ image[27][6])} + {7'd0,(kernel[4][1] ~^ image[27][7])} + {7'd0,(kernel[4][2] ~^ image[27][8])} + {7'd0,(kernel[4][3] ~^ image[27][9])} + {7'd0,(kernel[4][4] ~^ image[27][10])};
assign out_fmap[23][7][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[23][7])} + {7'd0,(kernel[0][1] ~^ image[23][8])} + {7'd0,(kernel[0][2] ~^ image[23][9])} + {7'd0,(kernel[0][3] ~^ image[23][10])} + {7'd0,(kernel[0][4] ~^ image[23][11])} + {7'd0,(kernel[1][0] ~^ image[24][7])} + {7'd0,(kernel[1][1] ~^ image[24][8])} + {7'd0,(kernel[1][2] ~^ image[24][9])} + {7'd0,(kernel[1][3] ~^ image[24][10])} + {7'd0,(kernel[1][4] ~^ image[24][11])} + {7'd0,(kernel[2][0] ~^ image[25][7])} + {7'd0,(kernel[2][1] ~^ image[25][8])} + {7'd0,(kernel[2][2] ~^ image[25][9])} + {7'd0,(kernel[2][3] ~^ image[25][10])} + {7'd0,(kernel[2][4] ~^ image[25][11])} + {7'd0,(kernel[3][0] ~^ image[26][7])} + {7'd0,(kernel[3][1] ~^ image[26][8])} + {7'd0,(kernel[3][2] ~^ image[26][9])} + {7'd0,(kernel[3][3] ~^ image[26][10])} + {7'd0,(kernel[3][4] ~^ image[26][11])} + {7'd0,(kernel[4][0] ~^ image[27][7])} + {7'd0,(kernel[4][1] ~^ image[27][8])} + {7'd0,(kernel[4][2] ~^ image[27][9])} + {7'd0,(kernel[4][3] ~^ image[27][10])} + {7'd0,(kernel[4][4] ~^ image[27][11])};
assign out_fmap[23][8][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[23][8])} + {7'd0,(kernel[0][1] ~^ image[23][9])} + {7'd0,(kernel[0][2] ~^ image[23][10])} + {7'd0,(kernel[0][3] ~^ image[23][11])} + {7'd0,(kernel[0][4] ~^ image[23][12])} + {7'd0,(kernel[1][0] ~^ image[24][8])} + {7'd0,(kernel[1][1] ~^ image[24][9])} + {7'd0,(kernel[1][2] ~^ image[24][10])} + {7'd0,(kernel[1][3] ~^ image[24][11])} + {7'd0,(kernel[1][4] ~^ image[24][12])} + {7'd0,(kernel[2][0] ~^ image[25][8])} + {7'd0,(kernel[2][1] ~^ image[25][9])} + {7'd0,(kernel[2][2] ~^ image[25][10])} + {7'd0,(kernel[2][3] ~^ image[25][11])} + {7'd0,(kernel[2][4] ~^ image[25][12])} + {7'd0,(kernel[3][0] ~^ image[26][8])} + {7'd0,(kernel[3][1] ~^ image[26][9])} + {7'd0,(kernel[3][2] ~^ image[26][10])} + {7'd0,(kernel[3][3] ~^ image[26][11])} + {7'd0,(kernel[3][4] ~^ image[26][12])} + {7'd0,(kernel[4][0] ~^ image[27][8])} + {7'd0,(kernel[4][1] ~^ image[27][9])} + {7'd0,(kernel[4][2] ~^ image[27][10])} + {7'd0,(kernel[4][3] ~^ image[27][11])} + {7'd0,(kernel[4][4] ~^ image[27][12])};
assign out_fmap[23][9][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[23][9])} + {7'd0,(kernel[0][1] ~^ image[23][10])} + {7'd0,(kernel[0][2] ~^ image[23][11])} + {7'd0,(kernel[0][3] ~^ image[23][12])} + {7'd0,(kernel[0][4] ~^ image[23][13])} + {7'd0,(kernel[1][0] ~^ image[24][9])} + {7'd0,(kernel[1][1] ~^ image[24][10])} + {7'd0,(kernel[1][2] ~^ image[24][11])} + {7'd0,(kernel[1][3] ~^ image[24][12])} + {7'd0,(kernel[1][4] ~^ image[24][13])} + {7'd0,(kernel[2][0] ~^ image[25][9])} + {7'd0,(kernel[2][1] ~^ image[25][10])} + {7'd0,(kernel[2][2] ~^ image[25][11])} + {7'd0,(kernel[2][3] ~^ image[25][12])} + {7'd0,(kernel[2][4] ~^ image[25][13])} + {7'd0,(kernel[3][0] ~^ image[26][9])} + {7'd0,(kernel[3][1] ~^ image[26][10])} + {7'd0,(kernel[3][2] ~^ image[26][11])} + {7'd0,(kernel[3][3] ~^ image[26][12])} + {7'd0,(kernel[3][4] ~^ image[26][13])} + {7'd0,(kernel[4][0] ~^ image[27][9])} + {7'd0,(kernel[4][1] ~^ image[27][10])} + {7'd0,(kernel[4][2] ~^ image[27][11])} + {7'd0,(kernel[4][3] ~^ image[27][12])} + {7'd0,(kernel[4][4] ~^ image[27][13])};
assign out_fmap[23][10][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[23][10])} + {7'd0,(kernel[0][1] ~^ image[23][11])} + {7'd0,(kernel[0][2] ~^ image[23][12])} + {7'd0,(kernel[0][3] ~^ image[23][13])} + {7'd0,(kernel[0][4] ~^ image[23][14])} + {7'd0,(kernel[1][0] ~^ image[24][10])} + {7'd0,(kernel[1][1] ~^ image[24][11])} + {7'd0,(kernel[1][2] ~^ image[24][12])} + {7'd0,(kernel[1][3] ~^ image[24][13])} + {7'd0,(kernel[1][4] ~^ image[24][14])} + {7'd0,(kernel[2][0] ~^ image[25][10])} + {7'd0,(kernel[2][1] ~^ image[25][11])} + {7'd0,(kernel[2][2] ~^ image[25][12])} + {7'd0,(kernel[2][3] ~^ image[25][13])} + {7'd0,(kernel[2][4] ~^ image[25][14])} + {7'd0,(kernel[3][0] ~^ image[26][10])} + {7'd0,(kernel[3][1] ~^ image[26][11])} + {7'd0,(kernel[3][2] ~^ image[26][12])} + {7'd0,(kernel[3][3] ~^ image[26][13])} + {7'd0,(kernel[3][4] ~^ image[26][14])} + {7'd0,(kernel[4][0] ~^ image[27][10])} + {7'd0,(kernel[4][1] ~^ image[27][11])} + {7'd0,(kernel[4][2] ~^ image[27][12])} + {7'd0,(kernel[4][3] ~^ image[27][13])} + {7'd0,(kernel[4][4] ~^ image[27][14])};
assign out_fmap[23][11][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[23][11])} + {7'd0,(kernel[0][1] ~^ image[23][12])} + {7'd0,(kernel[0][2] ~^ image[23][13])} + {7'd0,(kernel[0][3] ~^ image[23][14])} + {7'd0,(kernel[0][4] ~^ image[23][15])} + {7'd0,(kernel[1][0] ~^ image[24][11])} + {7'd0,(kernel[1][1] ~^ image[24][12])} + {7'd0,(kernel[1][2] ~^ image[24][13])} + {7'd0,(kernel[1][3] ~^ image[24][14])} + {7'd0,(kernel[1][4] ~^ image[24][15])} + {7'd0,(kernel[2][0] ~^ image[25][11])} + {7'd0,(kernel[2][1] ~^ image[25][12])} + {7'd0,(kernel[2][2] ~^ image[25][13])} + {7'd0,(kernel[2][3] ~^ image[25][14])} + {7'd0,(kernel[2][4] ~^ image[25][15])} + {7'd0,(kernel[3][0] ~^ image[26][11])} + {7'd0,(kernel[3][1] ~^ image[26][12])} + {7'd0,(kernel[3][2] ~^ image[26][13])} + {7'd0,(kernel[3][3] ~^ image[26][14])} + {7'd0,(kernel[3][4] ~^ image[26][15])} + {7'd0,(kernel[4][0] ~^ image[27][11])} + {7'd0,(kernel[4][1] ~^ image[27][12])} + {7'd0,(kernel[4][2] ~^ image[27][13])} + {7'd0,(kernel[4][3] ~^ image[27][14])} + {7'd0,(kernel[4][4] ~^ image[27][15])};
assign out_fmap[23][12][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[23][12])} + {7'd0,(kernel[0][1] ~^ image[23][13])} + {7'd0,(kernel[0][2] ~^ image[23][14])} + {7'd0,(kernel[0][3] ~^ image[23][15])} + {7'd0,(kernel[0][4] ~^ image[23][16])} + {7'd0,(kernel[1][0] ~^ image[24][12])} + {7'd0,(kernel[1][1] ~^ image[24][13])} + {7'd0,(kernel[1][2] ~^ image[24][14])} + {7'd0,(kernel[1][3] ~^ image[24][15])} + {7'd0,(kernel[1][4] ~^ image[24][16])} + {7'd0,(kernel[2][0] ~^ image[25][12])} + {7'd0,(kernel[2][1] ~^ image[25][13])} + {7'd0,(kernel[2][2] ~^ image[25][14])} + {7'd0,(kernel[2][3] ~^ image[25][15])} + {7'd0,(kernel[2][4] ~^ image[25][16])} + {7'd0,(kernel[3][0] ~^ image[26][12])} + {7'd0,(kernel[3][1] ~^ image[26][13])} + {7'd0,(kernel[3][2] ~^ image[26][14])} + {7'd0,(kernel[3][3] ~^ image[26][15])} + {7'd0,(kernel[3][4] ~^ image[26][16])} + {7'd0,(kernel[4][0] ~^ image[27][12])} + {7'd0,(kernel[4][1] ~^ image[27][13])} + {7'd0,(kernel[4][2] ~^ image[27][14])} + {7'd0,(kernel[4][3] ~^ image[27][15])} + {7'd0,(kernel[4][4] ~^ image[27][16])};
assign out_fmap[23][13][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[23][13])} + {7'd0,(kernel[0][1] ~^ image[23][14])} + {7'd0,(kernel[0][2] ~^ image[23][15])} + {7'd0,(kernel[0][3] ~^ image[23][16])} + {7'd0,(kernel[0][4] ~^ image[23][17])} + {7'd0,(kernel[1][0] ~^ image[24][13])} + {7'd0,(kernel[1][1] ~^ image[24][14])} + {7'd0,(kernel[1][2] ~^ image[24][15])} + {7'd0,(kernel[1][3] ~^ image[24][16])} + {7'd0,(kernel[1][4] ~^ image[24][17])} + {7'd0,(kernel[2][0] ~^ image[25][13])} + {7'd0,(kernel[2][1] ~^ image[25][14])} + {7'd0,(kernel[2][2] ~^ image[25][15])} + {7'd0,(kernel[2][3] ~^ image[25][16])} + {7'd0,(kernel[2][4] ~^ image[25][17])} + {7'd0,(kernel[3][0] ~^ image[26][13])} + {7'd0,(kernel[3][1] ~^ image[26][14])} + {7'd0,(kernel[3][2] ~^ image[26][15])} + {7'd0,(kernel[3][3] ~^ image[26][16])} + {7'd0,(kernel[3][4] ~^ image[26][17])} + {7'd0,(kernel[4][0] ~^ image[27][13])} + {7'd0,(kernel[4][1] ~^ image[27][14])} + {7'd0,(kernel[4][2] ~^ image[27][15])} + {7'd0,(kernel[4][3] ~^ image[27][16])} + {7'd0,(kernel[4][4] ~^ image[27][17])};
assign out_fmap[23][14][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[23][14])} + {7'd0,(kernel[0][1] ~^ image[23][15])} + {7'd0,(kernel[0][2] ~^ image[23][16])} + {7'd0,(kernel[0][3] ~^ image[23][17])} + {7'd0,(kernel[0][4] ~^ image[23][18])} + {7'd0,(kernel[1][0] ~^ image[24][14])} + {7'd0,(kernel[1][1] ~^ image[24][15])} + {7'd0,(kernel[1][2] ~^ image[24][16])} + {7'd0,(kernel[1][3] ~^ image[24][17])} + {7'd0,(kernel[1][4] ~^ image[24][18])} + {7'd0,(kernel[2][0] ~^ image[25][14])} + {7'd0,(kernel[2][1] ~^ image[25][15])} + {7'd0,(kernel[2][2] ~^ image[25][16])} + {7'd0,(kernel[2][3] ~^ image[25][17])} + {7'd0,(kernel[2][4] ~^ image[25][18])} + {7'd0,(kernel[3][0] ~^ image[26][14])} + {7'd0,(kernel[3][1] ~^ image[26][15])} + {7'd0,(kernel[3][2] ~^ image[26][16])} + {7'd0,(kernel[3][3] ~^ image[26][17])} + {7'd0,(kernel[3][4] ~^ image[26][18])} + {7'd0,(kernel[4][0] ~^ image[27][14])} + {7'd0,(kernel[4][1] ~^ image[27][15])} + {7'd0,(kernel[4][2] ~^ image[27][16])} + {7'd0,(kernel[4][3] ~^ image[27][17])} + {7'd0,(kernel[4][4] ~^ image[27][18])};
assign out_fmap[23][15][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[23][15])} + {7'd0,(kernel[0][1] ~^ image[23][16])} + {7'd0,(kernel[0][2] ~^ image[23][17])} + {7'd0,(kernel[0][3] ~^ image[23][18])} + {7'd0,(kernel[0][4] ~^ image[23][19])} + {7'd0,(kernel[1][0] ~^ image[24][15])} + {7'd0,(kernel[1][1] ~^ image[24][16])} + {7'd0,(kernel[1][2] ~^ image[24][17])} + {7'd0,(kernel[1][3] ~^ image[24][18])} + {7'd0,(kernel[1][4] ~^ image[24][19])} + {7'd0,(kernel[2][0] ~^ image[25][15])} + {7'd0,(kernel[2][1] ~^ image[25][16])} + {7'd0,(kernel[2][2] ~^ image[25][17])} + {7'd0,(kernel[2][3] ~^ image[25][18])} + {7'd0,(kernel[2][4] ~^ image[25][19])} + {7'd0,(kernel[3][0] ~^ image[26][15])} + {7'd0,(kernel[3][1] ~^ image[26][16])} + {7'd0,(kernel[3][2] ~^ image[26][17])} + {7'd0,(kernel[3][3] ~^ image[26][18])} + {7'd0,(kernel[3][4] ~^ image[26][19])} + {7'd0,(kernel[4][0] ~^ image[27][15])} + {7'd0,(kernel[4][1] ~^ image[27][16])} + {7'd0,(kernel[4][2] ~^ image[27][17])} + {7'd0,(kernel[4][3] ~^ image[27][18])} + {7'd0,(kernel[4][4] ~^ image[27][19])};
assign out_fmap[23][16][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[23][16])} + {7'd0,(kernel[0][1] ~^ image[23][17])} + {7'd0,(kernel[0][2] ~^ image[23][18])} + {7'd0,(kernel[0][3] ~^ image[23][19])} + {7'd0,(kernel[0][4] ~^ image[23][20])} + {7'd0,(kernel[1][0] ~^ image[24][16])} + {7'd0,(kernel[1][1] ~^ image[24][17])} + {7'd0,(kernel[1][2] ~^ image[24][18])} + {7'd0,(kernel[1][3] ~^ image[24][19])} + {7'd0,(kernel[1][4] ~^ image[24][20])} + {7'd0,(kernel[2][0] ~^ image[25][16])} + {7'd0,(kernel[2][1] ~^ image[25][17])} + {7'd0,(kernel[2][2] ~^ image[25][18])} + {7'd0,(kernel[2][3] ~^ image[25][19])} + {7'd0,(kernel[2][4] ~^ image[25][20])} + {7'd0,(kernel[3][0] ~^ image[26][16])} + {7'd0,(kernel[3][1] ~^ image[26][17])} + {7'd0,(kernel[3][2] ~^ image[26][18])} + {7'd0,(kernel[3][3] ~^ image[26][19])} + {7'd0,(kernel[3][4] ~^ image[26][20])} + {7'd0,(kernel[4][0] ~^ image[27][16])} + {7'd0,(kernel[4][1] ~^ image[27][17])} + {7'd0,(kernel[4][2] ~^ image[27][18])} + {7'd0,(kernel[4][3] ~^ image[27][19])} + {7'd0,(kernel[4][4] ~^ image[27][20])};
assign out_fmap[23][17][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[23][17])} + {7'd0,(kernel[0][1] ~^ image[23][18])} + {7'd0,(kernel[0][2] ~^ image[23][19])} + {7'd0,(kernel[0][3] ~^ image[23][20])} + {7'd0,(kernel[0][4] ~^ image[23][21])} + {7'd0,(kernel[1][0] ~^ image[24][17])} + {7'd0,(kernel[1][1] ~^ image[24][18])} + {7'd0,(kernel[1][2] ~^ image[24][19])} + {7'd0,(kernel[1][3] ~^ image[24][20])} + {7'd0,(kernel[1][4] ~^ image[24][21])} + {7'd0,(kernel[2][0] ~^ image[25][17])} + {7'd0,(kernel[2][1] ~^ image[25][18])} + {7'd0,(kernel[2][2] ~^ image[25][19])} + {7'd0,(kernel[2][3] ~^ image[25][20])} + {7'd0,(kernel[2][4] ~^ image[25][21])} + {7'd0,(kernel[3][0] ~^ image[26][17])} + {7'd0,(kernel[3][1] ~^ image[26][18])} + {7'd0,(kernel[3][2] ~^ image[26][19])} + {7'd0,(kernel[3][3] ~^ image[26][20])} + {7'd0,(kernel[3][4] ~^ image[26][21])} + {7'd0,(kernel[4][0] ~^ image[27][17])} + {7'd0,(kernel[4][1] ~^ image[27][18])} + {7'd0,(kernel[4][2] ~^ image[27][19])} + {7'd0,(kernel[4][3] ~^ image[27][20])} + {7'd0,(kernel[4][4] ~^ image[27][21])};
assign out_fmap[23][18][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[23][18])} + {7'd0,(kernel[0][1] ~^ image[23][19])} + {7'd0,(kernel[0][2] ~^ image[23][20])} + {7'd0,(kernel[0][3] ~^ image[23][21])} + {7'd0,(kernel[0][4] ~^ image[23][22])} + {7'd0,(kernel[1][0] ~^ image[24][18])} + {7'd0,(kernel[1][1] ~^ image[24][19])} + {7'd0,(kernel[1][2] ~^ image[24][20])} + {7'd0,(kernel[1][3] ~^ image[24][21])} + {7'd0,(kernel[1][4] ~^ image[24][22])} + {7'd0,(kernel[2][0] ~^ image[25][18])} + {7'd0,(kernel[2][1] ~^ image[25][19])} + {7'd0,(kernel[2][2] ~^ image[25][20])} + {7'd0,(kernel[2][3] ~^ image[25][21])} + {7'd0,(kernel[2][4] ~^ image[25][22])} + {7'd0,(kernel[3][0] ~^ image[26][18])} + {7'd0,(kernel[3][1] ~^ image[26][19])} + {7'd0,(kernel[3][2] ~^ image[26][20])} + {7'd0,(kernel[3][3] ~^ image[26][21])} + {7'd0,(kernel[3][4] ~^ image[26][22])} + {7'd0,(kernel[4][0] ~^ image[27][18])} + {7'd0,(kernel[4][1] ~^ image[27][19])} + {7'd0,(kernel[4][2] ~^ image[27][20])} + {7'd0,(kernel[4][3] ~^ image[27][21])} + {7'd0,(kernel[4][4] ~^ image[27][22])};
assign out_fmap[23][19][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[23][19])} + {7'd0,(kernel[0][1] ~^ image[23][20])} + {7'd0,(kernel[0][2] ~^ image[23][21])} + {7'd0,(kernel[0][3] ~^ image[23][22])} + {7'd0,(kernel[0][4] ~^ image[23][23])} + {7'd0,(kernel[1][0] ~^ image[24][19])} + {7'd0,(kernel[1][1] ~^ image[24][20])} + {7'd0,(kernel[1][2] ~^ image[24][21])} + {7'd0,(kernel[1][3] ~^ image[24][22])} + {7'd0,(kernel[1][4] ~^ image[24][23])} + {7'd0,(kernel[2][0] ~^ image[25][19])} + {7'd0,(kernel[2][1] ~^ image[25][20])} + {7'd0,(kernel[2][2] ~^ image[25][21])} + {7'd0,(kernel[2][3] ~^ image[25][22])} + {7'd0,(kernel[2][4] ~^ image[25][23])} + {7'd0,(kernel[3][0] ~^ image[26][19])} + {7'd0,(kernel[3][1] ~^ image[26][20])} + {7'd0,(kernel[3][2] ~^ image[26][21])} + {7'd0,(kernel[3][3] ~^ image[26][22])} + {7'd0,(kernel[3][4] ~^ image[26][23])} + {7'd0,(kernel[4][0] ~^ image[27][19])} + {7'd0,(kernel[4][1] ~^ image[27][20])} + {7'd0,(kernel[4][2] ~^ image[27][21])} + {7'd0,(kernel[4][3] ~^ image[27][22])} + {7'd0,(kernel[4][4] ~^ image[27][23])};
assign out_fmap[23][20][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[23][20])} + {7'd0,(kernel[0][1] ~^ image[23][21])} + {7'd0,(kernel[0][2] ~^ image[23][22])} + {7'd0,(kernel[0][3] ~^ image[23][23])} + {7'd0,(kernel[0][4] ~^ image[23][24])} + {7'd0,(kernel[1][0] ~^ image[24][20])} + {7'd0,(kernel[1][1] ~^ image[24][21])} + {7'd0,(kernel[1][2] ~^ image[24][22])} + {7'd0,(kernel[1][3] ~^ image[24][23])} + {7'd0,(kernel[1][4] ~^ image[24][24])} + {7'd0,(kernel[2][0] ~^ image[25][20])} + {7'd0,(kernel[2][1] ~^ image[25][21])} + {7'd0,(kernel[2][2] ~^ image[25][22])} + {7'd0,(kernel[2][3] ~^ image[25][23])} + {7'd0,(kernel[2][4] ~^ image[25][24])} + {7'd0,(kernel[3][0] ~^ image[26][20])} + {7'd0,(kernel[3][1] ~^ image[26][21])} + {7'd0,(kernel[3][2] ~^ image[26][22])} + {7'd0,(kernel[3][3] ~^ image[26][23])} + {7'd0,(kernel[3][4] ~^ image[26][24])} + {7'd0,(kernel[4][0] ~^ image[27][20])} + {7'd0,(kernel[4][1] ~^ image[27][21])} + {7'd0,(kernel[4][2] ~^ image[27][22])} + {7'd0,(kernel[4][3] ~^ image[27][23])} + {7'd0,(kernel[4][4] ~^ image[27][24])};
assign out_fmap[23][21][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[23][21])} + {7'd0,(kernel[0][1] ~^ image[23][22])} + {7'd0,(kernel[0][2] ~^ image[23][23])} + {7'd0,(kernel[0][3] ~^ image[23][24])} + {7'd0,(kernel[0][4] ~^ image[23][25])} + {7'd0,(kernel[1][0] ~^ image[24][21])} + {7'd0,(kernel[1][1] ~^ image[24][22])} + {7'd0,(kernel[1][2] ~^ image[24][23])} + {7'd0,(kernel[1][3] ~^ image[24][24])} + {7'd0,(kernel[1][4] ~^ image[24][25])} + {7'd0,(kernel[2][0] ~^ image[25][21])} + {7'd0,(kernel[2][1] ~^ image[25][22])} + {7'd0,(kernel[2][2] ~^ image[25][23])} + {7'd0,(kernel[2][3] ~^ image[25][24])} + {7'd0,(kernel[2][4] ~^ image[25][25])} + {7'd0,(kernel[3][0] ~^ image[26][21])} + {7'd0,(kernel[3][1] ~^ image[26][22])} + {7'd0,(kernel[3][2] ~^ image[26][23])} + {7'd0,(kernel[3][3] ~^ image[26][24])} + {7'd0,(kernel[3][4] ~^ image[26][25])} + {7'd0,(kernel[4][0] ~^ image[27][21])} + {7'd0,(kernel[4][1] ~^ image[27][22])} + {7'd0,(kernel[4][2] ~^ image[27][23])} + {7'd0,(kernel[4][3] ~^ image[27][24])} + {7'd0,(kernel[4][4] ~^ image[27][25])};
assign out_fmap[23][22][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[23][22])} + {7'd0,(kernel[0][1] ~^ image[23][23])} + {7'd0,(kernel[0][2] ~^ image[23][24])} + {7'd0,(kernel[0][3] ~^ image[23][25])} + {7'd0,(kernel[0][4] ~^ image[23][26])} + {7'd0,(kernel[1][0] ~^ image[24][22])} + {7'd0,(kernel[1][1] ~^ image[24][23])} + {7'd0,(kernel[1][2] ~^ image[24][24])} + {7'd0,(kernel[1][3] ~^ image[24][25])} + {7'd0,(kernel[1][4] ~^ image[24][26])} + {7'd0,(kernel[2][0] ~^ image[25][22])} + {7'd0,(kernel[2][1] ~^ image[25][23])} + {7'd0,(kernel[2][2] ~^ image[25][24])} + {7'd0,(kernel[2][3] ~^ image[25][25])} + {7'd0,(kernel[2][4] ~^ image[25][26])} + {7'd0,(kernel[3][0] ~^ image[26][22])} + {7'd0,(kernel[3][1] ~^ image[26][23])} + {7'd0,(kernel[3][2] ~^ image[26][24])} + {7'd0,(kernel[3][3] ~^ image[26][25])} + {7'd0,(kernel[3][4] ~^ image[26][26])} + {7'd0,(kernel[4][0] ~^ image[27][22])} + {7'd0,(kernel[4][1] ~^ image[27][23])} + {7'd0,(kernel[4][2] ~^ image[27][24])} + {7'd0,(kernel[4][3] ~^ image[27][25])} + {7'd0,(kernel[4][4] ~^ image[27][26])};
assign out_fmap[23][23][bW-1:0] = {7'd0,(kernel[0][0] ~^ image[23][23])} + {7'd0,(kernel[0][1] ~^ image[23][24])} + {7'd0,(kernel[0][2] ~^ image[23][25])} + {7'd0,(kernel[0][3] ~^ image[23][26])} + {7'd0,(kernel[0][4] ~^ image[23][27])} + {7'd0,(kernel[1][0] ~^ image[24][23])} + {7'd0,(kernel[1][1] ~^ image[24][24])} + {7'd0,(kernel[1][2] ~^ image[24][25])} + {7'd0,(kernel[1][3] ~^ image[24][26])} + {7'd0,(kernel[1][4] ~^ image[24][27])} + {7'd0,(kernel[2][0] ~^ image[25][23])} + {7'd0,(kernel[2][1] ~^ image[25][24])} + {7'd0,(kernel[2][2] ~^ image[25][25])} + {7'd0,(kernel[2][3] ~^ image[25][26])} + {7'd0,(kernel[2][4] ~^ image[25][27])} + {7'd0,(kernel[3][0] ~^ image[26][23])} + {7'd0,(kernel[3][1] ~^ image[26][24])} + {7'd0,(kernel[3][2] ~^ image[26][25])} + {7'd0,(kernel[3][3] ~^ image[26][26])} + {7'd0,(kernel[3][4] ~^ image[26][27])} + {7'd0,(kernel[4][0] ~^ image[27][23])} + {7'd0,(kernel[4][1] ~^ image[27][24])} + {7'd0,(kernel[4][2] ~^ image[27][25])} + {7'd0,(kernel[4][3] ~^ image[27][26])} + {7'd0,(kernel[4][4] ~^ image[27][27])};

endmodule