module conv2
    #( parameter bW = 8 )
    (
    input  logic [0:18*12*12 -1]      image         ,
    input  logic [0:18*60*5*5-1]      kernels       ,
    output logic [0:18*60*8*8*bW-1] xor_out 
    );

convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[1*5*5:2*5*5-1]), .o_out_fmap(xor_out[1*8*8*bW:2*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[2*5*5:3*5*5-1]), .o_out_fmap(xor_out[2*8*8*bW:3*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[3*5*5:4*5*5-1]), .o_out_fmap(xor_out[3*8*8*bW:4*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[4*5*5:5*5*5-1]), .o_out_fmap(xor_out[4*8*8*bW:5*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[5*5*5:6*5*5-1]), .o_out_fmap(xor_out[5*8*8*bW:6*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[6*5*5:7*5*5-1]), .o_out_fmap(xor_out[6*8*8*bW:7*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[7*5*5:8*5*5-1]), .o_out_fmap(xor_out[7*8*8*bW:8*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[8*5*5:9*5*5-1]), .o_out_fmap(xor_out[8*8*8*bW:9*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[9*5*5:10*5*5-1]), .o_out_fmap(xor_out[9*8*8*bW:10*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[10*5*5:11*5*5-1]), .o_out_fmap(xor_out[10*8*8*bW:11*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[11*5*5:12*5*5-1]), .o_out_fmap(xor_out[11*8*8*bW:12*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[12*5*5:13*5*5-1]), .o_out_fmap(xor_out[12*8*8*bW:13*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[13*5*5:14*5*5-1]), .o_out_fmap(xor_out[13*8*8*bW:14*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[14*5*5:15*5*5-1]), .o_out_fmap(xor_out[14*8*8*bW:15*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[15*5*5:16*5*5-1]), .o_out_fmap(xor_out[15*8*8*bW:16*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[16*5*5:17*5*5-1]), .o_out_fmap(xor_out[16*8*8*bW:17*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[17*5*5:18*5*5-1]), .o_out_fmap(xor_out[17*8*8*bW:18*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[18*5*5:19*5*5-1]), .o_out_fmap(xor_out[18*8*8*bW:19*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[19*5*5:20*5*5-1]), .o_out_fmap(xor_out[19*8*8*bW:20*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[20*5*5:21*5*5-1]), .o_out_fmap(xor_out[20*8*8*bW:21*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[21*5*5:22*5*5-1]), .o_out_fmap(xor_out[21*8*8*bW:22*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[22*5*5:23*5*5-1]), .o_out_fmap(xor_out[22*8*8*bW:23*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[23*5*5:24*5*5-1]), .o_out_fmap(xor_out[23*8*8*bW:24*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[24*5*5:25*5*5-1]), .o_out_fmap(xor_out[24*8*8*bW:25*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[25*5*5:26*5*5-1]), .o_out_fmap(xor_out[25*8*8*bW:26*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[26*5*5:27*5*5-1]), .o_out_fmap(xor_out[26*8*8*bW:27*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[27*5*5:28*5*5-1]), .o_out_fmap(xor_out[27*8*8*bW:28*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[28*5*5:29*5*5-1]), .o_out_fmap(xor_out[28*8*8*bW:29*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[29*5*5:30*5*5-1]), .o_out_fmap(xor_out[29*8*8*bW:30*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[30*5*5:31*5*5-1]), .o_out_fmap(xor_out[30*8*8*bW:31*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[31*5*5:32*5*5-1]), .o_out_fmap(xor_out[31*8*8*bW:32*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[32*5*5:33*5*5-1]), .o_out_fmap(xor_out[32*8*8*bW:33*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[33*5*5:34*5*5-1]), .o_out_fmap(xor_out[33*8*8*bW:34*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[34*5*5:35*5*5-1]), .o_out_fmap(xor_out[34*8*8*bW:35*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[35*5*5:36*5*5-1]), .o_out_fmap(xor_out[35*8*8*bW:36*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[36*5*5:37*5*5-1]), .o_out_fmap(xor_out[36*8*8*bW:37*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[37*5*5:38*5*5-1]), .o_out_fmap(xor_out[37*8*8*bW:38*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[38*5*5:39*5*5-1]), .o_out_fmap(xor_out[38*8*8*bW:39*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[39*5*5:40*5*5-1]), .o_out_fmap(xor_out[39*8*8*bW:40*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[40*5*5:41*5*5-1]), .o_out_fmap(xor_out[40*8*8*bW:41*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[41*5*5:42*5*5-1]), .o_out_fmap(xor_out[41*8*8*bW:42*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[42*5*5:43*5*5-1]), .o_out_fmap(xor_out[42*8*8*bW:43*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[43*5*5:44*5*5-1]), .o_out_fmap(xor_out[43*8*8*bW:44*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[44*5*5:45*5*5-1]), .o_out_fmap(xor_out[44*8*8*bW:45*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[45*5*5:46*5*5-1]), .o_out_fmap(xor_out[45*8*8*bW:46*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[46*5*5:47*5*5-1]), .o_out_fmap(xor_out[46*8*8*bW:47*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[47*5*5:48*5*5-1]), .o_out_fmap(xor_out[47*8*8*bW:48*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[48*5*5:49*5*5-1]), .o_out_fmap(xor_out[48*8*8*bW:49*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[49*5*5:50*5*5-1]), .o_out_fmap(xor_out[49*8*8*bW:50*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[50*5*5:51*5*5-1]), .o_out_fmap(xor_out[50*8*8*bW:51*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[51*5*5:52*5*5-1]), .o_out_fmap(xor_out[51*8*8*bW:52*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[52*5*5:53*5*5-1]), .o_out_fmap(xor_out[52*8*8*bW:53*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[53*5*5:54*5*5-1]), .o_out_fmap(xor_out[53*8*8*bW:54*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[54*5*5:55*5*5-1]), .o_out_fmap(xor_out[54*8*8*bW:55*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[55*5*5:56*5*5-1]), .o_out_fmap(xor_out[55*8*8*bW:56*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[56*5*5:57*5*5-1]), .o_out_fmap(xor_out[56*8*8*bW:57*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[57*5*5:58*5*5-1]), .o_out_fmap(xor_out[57*8*8*bW:58*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[58*5*5:59*5*5-1]), .o_out_fmap(xor_out[58*8*8*bW:59*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[59*5*5:60*5*5-1]), .o_out_fmap(xor_out[59*8*8*bW:60*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[2*5*5:3*5*5-1]), .o_out_fmap(xor_out[2*8*8*bW:3*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[4*5*5:5*5*5-1]), .o_out_fmap(xor_out[4*8*8*bW:5*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[6*5*5:7*5*5-1]), .o_out_fmap(xor_out[6*8*8*bW:7*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[8*5*5:9*5*5-1]), .o_out_fmap(xor_out[8*8*8*bW:9*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[10*5*5:11*5*5-1]), .o_out_fmap(xor_out[10*8*8*bW:11*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[12*5*5:13*5*5-1]), .o_out_fmap(xor_out[12*8*8*bW:13*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[14*5*5:15*5*5-1]), .o_out_fmap(xor_out[14*8*8*bW:15*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[16*5*5:17*5*5-1]), .o_out_fmap(xor_out[16*8*8*bW:17*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[18*5*5:19*5*5-1]), .o_out_fmap(xor_out[18*8*8*bW:19*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[20*5*5:21*5*5-1]), .o_out_fmap(xor_out[20*8*8*bW:21*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[22*5*5:23*5*5-1]), .o_out_fmap(xor_out[22*8*8*bW:23*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[24*5*5:25*5*5-1]), .o_out_fmap(xor_out[24*8*8*bW:25*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[26*5*5:27*5*5-1]), .o_out_fmap(xor_out[26*8*8*bW:27*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[28*5*5:29*5*5-1]), .o_out_fmap(xor_out[28*8*8*bW:29*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[30*5*5:31*5*5-1]), .o_out_fmap(xor_out[30*8*8*bW:31*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[32*5*5:33*5*5-1]), .o_out_fmap(xor_out[32*8*8*bW:33*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[34*5*5:35*5*5-1]), .o_out_fmap(xor_out[34*8*8*bW:35*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[36*5*5:37*5*5-1]), .o_out_fmap(xor_out[36*8*8*bW:37*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[38*5*5:39*5*5-1]), .o_out_fmap(xor_out[38*8*8*bW:39*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[40*5*5:41*5*5-1]), .o_out_fmap(xor_out[40*8*8*bW:41*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[42*5*5:43*5*5-1]), .o_out_fmap(xor_out[42*8*8*bW:43*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[44*5*5:45*5*5-1]), .o_out_fmap(xor_out[44*8*8*bW:45*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[46*5*5:47*5*5-1]), .o_out_fmap(xor_out[46*8*8*bW:47*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[48*5*5:49*5*5-1]), .o_out_fmap(xor_out[48*8*8*bW:49*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[50*5*5:51*5*5-1]), .o_out_fmap(xor_out[50*8*8*bW:51*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[52*5*5:53*5*5-1]), .o_out_fmap(xor_out[52*8*8*bW:53*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[54*5*5:55*5*5-1]), .o_out_fmap(xor_out[54*8*8*bW:55*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[56*5*5:57*5*5-1]), .o_out_fmap(xor_out[56*8*8*bW:57*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[58*5*5:59*5*5-1]), .o_out_fmap(xor_out[58*8*8*bW:59*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[60*5*5:61*5*5-1]), .o_out_fmap(xor_out[60*8*8*bW:61*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[62*5*5:63*5*5-1]), .o_out_fmap(xor_out[62*8*8*bW:63*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[64*5*5:65*5*5-1]), .o_out_fmap(xor_out[64*8*8*bW:65*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[66*5*5:67*5*5-1]), .o_out_fmap(xor_out[66*8*8*bW:67*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[68*5*5:69*5*5-1]), .o_out_fmap(xor_out[68*8*8*bW:69*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[70*5*5:71*5*5-1]), .o_out_fmap(xor_out[70*8*8*bW:71*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[72*5*5:73*5*5-1]), .o_out_fmap(xor_out[72*8*8*bW:73*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[74*5*5:75*5*5-1]), .o_out_fmap(xor_out[74*8*8*bW:75*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[76*5*5:77*5*5-1]), .o_out_fmap(xor_out[76*8*8*bW:77*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[78*5*5:79*5*5-1]), .o_out_fmap(xor_out[78*8*8*bW:79*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[80*5*5:81*5*5-1]), .o_out_fmap(xor_out[80*8*8*bW:81*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[82*5*5:83*5*5-1]), .o_out_fmap(xor_out[82*8*8*bW:83*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[84*5*5:85*5*5-1]), .o_out_fmap(xor_out[84*8*8*bW:85*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[86*5*5:87*5*5-1]), .o_out_fmap(xor_out[86*8*8*bW:87*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[88*5*5:89*5*5-1]), .o_out_fmap(xor_out[88*8*8*bW:89*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[90*5*5:91*5*5-1]), .o_out_fmap(xor_out[90*8*8*bW:91*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[92*5*5:93*5*5-1]), .o_out_fmap(xor_out[92*8*8*bW:93*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[94*5*5:95*5*5-1]), .o_out_fmap(xor_out[94*8*8*bW:95*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[96*5*5:97*5*5-1]), .o_out_fmap(xor_out[96*8*8*bW:97*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[98*5*5:99*5*5-1]), .o_out_fmap(xor_out[98*8*8*bW:99*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[100*5*5:101*5*5-1]), .o_out_fmap(xor_out[100*8*8*bW:101*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[102*5*5:103*5*5-1]), .o_out_fmap(xor_out[102*8*8*bW:103*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[104*5*5:105*5*5-1]), .o_out_fmap(xor_out[104*8*8*bW:105*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[106*5*5:107*5*5-1]), .o_out_fmap(xor_out[106*8*8*bW:107*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[108*5*5:109*5*5-1]), .o_out_fmap(xor_out[108*8*8*bW:109*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[110*5*5:111*5*5-1]), .o_out_fmap(xor_out[110*8*8*bW:111*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[112*5*5:113*5*5-1]), .o_out_fmap(xor_out[112*8*8*bW:113*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[114*5*5:115*5*5-1]), .o_out_fmap(xor_out[114*8*8*bW:115*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[116*5*5:117*5*5-1]), .o_out_fmap(xor_out[116*8*8*bW:117*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[118*5*5:119*5*5-1]), .o_out_fmap(xor_out[118*8*8*bW:119*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[3*5*5:4*5*5-1]), .o_out_fmap(xor_out[3*8*8*bW:4*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[6*5*5:7*5*5-1]), .o_out_fmap(xor_out[6*8*8*bW:7*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[9*5*5:10*5*5-1]), .o_out_fmap(xor_out[9*8*8*bW:10*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[12*5*5:13*5*5-1]), .o_out_fmap(xor_out[12*8*8*bW:13*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[15*5*5:16*5*5-1]), .o_out_fmap(xor_out[15*8*8*bW:16*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[18*5*5:19*5*5-1]), .o_out_fmap(xor_out[18*8*8*bW:19*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[21*5*5:22*5*5-1]), .o_out_fmap(xor_out[21*8*8*bW:22*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[24*5*5:25*5*5-1]), .o_out_fmap(xor_out[24*8*8*bW:25*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[27*5*5:28*5*5-1]), .o_out_fmap(xor_out[27*8*8*bW:28*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[30*5*5:31*5*5-1]), .o_out_fmap(xor_out[30*8*8*bW:31*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[33*5*5:34*5*5-1]), .o_out_fmap(xor_out[33*8*8*bW:34*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[36*5*5:37*5*5-1]), .o_out_fmap(xor_out[36*8*8*bW:37*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[39*5*5:40*5*5-1]), .o_out_fmap(xor_out[39*8*8*bW:40*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[42*5*5:43*5*5-1]), .o_out_fmap(xor_out[42*8*8*bW:43*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[45*5*5:46*5*5-1]), .o_out_fmap(xor_out[45*8*8*bW:46*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[48*5*5:49*5*5-1]), .o_out_fmap(xor_out[48*8*8*bW:49*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[51*5*5:52*5*5-1]), .o_out_fmap(xor_out[51*8*8*bW:52*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[54*5*5:55*5*5-1]), .o_out_fmap(xor_out[54*8*8*bW:55*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[57*5*5:58*5*5-1]), .o_out_fmap(xor_out[57*8*8*bW:58*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[60*5*5:61*5*5-1]), .o_out_fmap(xor_out[60*8*8*bW:61*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[63*5*5:64*5*5-1]), .o_out_fmap(xor_out[63*8*8*bW:64*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[66*5*5:67*5*5-1]), .o_out_fmap(xor_out[66*8*8*bW:67*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[69*5*5:70*5*5-1]), .o_out_fmap(xor_out[69*8*8*bW:70*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[72*5*5:73*5*5-1]), .o_out_fmap(xor_out[72*8*8*bW:73*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[75*5*5:76*5*5-1]), .o_out_fmap(xor_out[75*8*8*bW:76*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[78*5*5:79*5*5-1]), .o_out_fmap(xor_out[78*8*8*bW:79*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[81*5*5:82*5*5-1]), .o_out_fmap(xor_out[81*8*8*bW:82*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[84*5*5:85*5*5-1]), .o_out_fmap(xor_out[84*8*8*bW:85*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[87*5*5:88*5*5-1]), .o_out_fmap(xor_out[87*8*8*bW:88*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[90*5*5:91*5*5-1]), .o_out_fmap(xor_out[90*8*8*bW:91*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[93*5*5:94*5*5-1]), .o_out_fmap(xor_out[93*8*8*bW:94*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[96*5*5:97*5*5-1]), .o_out_fmap(xor_out[96*8*8*bW:97*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[99*5*5:100*5*5-1]), .o_out_fmap(xor_out[99*8*8*bW:100*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[102*5*5:103*5*5-1]), .o_out_fmap(xor_out[102*8*8*bW:103*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[105*5*5:106*5*5-1]), .o_out_fmap(xor_out[105*8*8*bW:106*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[108*5*5:109*5*5-1]), .o_out_fmap(xor_out[108*8*8*bW:109*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[111*5*5:112*5*5-1]), .o_out_fmap(xor_out[111*8*8*bW:112*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[114*5*5:115*5*5-1]), .o_out_fmap(xor_out[114*8*8*bW:115*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[117*5*5:118*5*5-1]), .o_out_fmap(xor_out[117*8*8*bW:118*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[120*5*5:121*5*5-1]), .o_out_fmap(xor_out[120*8*8*bW:121*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[123*5*5:124*5*5-1]), .o_out_fmap(xor_out[123*8*8*bW:124*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[126*5*5:127*5*5-1]), .o_out_fmap(xor_out[126*8*8*bW:127*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[129*5*5:130*5*5-1]), .o_out_fmap(xor_out[129*8*8*bW:130*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[132*5*5:133*5*5-1]), .o_out_fmap(xor_out[132*8*8*bW:133*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[135*5*5:136*5*5-1]), .o_out_fmap(xor_out[135*8*8*bW:136*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[138*5*5:139*5*5-1]), .o_out_fmap(xor_out[138*8*8*bW:139*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[141*5*5:142*5*5-1]), .o_out_fmap(xor_out[141*8*8*bW:142*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[144*5*5:145*5*5-1]), .o_out_fmap(xor_out[144*8*8*bW:145*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[147*5*5:148*5*5-1]), .o_out_fmap(xor_out[147*8*8*bW:148*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[150*5*5:151*5*5-1]), .o_out_fmap(xor_out[150*8*8*bW:151*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[153*5*5:154*5*5-1]), .o_out_fmap(xor_out[153*8*8*bW:154*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[156*5*5:157*5*5-1]), .o_out_fmap(xor_out[156*8*8*bW:157*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[159*5*5:160*5*5-1]), .o_out_fmap(xor_out[159*8*8*bW:160*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[162*5*5:163*5*5-1]), .o_out_fmap(xor_out[162*8*8*bW:163*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[165*5*5:166*5*5-1]), .o_out_fmap(xor_out[165*8*8*bW:166*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[168*5*5:169*5*5-1]), .o_out_fmap(xor_out[168*8*8*bW:169*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[171*5*5:172*5*5-1]), .o_out_fmap(xor_out[171*8*8*bW:172*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[174*5*5:175*5*5-1]), .o_out_fmap(xor_out[174*8*8*bW:175*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[177*5*5:178*5*5-1]), .o_out_fmap(xor_out[177*8*8*bW:178*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[4*5*5:5*5*5-1]), .o_out_fmap(xor_out[4*8*8*bW:5*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[8*5*5:9*5*5-1]), .o_out_fmap(xor_out[8*8*8*bW:9*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[12*5*5:13*5*5-1]), .o_out_fmap(xor_out[12*8*8*bW:13*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[16*5*5:17*5*5-1]), .o_out_fmap(xor_out[16*8*8*bW:17*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[20*5*5:21*5*5-1]), .o_out_fmap(xor_out[20*8*8*bW:21*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[24*5*5:25*5*5-1]), .o_out_fmap(xor_out[24*8*8*bW:25*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[28*5*5:29*5*5-1]), .o_out_fmap(xor_out[28*8*8*bW:29*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[32*5*5:33*5*5-1]), .o_out_fmap(xor_out[32*8*8*bW:33*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[36*5*5:37*5*5-1]), .o_out_fmap(xor_out[36*8*8*bW:37*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[40*5*5:41*5*5-1]), .o_out_fmap(xor_out[40*8*8*bW:41*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[44*5*5:45*5*5-1]), .o_out_fmap(xor_out[44*8*8*bW:45*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[48*5*5:49*5*5-1]), .o_out_fmap(xor_out[48*8*8*bW:49*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[52*5*5:53*5*5-1]), .o_out_fmap(xor_out[52*8*8*bW:53*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[56*5*5:57*5*5-1]), .o_out_fmap(xor_out[56*8*8*bW:57*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[60*5*5:61*5*5-1]), .o_out_fmap(xor_out[60*8*8*bW:61*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[64*5*5:65*5*5-1]), .o_out_fmap(xor_out[64*8*8*bW:65*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[68*5*5:69*5*5-1]), .o_out_fmap(xor_out[68*8*8*bW:69*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[72*5*5:73*5*5-1]), .o_out_fmap(xor_out[72*8*8*bW:73*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[76*5*5:77*5*5-1]), .o_out_fmap(xor_out[76*8*8*bW:77*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[80*5*5:81*5*5-1]), .o_out_fmap(xor_out[80*8*8*bW:81*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[84*5*5:85*5*5-1]), .o_out_fmap(xor_out[84*8*8*bW:85*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[88*5*5:89*5*5-1]), .o_out_fmap(xor_out[88*8*8*bW:89*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[92*5*5:93*5*5-1]), .o_out_fmap(xor_out[92*8*8*bW:93*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[96*5*5:97*5*5-1]), .o_out_fmap(xor_out[96*8*8*bW:97*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[100*5*5:101*5*5-1]), .o_out_fmap(xor_out[100*8*8*bW:101*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[104*5*5:105*5*5-1]), .o_out_fmap(xor_out[104*8*8*bW:105*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[108*5*5:109*5*5-1]), .o_out_fmap(xor_out[108*8*8*bW:109*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[112*5*5:113*5*5-1]), .o_out_fmap(xor_out[112*8*8*bW:113*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[116*5*5:117*5*5-1]), .o_out_fmap(xor_out[116*8*8*bW:117*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[120*5*5:121*5*5-1]), .o_out_fmap(xor_out[120*8*8*bW:121*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[124*5*5:125*5*5-1]), .o_out_fmap(xor_out[124*8*8*bW:125*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[128*5*5:129*5*5-1]), .o_out_fmap(xor_out[128*8*8*bW:129*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[132*5*5:133*5*5-1]), .o_out_fmap(xor_out[132*8*8*bW:133*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[136*5*5:137*5*5-1]), .o_out_fmap(xor_out[136*8*8*bW:137*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[140*5*5:141*5*5-1]), .o_out_fmap(xor_out[140*8*8*bW:141*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[144*5*5:145*5*5-1]), .o_out_fmap(xor_out[144*8*8*bW:145*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[148*5*5:149*5*5-1]), .o_out_fmap(xor_out[148*8*8*bW:149*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[152*5*5:153*5*5-1]), .o_out_fmap(xor_out[152*8*8*bW:153*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[156*5*5:157*5*5-1]), .o_out_fmap(xor_out[156*8*8*bW:157*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[160*5*5:161*5*5-1]), .o_out_fmap(xor_out[160*8*8*bW:161*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[164*5*5:165*5*5-1]), .o_out_fmap(xor_out[164*8*8*bW:165*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[168*5*5:169*5*5-1]), .o_out_fmap(xor_out[168*8*8*bW:169*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[172*5*5:173*5*5-1]), .o_out_fmap(xor_out[172*8*8*bW:173*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[176*5*5:177*5*5-1]), .o_out_fmap(xor_out[176*8*8*bW:177*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[180*5*5:181*5*5-1]), .o_out_fmap(xor_out[180*8*8*bW:181*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[184*5*5:185*5*5-1]), .o_out_fmap(xor_out[184*8*8*bW:185*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[188*5*5:189*5*5-1]), .o_out_fmap(xor_out[188*8*8*bW:189*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[192*5*5:193*5*5-1]), .o_out_fmap(xor_out[192*8*8*bW:193*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[196*5*5:197*5*5-1]), .o_out_fmap(xor_out[196*8*8*bW:197*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[200*5*5:201*5*5-1]), .o_out_fmap(xor_out[200*8*8*bW:201*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[204*5*5:205*5*5-1]), .o_out_fmap(xor_out[204*8*8*bW:205*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[208*5*5:209*5*5-1]), .o_out_fmap(xor_out[208*8*8*bW:209*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[212*5*5:213*5*5-1]), .o_out_fmap(xor_out[212*8*8*bW:213*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[216*5*5:217*5*5-1]), .o_out_fmap(xor_out[216*8*8*bW:217*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[220*5*5:221*5*5-1]), .o_out_fmap(xor_out[220*8*8*bW:221*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[224*5*5:225*5*5-1]), .o_out_fmap(xor_out[224*8*8*bW:225*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[228*5*5:229*5*5-1]), .o_out_fmap(xor_out[228*8*8*bW:229*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[232*5*5:233*5*5-1]), .o_out_fmap(xor_out[232*8*8*bW:233*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[236*5*5:237*5*5-1]), .o_out_fmap(xor_out[236*8*8*bW:237*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[5*5*5:6*5*5-1]), .o_out_fmap(xor_out[5*8*8*bW:6*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[10*5*5:11*5*5-1]), .o_out_fmap(xor_out[10*8*8*bW:11*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[15*5*5:16*5*5-1]), .o_out_fmap(xor_out[15*8*8*bW:16*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[20*5*5:21*5*5-1]), .o_out_fmap(xor_out[20*8*8*bW:21*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[25*5*5:26*5*5-1]), .o_out_fmap(xor_out[25*8*8*bW:26*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[30*5*5:31*5*5-1]), .o_out_fmap(xor_out[30*8*8*bW:31*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[35*5*5:36*5*5-1]), .o_out_fmap(xor_out[35*8*8*bW:36*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[40*5*5:41*5*5-1]), .o_out_fmap(xor_out[40*8*8*bW:41*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[45*5*5:46*5*5-1]), .o_out_fmap(xor_out[45*8*8*bW:46*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[50*5*5:51*5*5-1]), .o_out_fmap(xor_out[50*8*8*bW:51*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[55*5*5:56*5*5-1]), .o_out_fmap(xor_out[55*8*8*bW:56*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[60*5*5:61*5*5-1]), .o_out_fmap(xor_out[60*8*8*bW:61*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[65*5*5:66*5*5-1]), .o_out_fmap(xor_out[65*8*8*bW:66*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[70*5*5:71*5*5-1]), .o_out_fmap(xor_out[70*8*8*bW:71*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[75*5*5:76*5*5-1]), .o_out_fmap(xor_out[75*8*8*bW:76*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[80*5*5:81*5*5-1]), .o_out_fmap(xor_out[80*8*8*bW:81*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[85*5*5:86*5*5-1]), .o_out_fmap(xor_out[85*8*8*bW:86*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[90*5*5:91*5*5-1]), .o_out_fmap(xor_out[90*8*8*bW:91*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[95*5*5:96*5*5-1]), .o_out_fmap(xor_out[95*8*8*bW:96*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[100*5*5:101*5*5-1]), .o_out_fmap(xor_out[100*8*8*bW:101*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[105*5*5:106*5*5-1]), .o_out_fmap(xor_out[105*8*8*bW:106*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[110*5*5:111*5*5-1]), .o_out_fmap(xor_out[110*8*8*bW:111*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[115*5*5:116*5*5-1]), .o_out_fmap(xor_out[115*8*8*bW:116*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[120*5*5:121*5*5-1]), .o_out_fmap(xor_out[120*8*8*bW:121*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[125*5*5:126*5*5-1]), .o_out_fmap(xor_out[125*8*8*bW:126*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[130*5*5:131*5*5-1]), .o_out_fmap(xor_out[130*8*8*bW:131*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[135*5*5:136*5*5-1]), .o_out_fmap(xor_out[135*8*8*bW:136*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[140*5*5:141*5*5-1]), .o_out_fmap(xor_out[140*8*8*bW:141*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[145*5*5:146*5*5-1]), .o_out_fmap(xor_out[145*8*8*bW:146*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[150*5*5:151*5*5-1]), .o_out_fmap(xor_out[150*8*8*bW:151*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[155*5*5:156*5*5-1]), .o_out_fmap(xor_out[155*8*8*bW:156*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[160*5*5:161*5*5-1]), .o_out_fmap(xor_out[160*8*8*bW:161*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[165*5*5:166*5*5-1]), .o_out_fmap(xor_out[165*8*8*bW:166*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[170*5*5:171*5*5-1]), .o_out_fmap(xor_out[170*8*8*bW:171*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[175*5*5:176*5*5-1]), .o_out_fmap(xor_out[175*8*8*bW:176*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[180*5*5:181*5*5-1]), .o_out_fmap(xor_out[180*8*8*bW:181*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[185*5*5:186*5*5-1]), .o_out_fmap(xor_out[185*8*8*bW:186*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[190*5*5:191*5*5-1]), .o_out_fmap(xor_out[190*8*8*bW:191*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[195*5*5:196*5*5-1]), .o_out_fmap(xor_out[195*8*8*bW:196*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[200*5*5:201*5*5-1]), .o_out_fmap(xor_out[200*8*8*bW:201*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[205*5*5:206*5*5-1]), .o_out_fmap(xor_out[205*8*8*bW:206*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[210*5*5:211*5*5-1]), .o_out_fmap(xor_out[210*8*8*bW:211*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[215*5*5:216*5*5-1]), .o_out_fmap(xor_out[215*8*8*bW:216*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[220*5*5:221*5*5-1]), .o_out_fmap(xor_out[220*8*8*bW:221*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[225*5*5:226*5*5-1]), .o_out_fmap(xor_out[225*8*8*bW:226*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[230*5*5:231*5*5-1]), .o_out_fmap(xor_out[230*8*8*bW:231*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[235*5*5:236*5*5-1]), .o_out_fmap(xor_out[235*8*8*bW:236*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[240*5*5:241*5*5-1]), .o_out_fmap(xor_out[240*8*8*bW:241*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[245*5*5:246*5*5-1]), .o_out_fmap(xor_out[245*8*8*bW:246*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[250*5*5:251*5*5-1]), .o_out_fmap(xor_out[250*8*8*bW:251*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[255*5*5:256*5*5-1]), .o_out_fmap(xor_out[255*8*8*bW:256*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[260*5*5:261*5*5-1]), .o_out_fmap(xor_out[260*8*8*bW:261*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[265*5*5:266*5*5-1]), .o_out_fmap(xor_out[265*8*8*bW:266*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[270*5*5:271*5*5-1]), .o_out_fmap(xor_out[270*8*8*bW:271*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[275*5*5:276*5*5-1]), .o_out_fmap(xor_out[275*8*8*bW:276*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[280*5*5:281*5*5-1]), .o_out_fmap(xor_out[280*8*8*bW:281*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[285*5*5:286*5*5-1]), .o_out_fmap(xor_out[285*8*8*bW:286*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[290*5*5:291*5*5-1]), .o_out_fmap(xor_out[290*8*8*bW:291*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[295*5*5:296*5*5-1]), .o_out_fmap(xor_out[295*8*8*bW:296*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[6*5*5:7*5*5-1]), .o_out_fmap(xor_out[6*8*8*bW:7*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[12*5*5:13*5*5-1]), .o_out_fmap(xor_out[12*8*8*bW:13*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[18*5*5:19*5*5-1]), .o_out_fmap(xor_out[18*8*8*bW:19*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[24*5*5:25*5*5-1]), .o_out_fmap(xor_out[24*8*8*bW:25*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[30*5*5:31*5*5-1]), .o_out_fmap(xor_out[30*8*8*bW:31*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[36*5*5:37*5*5-1]), .o_out_fmap(xor_out[36*8*8*bW:37*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[42*5*5:43*5*5-1]), .o_out_fmap(xor_out[42*8*8*bW:43*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[48*5*5:49*5*5-1]), .o_out_fmap(xor_out[48*8*8*bW:49*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[54*5*5:55*5*5-1]), .o_out_fmap(xor_out[54*8*8*bW:55*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[60*5*5:61*5*5-1]), .o_out_fmap(xor_out[60*8*8*bW:61*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[66*5*5:67*5*5-1]), .o_out_fmap(xor_out[66*8*8*bW:67*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[72*5*5:73*5*5-1]), .o_out_fmap(xor_out[72*8*8*bW:73*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[78*5*5:79*5*5-1]), .o_out_fmap(xor_out[78*8*8*bW:79*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[84*5*5:85*5*5-1]), .o_out_fmap(xor_out[84*8*8*bW:85*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[90*5*5:91*5*5-1]), .o_out_fmap(xor_out[90*8*8*bW:91*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[96*5*5:97*5*5-1]), .o_out_fmap(xor_out[96*8*8*bW:97*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[102*5*5:103*5*5-1]), .o_out_fmap(xor_out[102*8*8*bW:103*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[108*5*5:109*5*5-1]), .o_out_fmap(xor_out[108*8*8*bW:109*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[114*5*5:115*5*5-1]), .o_out_fmap(xor_out[114*8*8*bW:115*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[120*5*5:121*5*5-1]), .o_out_fmap(xor_out[120*8*8*bW:121*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[126*5*5:127*5*5-1]), .o_out_fmap(xor_out[126*8*8*bW:127*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[132*5*5:133*5*5-1]), .o_out_fmap(xor_out[132*8*8*bW:133*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[138*5*5:139*5*5-1]), .o_out_fmap(xor_out[138*8*8*bW:139*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[144*5*5:145*5*5-1]), .o_out_fmap(xor_out[144*8*8*bW:145*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[150*5*5:151*5*5-1]), .o_out_fmap(xor_out[150*8*8*bW:151*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[156*5*5:157*5*5-1]), .o_out_fmap(xor_out[156*8*8*bW:157*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[162*5*5:163*5*5-1]), .o_out_fmap(xor_out[162*8*8*bW:163*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[168*5*5:169*5*5-1]), .o_out_fmap(xor_out[168*8*8*bW:169*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[174*5*5:175*5*5-1]), .o_out_fmap(xor_out[174*8*8*bW:175*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[180*5*5:181*5*5-1]), .o_out_fmap(xor_out[180*8*8*bW:181*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[186*5*5:187*5*5-1]), .o_out_fmap(xor_out[186*8*8*bW:187*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[192*5*5:193*5*5-1]), .o_out_fmap(xor_out[192*8*8*bW:193*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[198*5*5:199*5*5-1]), .o_out_fmap(xor_out[198*8*8*bW:199*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[204*5*5:205*5*5-1]), .o_out_fmap(xor_out[204*8*8*bW:205*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[210*5*5:211*5*5-1]), .o_out_fmap(xor_out[210*8*8*bW:211*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[216*5*5:217*5*5-1]), .o_out_fmap(xor_out[216*8*8*bW:217*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[222*5*5:223*5*5-1]), .o_out_fmap(xor_out[222*8*8*bW:223*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[228*5*5:229*5*5-1]), .o_out_fmap(xor_out[228*8*8*bW:229*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[234*5*5:235*5*5-1]), .o_out_fmap(xor_out[234*8*8*bW:235*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[240*5*5:241*5*5-1]), .o_out_fmap(xor_out[240*8*8*bW:241*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[246*5*5:247*5*5-1]), .o_out_fmap(xor_out[246*8*8*bW:247*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[252*5*5:253*5*5-1]), .o_out_fmap(xor_out[252*8*8*bW:253*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[258*5*5:259*5*5-1]), .o_out_fmap(xor_out[258*8*8*bW:259*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[264*5*5:265*5*5-1]), .o_out_fmap(xor_out[264*8*8*bW:265*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[270*5*5:271*5*5-1]), .o_out_fmap(xor_out[270*8*8*bW:271*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[276*5*5:277*5*5-1]), .o_out_fmap(xor_out[276*8*8*bW:277*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[282*5*5:283*5*5-1]), .o_out_fmap(xor_out[282*8*8*bW:283*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[288*5*5:289*5*5-1]), .o_out_fmap(xor_out[288*8*8*bW:289*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[294*5*5:295*5*5-1]), .o_out_fmap(xor_out[294*8*8*bW:295*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[300*5*5:301*5*5-1]), .o_out_fmap(xor_out[300*8*8*bW:301*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[306*5*5:307*5*5-1]), .o_out_fmap(xor_out[306*8*8*bW:307*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[312*5*5:313*5*5-1]), .o_out_fmap(xor_out[312*8*8*bW:313*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[318*5*5:319*5*5-1]), .o_out_fmap(xor_out[318*8*8*bW:319*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[324*5*5:325*5*5-1]), .o_out_fmap(xor_out[324*8*8*bW:325*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[330*5*5:331*5*5-1]), .o_out_fmap(xor_out[330*8*8*bW:331*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[336*5*5:337*5*5-1]), .o_out_fmap(xor_out[336*8*8*bW:337*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[342*5*5:343*5*5-1]), .o_out_fmap(xor_out[342*8*8*bW:343*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[348*5*5:349*5*5-1]), .o_out_fmap(xor_out[348*8*8*bW:349*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[354*5*5:355*5*5-1]), .o_out_fmap(xor_out[354*8*8*bW:355*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[7*5*5:8*5*5-1]), .o_out_fmap(xor_out[7*8*8*bW:8*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[14*5*5:15*5*5-1]), .o_out_fmap(xor_out[14*8*8*bW:15*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[21*5*5:22*5*5-1]), .o_out_fmap(xor_out[21*8*8*bW:22*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[28*5*5:29*5*5-1]), .o_out_fmap(xor_out[28*8*8*bW:29*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[35*5*5:36*5*5-1]), .o_out_fmap(xor_out[35*8*8*bW:36*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[42*5*5:43*5*5-1]), .o_out_fmap(xor_out[42*8*8*bW:43*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[49*5*5:50*5*5-1]), .o_out_fmap(xor_out[49*8*8*bW:50*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[56*5*5:57*5*5-1]), .o_out_fmap(xor_out[56*8*8*bW:57*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[63*5*5:64*5*5-1]), .o_out_fmap(xor_out[63*8*8*bW:64*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[70*5*5:71*5*5-1]), .o_out_fmap(xor_out[70*8*8*bW:71*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[77*5*5:78*5*5-1]), .o_out_fmap(xor_out[77*8*8*bW:78*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[84*5*5:85*5*5-1]), .o_out_fmap(xor_out[84*8*8*bW:85*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[91*5*5:92*5*5-1]), .o_out_fmap(xor_out[91*8*8*bW:92*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[98*5*5:99*5*5-1]), .o_out_fmap(xor_out[98*8*8*bW:99*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[105*5*5:106*5*5-1]), .o_out_fmap(xor_out[105*8*8*bW:106*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[112*5*5:113*5*5-1]), .o_out_fmap(xor_out[112*8*8*bW:113*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[119*5*5:120*5*5-1]), .o_out_fmap(xor_out[119*8*8*bW:120*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[126*5*5:127*5*5-1]), .o_out_fmap(xor_out[126*8*8*bW:127*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[133*5*5:134*5*5-1]), .o_out_fmap(xor_out[133*8*8*bW:134*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[140*5*5:141*5*5-1]), .o_out_fmap(xor_out[140*8*8*bW:141*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[147*5*5:148*5*5-1]), .o_out_fmap(xor_out[147*8*8*bW:148*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[154*5*5:155*5*5-1]), .o_out_fmap(xor_out[154*8*8*bW:155*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[161*5*5:162*5*5-1]), .o_out_fmap(xor_out[161*8*8*bW:162*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[168*5*5:169*5*5-1]), .o_out_fmap(xor_out[168*8*8*bW:169*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[175*5*5:176*5*5-1]), .o_out_fmap(xor_out[175*8*8*bW:176*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[182*5*5:183*5*5-1]), .o_out_fmap(xor_out[182*8*8*bW:183*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[189*5*5:190*5*5-1]), .o_out_fmap(xor_out[189*8*8*bW:190*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[196*5*5:197*5*5-1]), .o_out_fmap(xor_out[196*8*8*bW:197*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[203*5*5:204*5*5-1]), .o_out_fmap(xor_out[203*8*8*bW:204*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[210*5*5:211*5*5-1]), .o_out_fmap(xor_out[210*8*8*bW:211*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[217*5*5:218*5*5-1]), .o_out_fmap(xor_out[217*8*8*bW:218*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[224*5*5:225*5*5-1]), .o_out_fmap(xor_out[224*8*8*bW:225*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[231*5*5:232*5*5-1]), .o_out_fmap(xor_out[231*8*8*bW:232*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[238*5*5:239*5*5-1]), .o_out_fmap(xor_out[238*8*8*bW:239*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[245*5*5:246*5*5-1]), .o_out_fmap(xor_out[245*8*8*bW:246*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[252*5*5:253*5*5-1]), .o_out_fmap(xor_out[252*8*8*bW:253*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[259*5*5:260*5*5-1]), .o_out_fmap(xor_out[259*8*8*bW:260*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[266*5*5:267*5*5-1]), .o_out_fmap(xor_out[266*8*8*bW:267*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[273*5*5:274*5*5-1]), .o_out_fmap(xor_out[273*8*8*bW:274*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[280*5*5:281*5*5-1]), .o_out_fmap(xor_out[280*8*8*bW:281*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[287*5*5:288*5*5-1]), .o_out_fmap(xor_out[287*8*8*bW:288*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[294*5*5:295*5*5-1]), .o_out_fmap(xor_out[294*8*8*bW:295*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[301*5*5:302*5*5-1]), .o_out_fmap(xor_out[301*8*8*bW:302*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[308*5*5:309*5*5-1]), .o_out_fmap(xor_out[308*8*8*bW:309*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[315*5*5:316*5*5-1]), .o_out_fmap(xor_out[315*8*8*bW:316*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[322*5*5:323*5*5-1]), .o_out_fmap(xor_out[322*8*8*bW:323*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[329*5*5:330*5*5-1]), .o_out_fmap(xor_out[329*8*8*bW:330*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[336*5*5:337*5*5-1]), .o_out_fmap(xor_out[336*8*8*bW:337*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[343*5*5:344*5*5-1]), .o_out_fmap(xor_out[343*8*8*bW:344*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[350*5*5:351*5*5-1]), .o_out_fmap(xor_out[350*8*8*bW:351*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[357*5*5:358*5*5-1]), .o_out_fmap(xor_out[357*8*8*bW:358*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[364*5*5:365*5*5-1]), .o_out_fmap(xor_out[364*8*8*bW:365*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[371*5*5:372*5*5-1]), .o_out_fmap(xor_out[371*8*8*bW:372*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[378*5*5:379*5*5-1]), .o_out_fmap(xor_out[378*8*8*bW:379*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[385*5*5:386*5*5-1]), .o_out_fmap(xor_out[385*8*8*bW:386*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[392*5*5:393*5*5-1]), .o_out_fmap(xor_out[392*8*8*bW:393*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[399*5*5:400*5*5-1]), .o_out_fmap(xor_out[399*8*8*bW:400*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[406*5*5:407*5*5-1]), .o_out_fmap(xor_out[406*8*8*bW:407*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[413*5*5:414*5*5-1]), .o_out_fmap(xor_out[413*8*8*bW:414*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[8*5*5:9*5*5-1]), .o_out_fmap(xor_out[8*8*8*bW:9*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[16*5*5:17*5*5-1]), .o_out_fmap(xor_out[16*8*8*bW:17*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[24*5*5:25*5*5-1]), .o_out_fmap(xor_out[24*8*8*bW:25*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[32*5*5:33*5*5-1]), .o_out_fmap(xor_out[32*8*8*bW:33*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[40*5*5:41*5*5-1]), .o_out_fmap(xor_out[40*8*8*bW:41*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[48*5*5:49*5*5-1]), .o_out_fmap(xor_out[48*8*8*bW:49*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[56*5*5:57*5*5-1]), .o_out_fmap(xor_out[56*8*8*bW:57*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[64*5*5:65*5*5-1]), .o_out_fmap(xor_out[64*8*8*bW:65*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[72*5*5:73*5*5-1]), .o_out_fmap(xor_out[72*8*8*bW:73*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[80*5*5:81*5*5-1]), .o_out_fmap(xor_out[80*8*8*bW:81*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[88*5*5:89*5*5-1]), .o_out_fmap(xor_out[88*8*8*bW:89*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[96*5*5:97*5*5-1]), .o_out_fmap(xor_out[96*8*8*bW:97*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[104*5*5:105*5*5-1]), .o_out_fmap(xor_out[104*8*8*bW:105*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[112*5*5:113*5*5-1]), .o_out_fmap(xor_out[112*8*8*bW:113*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[120*5*5:121*5*5-1]), .o_out_fmap(xor_out[120*8*8*bW:121*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[128*5*5:129*5*5-1]), .o_out_fmap(xor_out[128*8*8*bW:129*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[136*5*5:137*5*5-1]), .o_out_fmap(xor_out[136*8*8*bW:137*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[144*5*5:145*5*5-1]), .o_out_fmap(xor_out[144*8*8*bW:145*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[152*5*5:153*5*5-1]), .o_out_fmap(xor_out[152*8*8*bW:153*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[160*5*5:161*5*5-1]), .o_out_fmap(xor_out[160*8*8*bW:161*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[168*5*5:169*5*5-1]), .o_out_fmap(xor_out[168*8*8*bW:169*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[176*5*5:177*5*5-1]), .o_out_fmap(xor_out[176*8*8*bW:177*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[184*5*5:185*5*5-1]), .o_out_fmap(xor_out[184*8*8*bW:185*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[192*5*5:193*5*5-1]), .o_out_fmap(xor_out[192*8*8*bW:193*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[200*5*5:201*5*5-1]), .o_out_fmap(xor_out[200*8*8*bW:201*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[208*5*5:209*5*5-1]), .o_out_fmap(xor_out[208*8*8*bW:209*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[216*5*5:217*5*5-1]), .o_out_fmap(xor_out[216*8*8*bW:217*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[224*5*5:225*5*5-1]), .o_out_fmap(xor_out[224*8*8*bW:225*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[232*5*5:233*5*5-1]), .o_out_fmap(xor_out[232*8*8*bW:233*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[240*5*5:241*5*5-1]), .o_out_fmap(xor_out[240*8*8*bW:241*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[248*5*5:249*5*5-1]), .o_out_fmap(xor_out[248*8*8*bW:249*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[256*5*5:257*5*5-1]), .o_out_fmap(xor_out[256*8*8*bW:257*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[264*5*5:265*5*5-1]), .o_out_fmap(xor_out[264*8*8*bW:265*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[272*5*5:273*5*5-1]), .o_out_fmap(xor_out[272*8*8*bW:273*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[280*5*5:281*5*5-1]), .o_out_fmap(xor_out[280*8*8*bW:281*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[288*5*5:289*5*5-1]), .o_out_fmap(xor_out[288*8*8*bW:289*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[296*5*5:297*5*5-1]), .o_out_fmap(xor_out[296*8*8*bW:297*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[304*5*5:305*5*5-1]), .o_out_fmap(xor_out[304*8*8*bW:305*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[312*5*5:313*5*5-1]), .o_out_fmap(xor_out[312*8*8*bW:313*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[320*5*5:321*5*5-1]), .o_out_fmap(xor_out[320*8*8*bW:321*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[328*5*5:329*5*5-1]), .o_out_fmap(xor_out[328*8*8*bW:329*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[336*5*5:337*5*5-1]), .o_out_fmap(xor_out[336*8*8*bW:337*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[344*5*5:345*5*5-1]), .o_out_fmap(xor_out[344*8*8*bW:345*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[352*5*5:353*5*5-1]), .o_out_fmap(xor_out[352*8*8*bW:353*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[360*5*5:361*5*5-1]), .o_out_fmap(xor_out[360*8*8*bW:361*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[368*5*5:369*5*5-1]), .o_out_fmap(xor_out[368*8*8*bW:369*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[376*5*5:377*5*5-1]), .o_out_fmap(xor_out[376*8*8*bW:377*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[384*5*5:385*5*5-1]), .o_out_fmap(xor_out[384*8*8*bW:385*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[392*5*5:393*5*5-1]), .o_out_fmap(xor_out[392*8*8*bW:393*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[400*5*5:401*5*5-1]), .o_out_fmap(xor_out[400*8*8*bW:401*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[408*5*5:409*5*5-1]), .o_out_fmap(xor_out[408*8*8*bW:409*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[416*5*5:417*5*5-1]), .o_out_fmap(xor_out[416*8*8*bW:417*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[424*5*5:425*5*5-1]), .o_out_fmap(xor_out[424*8*8*bW:425*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[432*5*5:433*5*5-1]), .o_out_fmap(xor_out[432*8*8*bW:433*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[440*5*5:441*5*5-1]), .o_out_fmap(xor_out[440*8*8*bW:441*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[448*5*5:449*5*5-1]), .o_out_fmap(xor_out[448*8*8*bW:449*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[456*5*5:457*5*5-1]), .o_out_fmap(xor_out[456*8*8*bW:457*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[464*5*5:465*5*5-1]), .o_out_fmap(xor_out[464*8*8*bW:465*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[472*5*5:473*5*5-1]), .o_out_fmap(xor_out[472*8*8*bW:473*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[9*5*5:10*5*5-1]), .o_out_fmap(xor_out[9*8*8*bW:10*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[18*5*5:19*5*5-1]), .o_out_fmap(xor_out[18*8*8*bW:19*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[27*5*5:28*5*5-1]), .o_out_fmap(xor_out[27*8*8*bW:28*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[36*5*5:37*5*5-1]), .o_out_fmap(xor_out[36*8*8*bW:37*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[45*5*5:46*5*5-1]), .o_out_fmap(xor_out[45*8*8*bW:46*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[54*5*5:55*5*5-1]), .o_out_fmap(xor_out[54*8*8*bW:55*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[63*5*5:64*5*5-1]), .o_out_fmap(xor_out[63*8*8*bW:64*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[72*5*5:73*5*5-1]), .o_out_fmap(xor_out[72*8*8*bW:73*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[81*5*5:82*5*5-1]), .o_out_fmap(xor_out[81*8*8*bW:82*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[90*5*5:91*5*5-1]), .o_out_fmap(xor_out[90*8*8*bW:91*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[99*5*5:100*5*5-1]), .o_out_fmap(xor_out[99*8*8*bW:100*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[108*5*5:109*5*5-1]), .o_out_fmap(xor_out[108*8*8*bW:109*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[117*5*5:118*5*5-1]), .o_out_fmap(xor_out[117*8*8*bW:118*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[126*5*5:127*5*5-1]), .o_out_fmap(xor_out[126*8*8*bW:127*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[135*5*5:136*5*5-1]), .o_out_fmap(xor_out[135*8*8*bW:136*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[144*5*5:145*5*5-1]), .o_out_fmap(xor_out[144*8*8*bW:145*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[153*5*5:154*5*5-1]), .o_out_fmap(xor_out[153*8*8*bW:154*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[162*5*5:163*5*5-1]), .o_out_fmap(xor_out[162*8*8*bW:163*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[171*5*5:172*5*5-1]), .o_out_fmap(xor_out[171*8*8*bW:172*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[180*5*5:181*5*5-1]), .o_out_fmap(xor_out[180*8*8*bW:181*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[189*5*5:190*5*5-1]), .o_out_fmap(xor_out[189*8*8*bW:190*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[198*5*5:199*5*5-1]), .o_out_fmap(xor_out[198*8*8*bW:199*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[207*5*5:208*5*5-1]), .o_out_fmap(xor_out[207*8*8*bW:208*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[216*5*5:217*5*5-1]), .o_out_fmap(xor_out[216*8*8*bW:217*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[225*5*5:226*5*5-1]), .o_out_fmap(xor_out[225*8*8*bW:226*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[234*5*5:235*5*5-1]), .o_out_fmap(xor_out[234*8*8*bW:235*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[243*5*5:244*5*5-1]), .o_out_fmap(xor_out[243*8*8*bW:244*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[252*5*5:253*5*5-1]), .o_out_fmap(xor_out[252*8*8*bW:253*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[261*5*5:262*5*5-1]), .o_out_fmap(xor_out[261*8*8*bW:262*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[270*5*5:271*5*5-1]), .o_out_fmap(xor_out[270*8*8*bW:271*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[279*5*5:280*5*5-1]), .o_out_fmap(xor_out[279*8*8*bW:280*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[288*5*5:289*5*5-1]), .o_out_fmap(xor_out[288*8*8*bW:289*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[297*5*5:298*5*5-1]), .o_out_fmap(xor_out[297*8*8*bW:298*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[306*5*5:307*5*5-1]), .o_out_fmap(xor_out[306*8*8*bW:307*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[315*5*5:316*5*5-1]), .o_out_fmap(xor_out[315*8*8*bW:316*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[324*5*5:325*5*5-1]), .o_out_fmap(xor_out[324*8*8*bW:325*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[333*5*5:334*5*5-1]), .o_out_fmap(xor_out[333*8*8*bW:334*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[342*5*5:343*5*5-1]), .o_out_fmap(xor_out[342*8*8*bW:343*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[351*5*5:352*5*5-1]), .o_out_fmap(xor_out[351*8*8*bW:352*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[360*5*5:361*5*5-1]), .o_out_fmap(xor_out[360*8*8*bW:361*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[369*5*5:370*5*5-1]), .o_out_fmap(xor_out[369*8*8*bW:370*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[378*5*5:379*5*5-1]), .o_out_fmap(xor_out[378*8*8*bW:379*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[387*5*5:388*5*5-1]), .o_out_fmap(xor_out[387*8*8*bW:388*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[396*5*5:397*5*5-1]), .o_out_fmap(xor_out[396*8*8*bW:397*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[405*5*5:406*5*5-1]), .o_out_fmap(xor_out[405*8*8*bW:406*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[414*5*5:415*5*5-1]), .o_out_fmap(xor_out[414*8*8*bW:415*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[423*5*5:424*5*5-1]), .o_out_fmap(xor_out[423*8*8*bW:424*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[432*5*5:433*5*5-1]), .o_out_fmap(xor_out[432*8*8*bW:433*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[441*5*5:442*5*5-1]), .o_out_fmap(xor_out[441*8*8*bW:442*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[450*5*5:451*5*5-1]), .o_out_fmap(xor_out[450*8*8*bW:451*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[459*5*5:460*5*5-1]), .o_out_fmap(xor_out[459*8*8*bW:460*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[468*5*5:469*5*5-1]), .o_out_fmap(xor_out[468*8*8*bW:469*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[477*5*5:478*5*5-1]), .o_out_fmap(xor_out[477*8*8*bW:478*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[486*5*5:487*5*5-1]), .o_out_fmap(xor_out[486*8*8*bW:487*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[495*5*5:496*5*5-1]), .o_out_fmap(xor_out[495*8*8*bW:496*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[504*5*5:505*5*5-1]), .o_out_fmap(xor_out[504*8*8*bW:505*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[513*5*5:514*5*5-1]), .o_out_fmap(xor_out[513*8*8*bW:514*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[522*5*5:523*5*5-1]), .o_out_fmap(xor_out[522*8*8*bW:523*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[531*5*5:532*5*5-1]), .o_out_fmap(xor_out[531*8*8*bW:532*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[10*5*5:11*5*5-1]), .o_out_fmap(xor_out[10*8*8*bW:11*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[20*5*5:21*5*5-1]), .o_out_fmap(xor_out[20*8*8*bW:21*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[30*5*5:31*5*5-1]), .o_out_fmap(xor_out[30*8*8*bW:31*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[40*5*5:41*5*5-1]), .o_out_fmap(xor_out[40*8*8*bW:41*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[50*5*5:51*5*5-1]), .o_out_fmap(xor_out[50*8*8*bW:51*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[60*5*5:61*5*5-1]), .o_out_fmap(xor_out[60*8*8*bW:61*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[70*5*5:71*5*5-1]), .o_out_fmap(xor_out[70*8*8*bW:71*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[80*5*5:81*5*5-1]), .o_out_fmap(xor_out[80*8*8*bW:81*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[90*5*5:91*5*5-1]), .o_out_fmap(xor_out[90*8*8*bW:91*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[100*5*5:101*5*5-1]), .o_out_fmap(xor_out[100*8*8*bW:101*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[110*5*5:111*5*5-1]), .o_out_fmap(xor_out[110*8*8*bW:111*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[120*5*5:121*5*5-1]), .o_out_fmap(xor_out[120*8*8*bW:121*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[130*5*5:131*5*5-1]), .o_out_fmap(xor_out[130*8*8*bW:131*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[140*5*5:141*5*5-1]), .o_out_fmap(xor_out[140*8*8*bW:141*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[150*5*5:151*5*5-1]), .o_out_fmap(xor_out[150*8*8*bW:151*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[160*5*5:161*5*5-1]), .o_out_fmap(xor_out[160*8*8*bW:161*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[170*5*5:171*5*5-1]), .o_out_fmap(xor_out[170*8*8*bW:171*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[180*5*5:181*5*5-1]), .o_out_fmap(xor_out[180*8*8*bW:181*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[190*5*5:191*5*5-1]), .o_out_fmap(xor_out[190*8*8*bW:191*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[200*5*5:201*5*5-1]), .o_out_fmap(xor_out[200*8*8*bW:201*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[210*5*5:211*5*5-1]), .o_out_fmap(xor_out[210*8*8*bW:211*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[220*5*5:221*5*5-1]), .o_out_fmap(xor_out[220*8*8*bW:221*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[230*5*5:231*5*5-1]), .o_out_fmap(xor_out[230*8*8*bW:231*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[240*5*5:241*5*5-1]), .o_out_fmap(xor_out[240*8*8*bW:241*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[250*5*5:251*5*5-1]), .o_out_fmap(xor_out[250*8*8*bW:251*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[260*5*5:261*5*5-1]), .o_out_fmap(xor_out[260*8*8*bW:261*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[270*5*5:271*5*5-1]), .o_out_fmap(xor_out[270*8*8*bW:271*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[280*5*5:281*5*5-1]), .o_out_fmap(xor_out[280*8*8*bW:281*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[290*5*5:291*5*5-1]), .o_out_fmap(xor_out[290*8*8*bW:291*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[300*5*5:301*5*5-1]), .o_out_fmap(xor_out[300*8*8*bW:301*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[310*5*5:311*5*5-1]), .o_out_fmap(xor_out[310*8*8*bW:311*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[320*5*5:321*5*5-1]), .o_out_fmap(xor_out[320*8*8*bW:321*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[330*5*5:331*5*5-1]), .o_out_fmap(xor_out[330*8*8*bW:331*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[340*5*5:341*5*5-1]), .o_out_fmap(xor_out[340*8*8*bW:341*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[350*5*5:351*5*5-1]), .o_out_fmap(xor_out[350*8*8*bW:351*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[360*5*5:361*5*5-1]), .o_out_fmap(xor_out[360*8*8*bW:361*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[370*5*5:371*5*5-1]), .o_out_fmap(xor_out[370*8*8*bW:371*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[380*5*5:381*5*5-1]), .o_out_fmap(xor_out[380*8*8*bW:381*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[390*5*5:391*5*5-1]), .o_out_fmap(xor_out[390*8*8*bW:391*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[400*5*5:401*5*5-1]), .o_out_fmap(xor_out[400*8*8*bW:401*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[410*5*5:411*5*5-1]), .o_out_fmap(xor_out[410*8*8*bW:411*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[420*5*5:421*5*5-1]), .o_out_fmap(xor_out[420*8*8*bW:421*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[430*5*5:431*5*5-1]), .o_out_fmap(xor_out[430*8*8*bW:431*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[440*5*5:441*5*5-1]), .o_out_fmap(xor_out[440*8*8*bW:441*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[450*5*5:451*5*5-1]), .o_out_fmap(xor_out[450*8*8*bW:451*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[460*5*5:461*5*5-1]), .o_out_fmap(xor_out[460*8*8*bW:461*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[470*5*5:471*5*5-1]), .o_out_fmap(xor_out[470*8*8*bW:471*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[480*5*5:481*5*5-1]), .o_out_fmap(xor_out[480*8*8*bW:481*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[490*5*5:491*5*5-1]), .o_out_fmap(xor_out[490*8*8*bW:491*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[500*5*5:501*5*5-1]), .o_out_fmap(xor_out[500*8*8*bW:501*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[510*5*5:511*5*5-1]), .o_out_fmap(xor_out[510*8*8*bW:511*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[520*5*5:521*5*5-1]), .o_out_fmap(xor_out[520*8*8*bW:521*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[530*5*5:531*5*5-1]), .o_out_fmap(xor_out[530*8*8*bW:531*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[540*5*5:541*5*5-1]), .o_out_fmap(xor_out[540*8*8*bW:541*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[550*5*5:551*5*5-1]), .o_out_fmap(xor_out[550*8*8*bW:551*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[560*5*5:561*5*5-1]), .o_out_fmap(xor_out[560*8*8*bW:561*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[570*5*5:571*5*5-1]), .o_out_fmap(xor_out[570*8*8*bW:571*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[580*5*5:581*5*5-1]), .o_out_fmap(xor_out[580*8*8*bW:581*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[590*5*5:591*5*5-1]), .o_out_fmap(xor_out[590*8*8*bW:591*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[11*5*5:12*5*5-1]), .o_out_fmap(xor_out[11*8*8*bW:12*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[22*5*5:23*5*5-1]), .o_out_fmap(xor_out[22*8*8*bW:23*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[33*5*5:34*5*5-1]), .o_out_fmap(xor_out[33*8*8*bW:34*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[44*5*5:45*5*5-1]), .o_out_fmap(xor_out[44*8*8*bW:45*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[55*5*5:56*5*5-1]), .o_out_fmap(xor_out[55*8*8*bW:56*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[66*5*5:67*5*5-1]), .o_out_fmap(xor_out[66*8*8*bW:67*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[77*5*5:78*5*5-1]), .o_out_fmap(xor_out[77*8*8*bW:78*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[88*5*5:89*5*5-1]), .o_out_fmap(xor_out[88*8*8*bW:89*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[99*5*5:100*5*5-1]), .o_out_fmap(xor_out[99*8*8*bW:100*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[110*5*5:111*5*5-1]), .o_out_fmap(xor_out[110*8*8*bW:111*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[121*5*5:122*5*5-1]), .o_out_fmap(xor_out[121*8*8*bW:122*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[132*5*5:133*5*5-1]), .o_out_fmap(xor_out[132*8*8*bW:133*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[143*5*5:144*5*5-1]), .o_out_fmap(xor_out[143*8*8*bW:144*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[154*5*5:155*5*5-1]), .o_out_fmap(xor_out[154*8*8*bW:155*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[165*5*5:166*5*5-1]), .o_out_fmap(xor_out[165*8*8*bW:166*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[176*5*5:177*5*5-1]), .o_out_fmap(xor_out[176*8*8*bW:177*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[187*5*5:188*5*5-1]), .o_out_fmap(xor_out[187*8*8*bW:188*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[198*5*5:199*5*5-1]), .o_out_fmap(xor_out[198*8*8*bW:199*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[209*5*5:210*5*5-1]), .o_out_fmap(xor_out[209*8*8*bW:210*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[220*5*5:221*5*5-1]), .o_out_fmap(xor_out[220*8*8*bW:221*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[231*5*5:232*5*5-1]), .o_out_fmap(xor_out[231*8*8*bW:232*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[242*5*5:243*5*5-1]), .o_out_fmap(xor_out[242*8*8*bW:243*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[253*5*5:254*5*5-1]), .o_out_fmap(xor_out[253*8*8*bW:254*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[264*5*5:265*5*5-1]), .o_out_fmap(xor_out[264*8*8*bW:265*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[275*5*5:276*5*5-1]), .o_out_fmap(xor_out[275*8*8*bW:276*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[286*5*5:287*5*5-1]), .o_out_fmap(xor_out[286*8*8*bW:287*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[297*5*5:298*5*5-1]), .o_out_fmap(xor_out[297*8*8*bW:298*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[308*5*5:309*5*5-1]), .o_out_fmap(xor_out[308*8*8*bW:309*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[319*5*5:320*5*5-1]), .o_out_fmap(xor_out[319*8*8*bW:320*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[330*5*5:331*5*5-1]), .o_out_fmap(xor_out[330*8*8*bW:331*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[341*5*5:342*5*5-1]), .o_out_fmap(xor_out[341*8*8*bW:342*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[352*5*5:353*5*5-1]), .o_out_fmap(xor_out[352*8*8*bW:353*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[363*5*5:364*5*5-1]), .o_out_fmap(xor_out[363*8*8*bW:364*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[374*5*5:375*5*5-1]), .o_out_fmap(xor_out[374*8*8*bW:375*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[385*5*5:386*5*5-1]), .o_out_fmap(xor_out[385*8*8*bW:386*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[396*5*5:397*5*5-1]), .o_out_fmap(xor_out[396*8*8*bW:397*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[407*5*5:408*5*5-1]), .o_out_fmap(xor_out[407*8*8*bW:408*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[418*5*5:419*5*5-1]), .o_out_fmap(xor_out[418*8*8*bW:419*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[429*5*5:430*5*5-1]), .o_out_fmap(xor_out[429*8*8*bW:430*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[440*5*5:441*5*5-1]), .o_out_fmap(xor_out[440*8*8*bW:441*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[451*5*5:452*5*5-1]), .o_out_fmap(xor_out[451*8*8*bW:452*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[462*5*5:463*5*5-1]), .o_out_fmap(xor_out[462*8*8*bW:463*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[473*5*5:474*5*5-1]), .o_out_fmap(xor_out[473*8*8*bW:474*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[484*5*5:485*5*5-1]), .o_out_fmap(xor_out[484*8*8*bW:485*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[495*5*5:496*5*5-1]), .o_out_fmap(xor_out[495*8*8*bW:496*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[506*5*5:507*5*5-1]), .o_out_fmap(xor_out[506*8*8*bW:507*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[517*5*5:518*5*5-1]), .o_out_fmap(xor_out[517*8*8*bW:518*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[528*5*5:529*5*5-1]), .o_out_fmap(xor_out[528*8*8*bW:529*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[539*5*5:540*5*5-1]), .o_out_fmap(xor_out[539*8*8*bW:540*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[550*5*5:551*5*5-1]), .o_out_fmap(xor_out[550*8*8*bW:551*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[561*5*5:562*5*5-1]), .o_out_fmap(xor_out[561*8*8*bW:562*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[572*5*5:573*5*5-1]), .o_out_fmap(xor_out[572*8*8*bW:573*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[583*5*5:584*5*5-1]), .o_out_fmap(xor_out[583*8*8*bW:584*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[594*5*5:595*5*5-1]), .o_out_fmap(xor_out[594*8*8*bW:595*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[605*5*5:606*5*5-1]), .o_out_fmap(xor_out[605*8*8*bW:606*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[616*5*5:617*5*5-1]), .o_out_fmap(xor_out[616*8*8*bW:617*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[627*5*5:628*5*5-1]), .o_out_fmap(xor_out[627*8*8*bW:628*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[638*5*5:639*5*5-1]), .o_out_fmap(xor_out[638*8*8*bW:639*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[649*5*5:650*5*5-1]), .o_out_fmap(xor_out[649*8*8*bW:650*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[12*5*5:13*5*5-1]), .o_out_fmap(xor_out[12*8*8*bW:13*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[24*5*5:25*5*5-1]), .o_out_fmap(xor_out[24*8*8*bW:25*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[36*5*5:37*5*5-1]), .o_out_fmap(xor_out[36*8*8*bW:37*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[48*5*5:49*5*5-1]), .o_out_fmap(xor_out[48*8*8*bW:49*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[60*5*5:61*5*5-1]), .o_out_fmap(xor_out[60*8*8*bW:61*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[72*5*5:73*5*5-1]), .o_out_fmap(xor_out[72*8*8*bW:73*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[84*5*5:85*5*5-1]), .o_out_fmap(xor_out[84*8*8*bW:85*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[96*5*5:97*5*5-1]), .o_out_fmap(xor_out[96*8*8*bW:97*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[108*5*5:109*5*5-1]), .o_out_fmap(xor_out[108*8*8*bW:109*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[120*5*5:121*5*5-1]), .o_out_fmap(xor_out[120*8*8*bW:121*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[132*5*5:133*5*5-1]), .o_out_fmap(xor_out[132*8*8*bW:133*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[144*5*5:145*5*5-1]), .o_out_fmap(xor_out[144*8*8*bW:145*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[156*5*5:157*5*5-1]), .o_out_fmap(xor_out[156*8*8*bW:157*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[168*5*5:169*5*5-1]), .o_out_fmap(xor_out[168*8*8*bW:169*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[180*5*5:181*5*5-1]), .o_out_fmap(xor_out[180*8*8*bW:181*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[192*5*5:193*5*5-1]), .o_out_fmap(xor_out[192*8*8*bW:193*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[204*5*5:205*5*5-1]), .o_out_fmap(xor_out[204*8*8*bW:205*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[216*5*5:217*5*5-1]), .o_out_fmap(xor_out[216*8*8*bW:217*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[228*5*5:229*5*5-1]), .o_out_fmap(xor_out[228*8*8*bW:229*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[240*5*5:241*5*5-1]), .o_out_fmap(xor_out[240*8*8*bW:241*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[252*5*5:253*5*5-1]), .o_out_fmap(xor_out[252*8*8*bW:253*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[264*5*5:265*5*5-1]), .o_out_fmap(xor_out[264*8*8*bW:265*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[276*5*5:277*5*5-1]), .o_out_fmap(xor_out[276*8*8*bW:277*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[288*5*5:289*5*5-1]), .o_out_fmap(xor_out[288*8*8*bW:289*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[300*5*5:301*5*5-1]), .o_out_fmap(xor_out[300*8*8*bW:301*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[312*5*5:313*5*5-1]), .o_out_fmap(xor_out[312*8*8*bW:313*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[324*5*5:325*5*5-1]), .o_out_fmap(xor_out[324*8*8*bW:325*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[336*5*5:337*5*5-1]), .o_out_fmap(xor_out[336*8*8*bW:337*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[348*5*5:349*5*5-1]), .o_out_fmap(xor_out[348*8*8*bW:349*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[360*5*5:361*5*5-1]), .o_out_fmap(xor_out[360*8*8*bW:361*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[372*5*5:373*5*5-1]), .o_out_fmap(xor_out[372*8*8*bW:373*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[384*5*5:385*5*5-1]), .o_out_fmap(xor_out[384*8*8*bW:385*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[396*5*5:397*5*5-1]), .o_out_fmap(xor_out[396*8*8*bW:397*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[408*5*5:409*5*5-1]), .o_out_fmap(xor_out[408*8*8*bW:409*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[420*5*5:421*5*5-1]), .o_out_fmap(xor_out[420*8*8*bW:421*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[432*5*5:433*5*5-1]), .o_out_fmap(xor_out[432*8*8*bW:433*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[444*5*5:445*5*5-1]), .o_out_fmap(xor_out[444*8*8*bW:445*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[456*5*5:457*5*5-1]), .o_out_fmap(xor_out[456*8*8*bW:457*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[468*5*5:469*5*5-1]), .o_out_fmap(xor_out[468*8*8*bW:469*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[480*5*5:481*5*5-1]), .o_out_fmap(xor_out[480*8*8*bW:481*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[492*5*5:493*5*5-1]), .o_out_fmap(xor_out[492*8*8*bW:493*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[504*5*5:505*5*5-1]), .o_out_fmap(xor_out[504*8*8*bW:505*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[516*5*5:517*5*5-1]), .o_out_fmap(xor_out[516*8*8*bW:517*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[528*5*5:529*5*5-1]), .o_out_fmap(xor_out[528*8*8*bW:529*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[540*5*5:541*5*5-1]), .o_out_fmap(xor_out[540*8*8*bW:541*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[552*5*5:553*5*5-1]), .o_out_fmap(xor_out[552*8*8*bW:553*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[564*5*5:565*5*5-1]), .o_out_fmap(xor_out[564*8*8*bW:565*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[576*5*5:577*5*5-1]), .o_out_fmap(xor_out[576*8*8*bW:577*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[588*5*5:589*5*5-1]), .o_out_fmap(xor_out[588*8*8*bW:589*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[600*5*5:601*5*5-1]), .o_out_fmap(xor_out[600*8*8*bW:601*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[612*5*5:613*5*5-1]), .o_out_fmap(xor_out[612*8*8*bW:613*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[624*5*5:625*5*5-1]), .o_out_fmap(xor_out[624*8*8*bW:625*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[636*5*5:637*5*5-1]), .o_out_fmap(xor_out[636*8*8*bW:637*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[648*5*5:649*5*5-1]), .o_out_fmap(xor_out[648*8*8*bW:649*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[660*5*5:661*5*5-1]), .o_out_fmap(xor_out[660*8*8*bW:661*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[672*5*5:673*5*5-1]), .o_out_fmap(xor_out[672*8*8*bW:673*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[684*5*5:685*5*5-1]), .o_out_fmap(xor_out[684*8*8*bW:685*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[696*5*5:697*5*5-1]), .o_out_fmap(xor_out[696*8*8*bW:697*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[708*5*5:709*5*5-1]), .o_out_fmap(xor_out[708*8*8*bW:709*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[13*5*5:14*5*5-1]), .o_out_fmap(xor_out[13*8*8*bW:14*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[26*5*5:27*5*5-1]), .o_out_fmap(xor_out[26*8*8*bW:27*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[39*5*5:40*5*5-1]), .o_out_fmap(xor_out[39*8*8*bW:40*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[52*5*5:53*5*5-1]), .o_out_fmap(xor_out[52*8*8*bW:53*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[65*5*5:66*5*5-1]), .o_out_fmap(xor_out[65*8*8*bW:66*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[78*5*5:79*5*5-1]), .o_out_fmap(xor_out[78*8*8*bW:79*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[91*5*5:92*5*5-1]), .o_out_fmap(xor_out[91*8*8*bW:92*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[104*5*5:105*5*5-1]), .o_out_fmap(xor_out[104*8*8*bW:105*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[117*5*5:118*5*5-1]), .o_out_fmap(xor_out[117*8*8*bW:118*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[130*5*5:131*5*5-1]), .o_out_fmap(xor_out[130*8*8*bW:131*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[143*5*5:144*5*5-1]), .o_out_fmap(xor_out[143*8*8*bW:144*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[156*5*5:157*5*5-1]), .o_out_fmap(xor_out[156*8*8*bW:157*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[169*5*5:170*5*5-1]), .o_out_fmap(xor_out[169*8*8*bW:170*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[182*5*5:183*5*5-1]), .o_out_fmap(xor_out[182*8*8*bW:183*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[195*5*5:196*5*5-1]), .o_out_fmap(xor_out[195*8*8*bW:196*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[208*5*5:209*5*5-1]), .o_out_fmap(xor_out[208*8*8*bW:209*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[221*5*5:222*5*5-1]), .o_out_fmap(xor_out[221*8*8*bW:222*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[234*5*5:235*5*5-1]), .o_out_fmap(xor_out[234*8*8*bW:235*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[247*5*5:248*5*5-1]), .o_out_fmap(xor_out[247*8*8*bW:248*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[260*5*5:261*5*5-1]), .o_out_fmap(xor_out[260*8*8*bW:261*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[273*5*5:274*5*5-1]), .o_out_fmap(xor_out[273*8*8*bW:274*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[286*5*5:287*5*5-1]), .o_out_fmap(xor_out[286*8*8*bW:287*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[299*5*5:300*5*5-1]), .o_out_fmap(xor_out[299*8*8*bW:300*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[312*5*5:313*5*5-1]), .o_out_fmap(xor_out[312*8*8*bW:313*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[325*5*5:326*5*5-1]), .o_out_fmap(xor_out[325*8*8*bW:326*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[338*5*5:339*5*5-1]), .o_out_fmap(xor_out[338*8*8*bW:339*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[351*5*5:352*5*5-1]), .o_out_fmap(xor_out[351*8*8*bW:352*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[364*5*5:365*5*5-1]), .o_out_fmap(xor_out[364*8*8*bW:365*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[377*5*5:378*5*5-1]), .o_out_fmap(xor_out[377*8*8*bW:378*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[390*5*5:391*5*5-1]), .o_out_fmap(xor_out[390*8*8*bW:391*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[403*5*5:404*5*5-1]), .o_out_fmap(xor_out[403*8*8*bW:404*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[416*5*5:417*5*5-1]), .o_out_fmap(xor_out[416*8*8*bW:417*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[429*5*5:430*5*5-1]), .o_out_fmap(xor_out[429*8*8*bW:430*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[442*5*5:443*5*5-1]), .o_out_fmap(xor_out[442*8*8*bW:443*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[455*5*5:456*5*5-1]), .o_out_fmap(xor_out[455*8*8*bW:456*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[468*5*5:469*5*5-1]), .o_out_fmap(xor_out[468*8*8*bW:469*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[481*5*5:482*5*5-1]), .o_out_fmap(xor_out[481*8*8*bW:482*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[494*5*5:495*5*5-1]), .o_out_fmap(xor_out[494*8*8*bW:495*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[507*5*5:508*5*5-1]), .o_out_fmap(xor_out[507*8*8*bW:508*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[520*5*5:521*5*5-1]), .o_out_fmap(xor_out[520*8*8*bW:521*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[533*5*5:534*5*5-1]), .o_out_fmap(xor_out[533*8*8*bW:534*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[546*5*5:547*5*5-1]), .o_out_fmap(xor_out[546*8*8*bW:547*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[559*5*5:560*5*5-1]), .o_out_fmap(xor_out[559*8*8*bW:560*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[572*5*5:573*5*5-1]), .o_out_fmap(xor_out[572*8*8*bW:573*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[585*5*5:586*5*5-1]), .o_out_fmap(xor_out[585*8*8*bW:586*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[598*5*5:599*5*5-1]), .o_out_fmap(xor_out[598*8*8*bW:599*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[611*5*5:612*5*5-1]), .o_out_fmap(xor_out[611*8*8*bW:612*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[624*5*5:625*5*5-1]), .o_out_fmap(xor_out[624*8*8*bW:625*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[637*5*5:638*5*5-1]), .o_out_fmap(xor_out[637*8*8*bW:638*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[650*5*5:651*5*5-1]), .o_out_fmap(xor_out[650*8*8*bW:651*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[663*5*5:664*5*5-1]), .o_out_fmap(xor_out[663*8*8*bW:664*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[676*5*5:677*5*5-1]), .o_out_fmap(xor_out[676*8*8*bW:677*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[689*5*5:690*5*5-1]), .o_out_fmap(xor_out[689*8*8*bW:690*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[702*5*5:703*5*5-1]), .o_out_fmap(xor_out[702*8*8*bW:703*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[715*5*5:716*5*5-1]), .o_out_fmap(xor_out[715*8*8*bW:716*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[728*5*5:729*5*5-1]), .o_out_fmap(xor_out[728*8*8*bW:729*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[741*5*5:742*5*5-1]), .o_out_fmap(xor_out[741*8*8*bW:742*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[754*5*5:755*5*5-1]), .o_out_fmap(xor_out[754*8*8*bW:755*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[767*5*5:768*5*5-1]), .o_out_fmap(xor_out[767*8*8*bW:768*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[14*5*5:15*5*5-1]), .o_out_fmap(xor_out[14*8*8*bW:15*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[28*5*5:29*5*5-1]), .o_out_fmap(xor_out[28*8*8*bW:29*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[42*5*5:43*5*5-1]), .o_out_fmap(xor_out[42*8*8*bW:43*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[56*5*5:57*5*5-1]), .o_out_fmap(xor_out[56*8*8*bW:57*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[70*5*5:71*5*5-1]), .o_out_fmap(xor_out[70*8*8*bW:71*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[84*5*5:85*5*5-1]), .o_out_fmap(xor_out[84*8*8*bW:85*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[98*5*5:99*5*5-1]), .o_out_fmap(xor_out[98*8*8*bW:99*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[112*5*5:113*5*5-1]), .o_out_fmap(xor_out[112*8*8*bW:113*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[126*5*5:127*5*5-1]), .o_out_fmap(xor_out[126*8*8*bW:127*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[140*5*5:141*5*5-1]), .o_out_fmap(xor_out[140*8*8*bW:141*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[154*5*5:155*5*5-1]), .o_out_fmap(xor_out[154*8*8*bW:155*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[168*5*5:169*5*5-1]), .o_out_fmap(xor_out[168*8*8*bW:169*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[182*5*5:183*5*5-1]), .o_out_fmap(xor_out[182*8*8*bW:183*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[196*5*5:197*5*5-1]), .o_out_fmap(xor_out[196*8*8*bW:197*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[210*5*5:211*5*5-1]), .o_out_fmap(xor_out[210*8*8*bW:211*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[224*5*5:225*5*5-1]), .o_out_fmap(xor_out[224*8*8*bW:225*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[238*5*5:239*5*5-1]), .o_out_fmap(xor_out[238*8*8*bW:239*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[252*5*5:253*5*5-1]), .o_out_fmap(xor_out[252*8*8*bW:253*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[266*5*5:267*5*5-1]), .o_out_fmap(xor_out[266*8*8*bW:267*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[280*5*5:281*5*5-1]), .o_out_fmap(xor_out[280*8*8*bW:281*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[294*5*5:295*5*5-1]), .o_out_fmap(xor_out[294*8*8*bW:295*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[308*5*5:309*5*5-1]), .o_out_fmap(xor_out[308*8*8*bW:309*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[322*5*5:323*5*5-1]), .o_out_fmap(xor_out[322*8*8*bW:323*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[336*5*5:337*5*5-1]), .o_out_fmap(xor_out[336*8*8*bW:337*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[350*5*5:351*5*5-1]), .o_out_fmap(xor_out[350*8*8*bW:351*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[364*5*5:365*5*5-1]), .o_out_fmap(xor_out[364*8*8*bW:365*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[378*5*5:379*5*5-1]), .o_out_fmap(xor_out[378*8*8*bW:379*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[392*5*5:393*5*5-1]), .o_out_fmap(xor_out[392*8*8*bW:393*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[406*5*5:407*5*5-1]), .o_out_fmap(xor_out[406*8*8*bW:407*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[420*5*5:421*5*5-1]), .o_out_fmap(xor_out[420*8*8*bW:421*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[434*5*5:435*5*5-1]), .o_out_fmap(xor_out[434*8*8*bW:435*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[448*5*5:449*5*5-1]), .o_out_fmap(xor_out[448*8*8*bW:449*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[462*5*5:463*5*5-1]), .o_out_fmap(xor_out[462*8*8*bW:463*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[476*5*5:477*5*5-1]), .o_out_fmap(xor_out[476*8*8*bW:477*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[490*5*5:491*5*5-1]), .o_out_fmap(xor_out[490*8*8*bW:491*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[504*5*5:505*5*5-1]), .o_out_fmap(xor_out[504*8*8*bW:505*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[518*5*5:519*5*5-1]), .o_out_fmap(xor_out[518*8*8*bW:519*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[532*5*5:533*5*5-1]), .o_out_fmap(xor_out[532*8*8*bW:533*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[546*5*5:547*5*5-1]), .o_out_fmap(xor_out[546*8*8*bW:547*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[560*5*5:561*5*5-1]), .o_out_fmap(xor_out[560*8*8*bW:561*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[574*5*5:575*5*5-1]), .o_out_fmap(xor_out[574*8*8*bW:575*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[588*5*5:589*5*5-1]), .o_out_fmap(xor_out[588*8*8*bW:589*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[602*5*5:603*5*5-1]), .o_out_fmap(xor_out[602*8*8*bW:603*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[616*5*5:617*5*5-1]), .o_out_fmap(xor_out[616*8*8*bW:617*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[630*5*5:631*5*5-1]), .o_out_fmap(xor_out[630*8*8*bW:631*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[644*5*5:645*5*5-1]), .o_out_fmap(xor_out[644*8*8*bW:645*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[658*5*5:659*5*5-1]), .o_out_fmap(xor_out[658*8*8*bW:659*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[672*5*5:673*5*5-1]), .o_out_fmap(xor_out[672*8*8*bW:673*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[686*5*5:687*5*5-1]), .o_out_fmap(xor_out[686*8*8*bW:687*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[700*5*5:701*5*5-1]), .o_out_fmap(xor_out[700*8*8*bW:701*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[714*5*5:715*5*5-1]), .o_out_fmap(xor_out[714*8*8*bW:715*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[728*5*5:729*5*5-1]), .o_out_fmap(xor_out[728*8*8*bW:729*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[742*5*5:743*5*5-1]), .o_out_fmap(xor_out[742*8*8*bW:743*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[756*5*5:757*5*5-1]), .o_out_fmap(xor_out[756*8*8*bW:757*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[770*5*5:771*5*5-1]), .o_out_fmap(xor_out[770*8*8*bW:771*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[784*5*5:785*5*5-1]), .o_out_fmap(xor_out[784*8*8*bW:785*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[798*5*5:799*5*5-1]), .o_out_fmap(xor_out[798*8*8*bW:799*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[812*5*5:813*5*5-1]), .o_out_fmap(xor_out[812*8*8*bW:813*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[826*5*5:827*5*5-1]), .o_out_fmap(xor_out[826*8*8*bW:827*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[15*5*5:16*5*5-1]), .o_out_fmap(xor_out[15*8*8*bW:16*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[30*5*5:31*5*5-1]), .o_out_fmap(xor_out[30*8*8*bW:31*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[45*5*5:46*5*5-1]), .o_out_fmap(xor_out[45*8*8*bW:46*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[60*5*5:61*5*5-1]), .o_out_fmap(xor_out[60*8*8*bW:61*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[75*5*5:76*5*5-1]), .o_out_fmap(xor_out[75*8*8*bW:76*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[90*5*5:91*5*5-1]), .o_out_fmap(xor_out[90*8*8*bW:91*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[105*5*5:106*5*5-1]), .o_out_fmap(xor_out[105*8*8*bW:106*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[120*5*5:121*5*5-1]), .o_out_fmap(xor_out[120*8*8*bW:121*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[135*5*5:136*5*5-1]), .o_out_fmap(xor_out[135*8*8*bW:136*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[150*5*5:151*5*5-1]), .o_out_fmap(xor_out[150*8*8*bW:151*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[165*5*5:166*5*5-1]), .o_out_fmap(xor_out[165*8*8*bW:166*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[180*5*5:181*5*5-1]), .o_out_fmap(xor_out[180*8*8*bW:181*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[195*5*5:196*5*5-1]), .o_out_fmap(xor_out[195*8*8*bW:196*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[210*5*5:211*5*5-1]), .o_out_fmap(xor_out[210*8*8*bW:211*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[225*5*5:226*5*5-1]), .o_out_fmap(xor_out[225*8*8*bW:226*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[240*5*5:241*5*5-1]), .o_out_fmap(xor_out[240*8*8*bW:241*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[255*5*5:256*5*5-1]), .o_out_fmap(xor_out[255*8*8*bW:256*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[270*5*5:271*5*5-1]), .o_out_fmap(xor_out[270*8*8*bW:271*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[285*5*5:286*5*5-1]), .o_out_fmap(xor_out[285*8*8*bW:286*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[300*5*5:301*5*5-1]), .o_out_fmap(xor_out[300*8*8*bW:301*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[315*5*5:316*5*5-1]), .o_out_fmap(xor_out[315*8*8*bW:316*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[330*5*5:331*5*5-1]), .o_out_fmap(xor_out[330*8*8*bW:331*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[345*5*5:346*5*5-1]), .o_out_fmap(xor_out[345*8*8*bW:346*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[360*5*5:361*5*5-1]), .o_out_fmap(xor_out[360*8*8*bW:361*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[375*5*5:376*5*5-1]), .o_out_fmap(xor_out[375*8*8*bW:376*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[390*5*5:391*5*5-1]), .o_out_fmap(xor_out[390*8*8*bW:391*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[405*5*5:406*5*5-1]), .o_out_fmap(xor_out[405*8*8*bW:406*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[420*5*5:421*5*5-1]), .o_out_fmap(xor_out[420*8*8*bW:421*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[435*5*5:436*5*5-1]), .o_out_fmap(xor_out[435*8*8*bW:436*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[450*5*5:451*5*5-1]), .o_out_fmap(xor_out[450*8*8*bW:451*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[465*5*5:466*5*5-1]), .o_out_fmap(xor_out[465*8*8*bW:466*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[480*5*5:481*5*5-1]), .o_out_fmap(xor_out[480*8*8*bW:481*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[495*5*5:496*5*5-1]), .o_out_fmap(xor_out[495*8*8*bW:496*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[510*5*5:511*5*5-1]), .o_out_fmap(xor_out[510*8*8*bW:511*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[525*5*5:526*5*5-1]), .o_out_fmap(xor_out[525*8*8*bW:526*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[540*5*5:541*5*5-1]), .o_out_fmap(xor_out[540*8*8*bW:541*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[555*5*5:556*5*5-1]), .o_out_fmap(xor_out[555*8*8*bW:556*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[570*5*5:571*5*5-1]), .o_out_fmap(xor_out[570*8*8*bW:571*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[585*5*5:586*5*5-1]), .o_out_fmap(xor_out[585*8*8*bW:586*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[600*5*5:601*5*5-1]), .o_out_fmap(xor_out[600*8*8*bW:601*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[615*5*5:616*5*5-1]), .o_out_fmap(xor_out[615*8*8*bW:616*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[630*5*5:631*5*5-1]), .o_out_fmap(xor_out[630*8*8*bW:631*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[645*5*5:646*5*5-1]), .o_out_fmap(xor_out[645*8*8*bW:646*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[660*5*5:661*5*5-1]), .o_out_fmap(xor_out[660*8*8*bW:661*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[675*5*5:676*5*5-1]), .o_out_fmap(xor_out[675*8*8*bW:676*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[690*5*5:691*5*5-1]), .o_out_fmap(xor_out[690*8*8*bW:691*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[705*5*5:706*5*5-1]), .o_out_fmap(xor_out[705*8*8*bW:706*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[720*5*5:721*5*5-1]), .o_out_fmap(xor_out[720*8*8*bW:721*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[735*5*5:736*5*5-1]), .o_out_fmap(xor_out[735*8*8*bW:736*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[750*5*5:751*5*5-1]), .o_out_fmap(xor_out[750*8*8*bW:751*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[765*5*5:766*5*5-1]), .o_out_fmap(xor_out[765*8*8*bW:766*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[780*5*5:781*5*5-1]), .o_out_fmap(xor_out[780*8*8*bW:781*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[795*5*5:796*5*5-1]), .o_out_fmap(xor_out[795*8*8*bW:796*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[810*5*5:811*5*5-1]), .o_out_fmap(xor_out[810*8*8*bW:811*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[825*5*5:826*5*5-1]), .o_out_fmap(xor_out[825*8*8*bW:826*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[840*5*5:841*5*5-1]), .o_out_fmap(xor_out[840*8*8*bW:841*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[855*5*5:856*5*5-1]), .o_out_fmap(xor_out[855*8*8*bW:856*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[870*5*5:871*5*5-1]), .o_out_fmap(xor_out[870*8*8*bW:871*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[885*5*5:886*5*5-1]), .o_out_fmap(xor_out[885*8*8*bW:886*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[16*5*5:17*5*5-1]), .o_out_fmap(xor_out[16*8*8*bW:17*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[32*5*5:33*5*5-1]), .o_out_fmap(xor_out[32*8*8*bW:33*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[48*5*5:49*5*5-1]), .o_out_fmap(xor_out[48*8*8*bW:49*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[64*5*5:65*5*5-1]), .o_out_fmap(xor_out[64*8*8*bW:65*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[80*5*5:81*5*5-1]), .o_out_fmap(xor_out[80*8*8*bW:81*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[96*5*5:97*5*5-1]), .o_out_fmap(xor_out[96*8*8*bW:97*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[112*5*5:113*5*5-1]), .o_out_fmap(xor_out[112*8*8*bW:113*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[128*5*5:129*5*5-1]), .o_out_fmap(xor_out[128*8*8*bW:129*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[144*5*5:145*5*5-1]), .o_out_fmap(xor_out[144*8*8*bW:145*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[160*5*5:161*5*5-1]), .o_out_fmap(xor_out[160*8*8*bW:161*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[176*5*5:177*5*5-1]), .o_out_fmap(xor_out[176*8*8*bW:177*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[192*5*5:193*5*5-1]), .o_out_fmap(xor_out[192*8*8*bW:193*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[208*5*5:209*5*5-1]), .o_out_fmap(xor_out[208*8*8*bW:209*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[224*5*5:225*5*5-1]), .o_out_fmap(xor_out[224*8*8*bW:225*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[240*5*5:241*5*5-1]), .o_out_fmap(xor_out[240*8*8*bW:241*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[256*5*5:257*5*5-1]), .o_out_fmap(xor_out[256*8*8*bW:257*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[272*5*5:273*5*5-1]), .o_out_fmap(xor_out[272*8*8*bW:273*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[288*5*5:289*5*5-1]), .o_out_fmap(xor_out[288*8*8*bW:289*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[304*5*5:305*5*5-1]), .o_out_fmap(xor_out[304*8*8*bW:305*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[320*5*5:321*5*5-1]), .o_out_fmap(xor_out[320*8*8*bW:321*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[336*5*5:337*5*5-1]), .o_out_fmap(xor_out[336*8*8*bW:337*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[352*5*5:353*5*5-1]), .o_out_fmap(xor_out[352*8*8*bW:353*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[368*5*5:369*5*5-1]), .o_out_fmap(xor_out[368*8*8*bW:369*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[384*5*5:385*5*5-1]), .o_out_fmap(xor_out[384*8*8*bW:385*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[400*5*5:401*5*5-1]), .o_out_fmap(xor_out[400*8*8*bW:401*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[416*5*5:417*5*5-1]), .o_out_fmap(xor_out[416*8*8*bW:417*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[432*5*5:433*5*5-1]), .o_out_fmap(xor_out[432*8*8*bW:433*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[448*5*5:449*5*5-1]), .o_out_fmap(xor_out[448*8*8*bW:449*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[464*5*5:465*5*5-1]), .o_out_fmap(xor_out[464*8*8*bW:465*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[480*5*5:481*5*5-1]), .o_out_fmap(xor_out[480*8*8*bW:481*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[496*5*5:497*5*5-1]), .o_out_fmap(xor_out[496*8*8*bW:497*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[512*5*5:513*5*5-1]), .o_out_fmap(xor_out[512*8*8*bW:513*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[528*5*5:529*5*5-1]), .o_out_fmap(xor_out[528*8*8*bW:529*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[544*5*5:545*5*5-1]), .o_out_fmap(xor_out[544*8*8*bW:545*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[560*5*5:561*5*5-1]), .o_out_fmap(xor_out[560*8*8*bW:561*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[576*5*5:577*5*5-1]), .o_out_fmap(xor_out[576*8*8*bW:577*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[592*5*5:593*5*5-1]), .o_out_fmap(xor_out[592*8*8*bW:593*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[608*5*5:609*5*5-1]), .o_out_fmap(xor_out[608*8*8*bW:609*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[624*5*5:625*5*5-1]), .o_out_fmap(xor_out[624*8*8*bW:625*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[640*5*5:641*5*5-1]), .o_out_fmap(xor_out[640*8*8*bW:641*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[656*5*5:657*5*5-1]), .o_out_fmap(xor_out[656*8*8*bW:657*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[672*5*5:673*5*5-1]), .o_out_fmap(xor_out[672*8*8*bW:673*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[688*5*5:689*5*5-1]), .o_out_fmap(xor_out[688*8*8*bW:689*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[704*5*5:705*5*5-1]), .o_out_fmap(xor_out[704*8*8*bW:705*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[720*5*5:721*5*5-1]), .o_out_fmap(xor_out[720*8*8*bW:721*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[736*5*5:737*5*5-1]), .o_out_fmap(xor_out[736*8*8*bW:737*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[752*5*5:753*5*5-1]), .o_out_fmap(xor_out[752*8*8*bW:753*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[768*5*5:769*5*5-1]), .o_out_fmap(xor_out[768*8*8*bW:769*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[784*5*5:785*5*5-1]), .o_out_fmap(xor_out[784*8*8*bW:785*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[800*5*5:801*5*5-1]), .o_out_fmap(xor_out[800*8*8*bW:801*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[816*5*5:817*5*5-1]), .o_out_fmap(xor_out[816*8*8*bW:817*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[832*5*5:833*5*5-1]), .o_out_fmap(xor_out[832*8*8*bW:833*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[848*5*5:849*5*5-1]), .o_out_fmap(xor_out[848*8*8*bW:849*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[864*5*5:865*5*5-1]), .o_out_fmap(xor_out[864*8*8*bW:865*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[880*5*5:881*5*5-1]), .o_out_fmap(xor_out[880*8*8*bW:881*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[896*5*5:897*5*5-1]), .o_out_fmap(xor_out[896*8*8*bW:897*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[912*5*5:913*5*5-1]), .o_out_fmap(xor_out[912*8*8*bW:913*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[928*5*5:929*5*5-1]), .o_out_fmap(xor_out[928*8*8*bW:929*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[944*5*5:945*5*5-1]), .o_out_fmap(xor_out[944*8*8*bW:945*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[17*5*5:18*5*5-1]), .o_out_fmap(xor_out[17*8*8*bW:18*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[34*5*5:35*5*5-1]), .o_out_fmap(xor_out[34*8*8*bW:35*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[51*5*5:52*5*5-1]), .o_out_fmap(xor_out[51*8*8*bW:52*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[68*5*5:69*5*5-1]), .o_out_fmap(xor_out[68*8*8*bW:69*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[85*5*5:86*5*5-1]), .o_out_fmap(xor_out[85*8*8*bW:86*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[102*5*5:103*5*5-1]), .o_out_fmap(xor_out[102*8*8*bW:103*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[119*5*5:120*5*5-1]), .o_out_fmap(xor_out[119*8*8*bW:120*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[136*5*5:137*5*5-1]), .o_out_fmap(xor_out[136*8*8*bW:137*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[153*5*5:154*5*5-1]), .o_out_fmap(xor_out[153*8*8*bW:154*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[170*5*5:171*5*5-1]), .o_out_fmap(xor_out[170*8*8*bW:171*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[187*5*5:188*5*5-1]), .o_out_fmap(xor_out[187*8*8*bW:188*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[204*5*5:205*5*5-1]), .o_out_fmap(xor_out[204*8*8*bW:205*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[221*5*5:222*5*5-1]), .o_out_fmap(xor_out[221*8*8*bW:222*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[238*5*5:239*5*5-1]), .o_out_fmap(xor_out[238*8*8*bW:239*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[255*5*5:256*5*5-1]), .o_out_fmap(xor_out[255*8*8*bW:256*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[272*5*5:273*5*5-1]), .o_out_fmap(xor_out[272*8*8*bW:273*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[289*5*5:290*5*5-1]), .o_out_fmap(xor_out[289*8*8*bW:290*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[306*5*5:307*5*5-1]), .o_out_fmap(xor_out[306*8*8*bW:307*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[323*5*5:324*5*5-1]), .o_out_fmap(xor_out[323*8*8*bW:324*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[340*5*5:341*5*5-1]), .o_out_fmap(xor_out[340*8*8*bW:341*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[357*5*5:358*5*5-1]), .o_out_fmap(xor_out[357*8*8*bW:358*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[374*5*5:375*5*5-1]), .o_out_fmap(xor_out[374*8*8*bW:375*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[391*5*5:392*5*5-1]), .o_out_fmap(xor_out[391*8*8*bW:392*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[408*5*5:409*5*5-1]), .o_out_fmap(xor_out[408*8*8*bW:409*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[425*5*5:426*5*5-1]), .o_out_fmap(xor_out[425*8*8*bW:426*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[442*5*5:443*5*5-1]), .o_out_fmap(xor_out[442*8*8*bW:443*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[459*5*5:460*5*5-1]), .o_out_fmap(xor_out[459*8*8*bW:460*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[476*5*5:477*5*5-1]), .o_out_fmap(xor_out[476*8*8*bW:477*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[493*5*5:494*5*5-1]), .o_out_fmap(xor_out[493*8*8*bW:494*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[510*5*5:511*5*5-1]), .o_out_fmap(xor_out[510*8*8*bW:511*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[527*5*5:528*5*5-1]), .o_out_fmap(xor_out[527*8*8*bW:528*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[544*5*5:545*5*5-1]), .o_out_fmap(xor_out[544*8*8*bW:545*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[561*5*5:562*5*5-1]), .o_out_fmap(xor_out[561*8*8*bW:562*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[578*5*5:579*5*5-1]), .o_out_fmap(xor_out[578*8*8*bW:579*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[595*5*5:596*5*5-1]), .o_out_fmap(xor_out[595*8*8*bW:596*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[612*5*5:613*5*5-1]), .o_out_fmap(xor_out[612*8*8*bW:613*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[629*5*5:630*5*5-1]), .o_out_fmap(xor_out[629*8*8*bW:630*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[646*5*5:647*5*5-1]), .o_out_fmap(xor_out[646*8*8*bW:647*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[663*5*5:664*5*5-1]), .o_out_fmap(xor_out[663*8*8*bW:664*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[680*5*5:681*5*5-1]), .o_out_fmap(xor_out[680*8*8*bW:681*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[697*5*5:698*5*5-1]), .o_out_fmap(xor_out[697*8*8*bW:698*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[714*5*5:715*5*5-1]), .o_out_fmap(xor_out[714*8*8*bW:715*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[731*5*5:732*5*5-1]), .o_out_fmap(xor_out[731*8*8*bW:732*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[748*5*5:749*5*5-1]), .o_out_fmap(xor_out[748*8*8*bW:749*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[765*5*5:766*5*5-1]), .o_out_fmap(xor_out[765*8*8*bW:766*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[782*5*5:783*5*5-1]), .o_out_fmap(xor_out[782*8*8*bW:783*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[799*5*5:800*5*5-1]), .o_out_fmap(xor_out[799*8*8*bW:800*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[816*5*5:817*5*5-1]), .o_out_fmap(xor_out[816*8*8*bW:817*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[833*5*5:834*5*5-1]), .o_out_fmap(xor_out[833*8*8*bW:834*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[850*5*5:851*5*5-1]), .o_out_fmap(xor_out[850*8*8*bW:851*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[867*5*5:868*5*5-1]), .o_out_fmap(xor_out[867*8*8*bW:868*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[884*5*5:885*5*5-1]), .o_out_fmap(xor_out[884*8*8*bW:885*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[901*5*5:902*5*5-1]), .o_out_fmap(xor_out[901*8*8*bW:902*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[918*5*5:919*5*5-1]), .o_out_fmap(xor_out[918*8*8*bW:919*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[935*5*5:936*5*5-1]), .o_out_fmap(xor_out[935*8*8*bW:936*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[952*5*5:953*5*5-1]), .o_out_fmap(xor_out[952*8*8*bW:953*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[969*5*5:970*5*5-1]), .o_out_fmap(xor_out[969*8*8*bW:970*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[986*5*5:987*5*5-1]), .o_out_fmap(xor_out[986*8*8*bW:987*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1003*5*5:1004*5*5-1]), .o_out_fmap(xor_out[1003*8*8*bW:1004*8*8*bW-1]));

endmodule