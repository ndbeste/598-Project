module conv2
    #( parameter bW = 8 )
    (
    input  logic [0:18*12*12 -1]      image         ,
    input  logic [0:18*60*5*5-1]      kernels       ,
    output logic [0:18*60*24*24*bW-1] xor_out 
    );

convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[1*5*5:2*5*5-1]), .o_out_fmap(xor_out[1*24*24*bW:2*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[2*5*5:3*5*5-1]), .o_out_fmap(xor_out[2*24*24*bW:3*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[3*5*5:4*5*5-1]), .o_out_fmap(xor_out[3*24*24*bW:4*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[4*5*5:5*5*5-1]), .o_out_fmap(xor_out[4*24*24*bW:5*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[5*5*5:6*5*5-1]), .o_out_fmap(xor_out[5*24*24*bW:6*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[6*5*5:7*5*5-1]), .o_out_fmap(xor_out[6*24*24*bW:7*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[7*5*5:8*5*5-1]), .o_out_fmap(xor_out[7*24*24*bW:8*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[8*5*5:9*5*5-1]), .o_out_fmap(xor_out[8*24*24*bW:9*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[9*5*5:10*5*5-1]), .o_out_fmap(xor_out[9*24*24*bW:10*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[10*5*5:11*5*5-1]), .o_out_fmap(xor_out[10*24*24*bW:11*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[11*5*5:12*5*5-1]), .o_out_fmap(xor_out[11*24*24*bW:12*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[12*5*5:13*5*5-1]), .o_out_fmap(xor_out[12*24*24*bW:13*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[13*5*5:14*5*5-1]), .o_out_fmap(xor_out[13*24*24*bW:14*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[14*5*5:15*5*5-1]), .o_out_fmap(xor_out[14*24*24*bW:15*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[15*5*5:16*5*5-1]), .o_out_fmap(xor_out[15*24*24*bW:16*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[16*5*5:17*5*5-1]), .o_out_fmap(xor_out[16*24*24*bW:17*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[17*5*5:18*5*5-1]), .o_out_fmap(xor_out[17*24*24*bW:18*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[18*5*5:19*5*5-1]), .o_out_fmap(xor_out[18*24*24*bW:19*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[19*5*5:20*5*5-1]), .o_out_fmap(xor_out[19*24*24*bW:20*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[20*5*5:21*5*5-1]), .o_out_fmap(xor_out[20*24*24*bW:21*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[21*5*5:22*5*5-1]), .o_out_fmap(xor_out[21*24*24*bW:22*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[22*5*5:23*5*5-1]), .o_out_fmap(xor_out[22*24*24*bW:23*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[23*5*5:24*5*5-1]), .o_out_fmap(xor_out[23*24*24*bW:24*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[24*5*5:25*5*5-1]), .o_out_fmap(xor_out[24*24*24*bW:25*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[25*5*5:26*5*5-1]), .o_out_fmap(xor_out[25*24*24*bW:26*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[26*5*5:27*5*5-1]), .o_out_fmap(xor_out[26*24*24*bW:27*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[27*5*5:28*5*5-1]), .o_out_fmap(xor_out[27*24*24*bW:28*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[28*5*5:29*5*5-1]), .o_out_fmap(xor_out[28*24*24*bW:29*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[29*5*5:30*5*5-1]), .o_out_fmap(xor_out[29*24*24*bW:30*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[30*5*5:31*5*5-1]), .o_out_fmap(xor_out[30*24*24*bW:31*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[31*5*5:32*5*5-1]), .o_out_fmap(xor_out[31*24*24*bW:32*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[32*5*5:33*5*5-1]), .o_out_fmap(xor_out[32*24*24*bW:33*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[33*5*5:34*5*5-1]), .o_out_fmap(xor_out[33*24*24*bW:34*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[34*5*5:35*5*5-1]), .o_out_fmap(xor_out[34*24*24*bW:35*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[35*5*5:36*5*5-1]), .o_out_fmap(xor_out[35*24*24*bW:36*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[36*5*5:37*5*5-1]), .o_out_fmap(xor_out[36*24*24*bW:37*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[37*5*5:38*5*5-1]), .o_out_fmap(xor_out[37*24*24*bW:38*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[38*5*5:39*5*5-1]), .o_out_fmap(xor_out[38*24*24*bW:39*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[39*5*5:40*5*5-1]), .o_out_fmap(xor_out[39*24*24*bW:40*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[40*5*5:41*5*5-1]), .o_out_fmap(xor_out[40*24*24*bW:41*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[41*5*5:42*5*5-1]), .o_out_fmap(xor_out[41*24*24*bW:42*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[42*5*5:43*5*5-1]), .o_out_fmap(xor_out[42*24*24*bW:43*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[43*5*5:44*5*5-1]), .o_out_fmap(xor_out[43*24*24*bW:44*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[44*5*5:45*5*5-1]), .o_out_fmap(xor_out[44*24*24*bW:45*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[45*5*5:46*5*5-1]), .o_out_fmap(xor_out[45*24*24*bW:46*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[46*5*5:47*5*5-1]), .o_out_fmap(xor_out[46*24*24*bW:47*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[47*5*5:48*5*5-1]), .o_out_fmap(xor_out[47*24*24*bW:48*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[48*5*5:49*5*5-1]), .o_out_fmap(xor_out[48*24*24*bW:49*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[49*5*5:50*5*5-1]), .o_out_fmap(xor_out[49*24*24*bW:50*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[50*5*5:51*5*5-1]), .o_out_fmap(xor_out[50*24*24*bW:51*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[51*5*5:52*5*5-1]), .o_out_fmap(xor_out[51*24*24*bW:52*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[52*5*5:53*5*5-1]), .o_out_fmap(xor_out[52*24*24*bW:53*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[53*5*5:54*5*5-1]), .o_out_fmap(xor_out[53*24*24*bW:54*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[54*5*5:55*5*5-1]), .o_out_fmap(xor_out[54*24*24*bW:55*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[55*5*5:56*5*5-1]), .o_out_fmap(xor_out[55*24*24*bW:56*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[56*5*5:57*5*5-1]), .o_out_fmap(xor_out[56*24*24*bW:57*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[57*5*5:58*5*5-1]), .o_out_fmap(xor_out[57*24*24*bW:58*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[58*5*5:59*5*5-1]), .o_out_fmap(xor_out[58*24*24*bW:59*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[59*5*5:60*5*5-1]), .o_out_fmap(xor_out[59*24*24*bW:60*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[2*5*5:3*5*5-1]), .o_out_fmap(xor_out[2*24*24*bW:3*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[4*5*5:5*5*5-1]), .o_out_fmap(xor_out[4*24*24*bW:5*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[6*5*5:7*5*5-1]), .o_out_fmap(xor_out[6*24*24*bW:7*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[8*5*5:9*5*5-1]), .o_out_fmap(xor_out[8*24*24*bW:9*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[10*5*5:11*5*5-1]), .o_out_fmap(xor_out[10*24*24*bW:11*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[12*5*5:13*5*5-1]), .o_out_fmap(xor_out[12*24*24*bW:13*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[14*5*5:15*5*5-1]), .o_out_fmap(xor_out[14*24*24*bW:15*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[16*5*5:17*5*5-1]), .o_out_fmap(xor_out[16*24*24*bW:17*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[18*5*5:19*5*5-1]), .o_out_fmap(xor_out[18*24*24*bW:19*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[20*5*5:21*5*5-1]), .o_out_fmap(xor_out[20*24*24*bW:21*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[22*5*5:23*5*5-1]), .o_out_fmap(xor_out[22*24*24*bW:23*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[24*5*5:25*5*5-1]), .o_out_fmap(xor_out[24*24*24*bW:25*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[26*5*5:27*5*5-1]), .o_out_fmap(xor_out[26*24*24*bW:27*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[28*5*5:29*5*5-1]), .o_out_fmap(xor_out[28*24*24*bW:29*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[30*5*5:31*5*5-1]), .o_out_fmap(xor_out[30*24*24*bW:31*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[32*5*5:33*5*5-1]), .o_out_fmap(xor_out[32*24*24*bW:33*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[34*5*5:35*5*5-1]), .o_out_fmap(xor_out[34*24*24*bW:35*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[36*5*5:37*5*5-1]), .o_out_fmap(xor_out[36*24*24*bW:37*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[38*5*5:39*5*5-1]), .o_out_fmap(xor_out[38*24*24*bW:39*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[40*5*5:41*5*5-1]), .o_out_fmap(xor_out[40*24*24*bW:41*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[42*5*5:43*5*5-1]), .o_out_fmap(xor_out[42*24*24*bW:43*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[44*5*5:45*5*5-1]), .o_out_fmap(xor_out[44*24*24*bW:45*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[46*5*5:47*5*5-1]), .o_out_fmap(xor_out[46*24*24*bW:47*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[48*5*5:49*5*5-1]), .o_out_fmap(xor_out[48*24*24*bW:49*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[50*5*5:51*5*5-1]), .o_out_fmap(xor_out[50*24*24*bW:51*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[52*5*5:53*5*5-1]), .o_out_fmap(xor_out[52*24*24*bW:53*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[54*5*5:55*5*5-1]), .o_out_fmap(xor_out[54*24*24*bW:55*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[56*5*5:57*5*5-1]), .o_out_fmap(xor_out[56*24*24*bW:57*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[58*5*5:59*5*5-1]), .o_out_fmap(xor_out[58*24*24*bW:59*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[60*5*5:61*5*5-1]), .o_out_fmap(xor_out[60*24*24*bW:61*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[62*5*5:63*5*5-1]), .o_out_fmap(xor_out[62*24*24*bW:63*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[64*5*5:65*5*5-1]), .o_out_fmap(xor_out[64*24*24*bW:65*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[66*5*5:67*5*5-1]), .o_out_fmap(xor_out[66*24*24*bW:67*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[68*5*5:69*5*5-1]), .o_out_fmap(xor_out[68*24*24*bW:69*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[70*5*5:71*5*5-1]), .o_out_fmap(xor_out[70*24*24*bW:71*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[72*5*5:73*5*5-1]), .o_out_fmap(xor_out[72*24*24*bW:73*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[74*5*5:75*5*5-1]), .o_out_fmap(xor_out[74*24*24*bW:75*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[76*5*5:77*5*5-1]), .o_out_fmap(xor_out[76*24*24*bW:77*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[78*5*5:79*5*5-1]), .o_out_fmap(xor_out[78*24*24*bW:79*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[80*5*5:81*5*5-1]), .o_out_fmap(xor_out[80*24*24*bW:81*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[82*5*5:83*5*5-1]), .o_out_fmap(xor_out[82*24*24*bW:83*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[84*5*5:85*5*5-1]), .o_out_fmap(xor_out[84*24*24*bW:85*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[86*5*5:87*5*5-1]), .o_out_fmap(xor_out[86*24*24*bW:87*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[88*5*5:89*5*5-1]), .o_out_fmap(xor_out[88*24*24*bW:89*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[90*5*5:91*5*5-1]), .o_out_fmap(xor_out[90*24*24*bW:91*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[92*5*5:93*5*5-1]), .o_out_fmap(xor_out[92*24*24*bW:93*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[94*5*5:95*5*5-1]), .o_out_fmap(xor_out[94*24*24*bW:95*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[96*5*5:97*5*5-1]), .o_out_fmap(xor_out[96*24*24*bW:97*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[98*5*5:99*5*5-1]), .o_out_fmap(xor_out[98*24*24*bW:99*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[100*5*5:101*5*5-1]), .o_out_fmap(xor_out[100*24*24*bW:101*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[102*5*5:103*5*5-1]), .o_out_fmap(xor_out[102*24*24*bW:103*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[104*5*5:105*5*5-1]), .o_out_fmap(xor_out[104*24*24*bW:105*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[106*5*5:107*5*5-1]), .o_out_fmap(xor_out[106*24*24*bW:107*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[108*5*5:109*5*5-1]), .o_out_fmap(xor_out[108*24*24*bW:109*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[110*5*5:111*5*5-1]), .o_out_fmap(xor_out[110*24*24*bW:111*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[112*5*5:113*5*5-1]), .o_out_fmap(xor_out[112*24*24*bW:113*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[114*5*5:115*5*5-1]), .o_out_fmap(xor_out[114*24*24*bW:115*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[116*5*5:117*5*5-1]), .o_out_fmap(xor_out[116*24*24*bW:117*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[2*12*12:3*12*12-1]), .i_kernel(kernels[118*5*5:119*5*5-1]), .o_out_fmap(xor_out[118*24*24*bW:119*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[3*5*5:4*5*5-1]), .o_out_fmap(xor_out[3*24*24*bW:4*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[6*5*5:7*5*5-1]), .o_out_fmap(xor_out[6*24*24*bW:7*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[9*5*5:10*5*5-1]), .o_out_fmap(xor_out[9*24*24*bW:10*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[12*5*5:13*5*5-1]), .o_out_fmap(xor_out[12*24*24*bW:13*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[15*5*5:16*5*5-1]), .o_out_fmap(xor_out[15*24*24*bW:16*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[18*5*5:19*5*5-1]), .o_out_fmap(xor_out[18*24*24*bW:19*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[21*5*5:22*5*5-1]), .o_out_fmap(xor_out[21*24*24*bW:22*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[24*5*5:25*5*5-1]), .o_out_fmap(xor_out[24*24*24*bW:25*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[27*5*5:28*5*5-1]), .o_out_fmap(xor_out[27*24*24*bW:28*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[30*5*5:31*5*5-1]), .o_out_fmap(xor_out[30*24*24*bW:31*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[33*5*5:34*5*5-1]), .o_out_fmap(xor_out[33*24*24*bW:34*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[36*5*5:37*5*5-1]), .o_out_fmap(xor_out[36*24*24*bW:37*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[39*5*5:40*5*5-1]), .o_out_fmap(xor_out[39*24*24*bW:40*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[42*5*5:43*5*5-1]), .o_out_fmap(xor_out[42*24*24*bW:43*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[45*5*5:46*5*5-1]), .o_out_fmap(xor_out[45*24*24*bW:46*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[48*5*5:49*5*5-1]), .o_out_fmap(xor_out[48*24*24*bW:49*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[51*5*5:52*5*5-1]), .o_out_fmap(xor_out[51*24*24*bW:52*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[54*5*5:55*5*5-1]), .o_out_fmap(xor_out[54*24*24*bW:55*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[57*5*5:58*5*5-1]), .o_out_fmap(xor_out[57*24*24*bW:58*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[60*5*5:61*5*5-1]), .o_out_fmap(xor_out[60*24*24*bW:61*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[63*5*5:64*5*5-1]), .o_out_fmap(xor_out[63*24*24*bW:64*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[66*5*5:67*5*5-1]), .o_out_fmap(xor_out[66*24*24*bW:67*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[69*5*5:70*5*5-1]), .o_out_fmap(xor_out[69*24*24*bW:70*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[72*5*5:73*5*5-1]), .o_out_fmap(xor_out[72*24*24*bW:73*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[75*5*5:76*5*5-1]), .o_out_fmap(xor_out[75*24*24*bW:76*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[78*5*5:79*5*5-1]), .o_out_fmap(xor_out[78*24*24*bW:79*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[81*5*5:82*5*5-1]), .o_out_fmap(xor_out[81*24*24*bW:82*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[84*5*5:85*5*5-1]), .o_out_fmap(xor_out[84*24*24*bW:85*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[87*5*5:88*5*5-1]), .o_out_fmap(xor_out[87*24*24*bW:88*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[90*5*5:91*5*5-1]), .o_out_fmap(xor_out[90*24*24*bW:91*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[93*5*5:94*5*5-1]), .o_out_fmap(xor_out[93*24*24*bW:94*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[96*5*5:97*5*5-1]), .o_out_fmap(xor_out[96*24*24*bW:97*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[99*5*5:100*5*5-1]), .o_out_fmap(xor_out[99*24*24*bW:100*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[102*5*5:103*5*5-1]), .o_out_fmap(xor_out[102*24*24*bW:103*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[105*5*5:106*5*5-1]), .o_out_fmap(xor_out[105*24*24*bW:106*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[108*5*5:109*5*5-1]), .o_out_fmap(xor_out[108*24*24*bW:109*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[111*5*5:112*5*5-1]), .o_out_fmap(xor_out[111*24*24*bW:112*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[114*5*5:115*5*5-1]), .o_out_fmap(xor_out[114*24*24*bW:115*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[117*5*5:118*5*5-1]), .o_out_fmap(xor_out[117*24*24*bW:118*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[120*5*5:121*5*5-1]), .o_out_fmap(xor_out[120*24*24*bW:121*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[123*5*5:124*5*5-1]), .o_out_fmap(xor_out[123*24*24*bW:124*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[126*5*5:127*5*5-1]), .o_out_fmap(xor_out[126*24*24*bW:127*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[129*5*5:130*5*5-1]), .o_out_fmap(xor_out[129*24*24*bW:130*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[132*5*5:133*5*5-1]), .o_out_fmap(xor_out[132*24*24*bW:133*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[135*5*5:136*5*5-1]), .o_out_fmap(xor_out[135*24*24*bW:136*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[138*5*5:139*5*5-1]), .o_out_fmap(xor_out[138*24*24*bW:139*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[141*5*5:142*5*5-1]), .o_out_fmap(xor_out[141*24*24*bW:142*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[144*5*5:145*5*5-1]), .o_out_fmap(xor_out[144*24*24*bW:145*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[147*5*5:148*5*5-1]), .o_out_fmap(xor_out[147*24*24*bW:148*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[150*5*5:151*5*5-1]), .o_out_fmap(xor_out[150*24*24*bW:151*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[153*5*5:154*5*5-1]), .o_out_fmap(xor_out[153*24*24*bW:154*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[156*5*5:157*5*5-1]), .o_out_fmap(xor_out[156*24*24*bW:157*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[159*5*5:160*5*5-1]), .o_out_fmap(xor_out[159*24*24*bW:160*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[162*5*5:163*5*5-1]), .o_out_fmap(xor_out[162*24*24*bW:163*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[165*5*5:166*5*5-1]), .o_out_fmap(xor_out[165*24*24*bW:166*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[168*5*5:169*5*5-1]), .o_out_fmap(xor_out[168*24*24*bW:169*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[171*5*5:172*5*5-1]), .o_out_fmap(xor_out[171*24*24*bW:172*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[174*5*5:175*5*5-1]), .o_out_fmap(xor_out[174*24*24*bW:175*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[3*12*12:4*12*12-1]), .i_kernel(kernels[177*5*5:178*5*5-1]), .o_out_fmap(xor_out[177*24*24*bW:178*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[4*5*5:5*5*5-1]), .o_out_fmap(xor_out[4*24*24*bW:5*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[8*5*5:9*5*5-1]), .o_out_fmap(xor_out[8*24*24*bW:9*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[12*5*5:13*5*5-1]), .o_out_fmap(xor_out[12*24*24*bW:13*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[16*5*5:17*5*5-1]), .o_out_fmap(xor_out[16*24*24*bW:17*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[20*5*5:21*5*5-1]), .o_out_fmap(xor_out[20*24*24*bW:21*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[24*5*5:25*5*5-1]), .o_out_fmap(xor_out[24*24*24*bW:25*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[28*5*5:29*5*5-1]), .o_out_fmap(xor_out[28*24*24*bW:29*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[32*5*5:33*5*5-1]), .o_out_fmap(xor_out[32*24*24*bW:33*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[36*5*5:37*5*5-1]), .o_out_fmap(xor_out[36*24*24*bW:37*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[40*5*5:41*5*5-1]), .o_out_fmap(xor_out[40*24*24*bW:41*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[44*5*5:45*5*5-1]), .o_out_fmap(xor_out[44*24*24*bW:45*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[48*5*5:49*5*5-1]), .o_out_fmap(xor_out[48*24*24*bW:49*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[52*5*5:53*5*5-1]), .o_out_fmap(xor_out[52*24*24*bW:53*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[56*5*5:57*5*5-1]), .o_out_fmap(xor_out[56*24*24*bW:57*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[60*5*5:61*5*5-1]), .o_out_fmap(xor_out[60*24*24*bW:61*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[64*5*5:65*5*5-1]), .o_out_fmap(xor_out[64*24*24*bW:65*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[68*5*5:69*5*5-1]), .o_out_fmap(xor_out[68*24*24*bW:69*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[72*5*5:73*5*5-1]), .o_out_fmap(xor_out[72*24*24*bW:73*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[76*5*5:77*5*5-1]), .o_out_fmap(xor_out[76*24*24*bW:77*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[80*5*5:81*5*5-1]), .o_out_fmap(xor_out[80*24*24*bW:81*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[84*5*5:85*5*5-1]), .o_out_fmap(xor_out[84*24*24*bW:85*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[88*5*5:89*5*5-1]), .o_out_fmap(xor_out[88*24*24*bW:89*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[92*5*5:93*5*5-1]), .o_out_fmap(xor_out[92*24*24*bW:93*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[96*5*5:97*5*5-1]), .o_out_fmap(xor_out[96*24*24*bW:97*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[100*5*5:101*5*5-1]), .o_out_fmap(xor_out[100*24*24*bW:101*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[104*5*5:105*5*5-1]), .o_out_fmap(xor_out[104*24*24*bW:105*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[108*5*5:109*5*5-1]), .o_out_fmap(xor_out[108*24*24*bW:109*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[112*5*5:113*5*5-1]), .o_out_fmap(xor_out[112*24*24*bW:113*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[116*5*5:117*5*5-1]), .o_out_fmap(xor_out[116*24*24*bW:117*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[120*5*5:121*5*5-1]), .o_out_fmap(xor_out[120*24*24*bW:121*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[124*5*5:125*5*5-1]), .o_out_fmap(xor_out[124*24*24*bW:125*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[128*5*5:129*5*5-1]), .o_out_fmap(xor_out[128*24*24*bW:129*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[132*5*5:133*5*5-1]), .o_out_fmap(xor_out[132*24*24*bW:133*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[136*5*5:137*5*5-1]), .o_out_fmap(xor_out[136*24*24*bW:137*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[140*5*5:141*5*5-1]), .o_out_fmap(xor_out[140*24*24*bW:141*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[144*5*5:145*5*5-1]), .o_out_fmap(xor_out[144*24*24*bW:145*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[148*5*5:149*5*5-1]), .o_out_fmap(xor_out[148*24*24*bW:149*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[152*5*5:153*5*5-1]), .o_out_fmap(xor_out[152*24*24*bW:153*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[156*5*5:157*5*5-1]), .o_out_fmap(xor_out[156*24*24*bW:157*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[160*5*5:161*5*5-1]), .o_out_fmap(xor_out[160*24*24*bW:161*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[164*5*5:165*5*5-1]), .o_out_fmap(xor_out[164*24*24*bW:165*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[168*5*5:169*5*5-1]), .o_out_fmap(xor_out[168*24*24*bW:169*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[172*5*5:173*5*5-1]), .o_out_fmap(xor_out[172*24*24*bW:173*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[176*5*5:177*5*5-1]), .o_out_fmap(xor_out[176*24*24*bW:177*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[180*5*5:181*5*5-1]), .o_out_fmap(xor_out[180*24*24*bW:181*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[184*5*5:185*5*5-1]), .o_out_fmap(xor_out[184*24*24*bW:185*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[188*5*5:189*5*5-1]), .o_out_fmap(xor_out[188*24*24*bW:189*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[192*5*5:193*5*5-1]), .o_out_fmap(xor_out[192*24*24*bW:193*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[196*5*5:197*5*5-1]), .o_out_fmap(xor_out[196*24*24*bW:197*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[200*5*5:201*5*5-1]), .o_out_fmap(xor_out[200*24*24*bW:201*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[204*5*5:205*5*5-1]), .o_out_fmap(xor_out[204*24*24*bW:205*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[208*5*5:209*5*5-1]), .o_out_fmap(xor_out[208*24*24*bW:209*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[212*5*5:213*5*5-1]), .o_out_fmap(xor_out[212*24*24*bW:213*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[216*5*5:217*5*5-1]), .o_out_fmap(xor_out[216*24*24*bW:217*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[220*5*5:221*5*5-1]), .o_out_fmap(xor_out[220*24*24*bW:221*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[224*5*5:225*5*5-1]), .o_out_fmap(xor_out[224*24*24*bW:225*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[228*5*5:229*5*5-1]), .o_out_fmap(xor_out[228*24*24*bW:229*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[232*5*5:233*5*5-1]), .o_out_fmap(xor_out[232*24*24*bW:233*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[4*12*12:5*12*12-1]), .i_kernel(kernels[236*5*5:237*5*5-1]), .o_out_fmap(xor_out[236*24*24*bW:237*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[5*5*5:6*5*5-1]), .o_out_fmap(xor_out[5*24*24*bW:6*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[10*5*5:11*5*5-1]), .o_out_fmap(xor_out[10*24*24*bW:11*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[15*5*5:16*5*5-1]), .o_out_fmap(xor_out[15*24*24*bW:16*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[20*5*5:21*5*5-1]), .o_out_fmap(xor_out[20*24*24*bW:21*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[25*5*5:26*5*5-1]), .o_out_fmap(xor_out[25*24*24*bW:26*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[30*5*5:31*5*5-1]), .o_out_fmap(xor_out[30*24*24*bW:31*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[35*5*5:36*5*5-1]), .o_out_fmap(xor_out[35*24*24*bW:36*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[40*5*5:41*5*5-1]), .o_out_fmap(xor_out[40*24*24*bW:41*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[45*5*5:46*5*5-1]), .o_out_fmap(xor_out[45*24*24*bW:46*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[50*5*5:51*5*5-1]), .o_out_fmap(xor_out[50*24*24*bW:51*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[55*5*5:56*5*5-1]), .o_out_fmap(xor_out[55*24*24*bW:56*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[60*5*5:61*5*5-1]), .o_out_fmap(xor_out[60*24*24*bW:61*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[65*5*5:66*5*5-1]), .o_out_fmap(xor_out[65*24*24*bW:66*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[70*5*5:71*5*5-1]), .o_out_fmap(xor_out[70*24*24*bW:71*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[75*5*5:76*5*5-1]), .o_out_fmap(xor_out[75*24*24*bW:76*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[80*5*5:81*5*5-1]), .o_out_fmap(xor_out[80*24*24*bW:81*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[85*5*5:86*5*5-1]), .o_out_fmap(xor_out[85*24*24*bW:86*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[90*5*5:91*5*5-1]), .o_out_fmap(xor_out[90*24*24*bW:91*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[95*5*5:96*5*5-1]), .o_out_fmap(xor_out[95*24*24*bW:96*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[100*5*5:101*5*5-1]), .o_out_fmap(xor_out[100*24*24*bW:101*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[105*5*5:106*5*5-1]), .o_out_fmap(xor_out[105*24*24*bW:106*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[110*5*5:111*5*5-1]), .o_out_fmap(xor_out[110*24*24*bW:111*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[115*5*5:116*5*5-1]), .o_out_fmap(xor_out[115*24*24*bW:116*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[120*5*5:121*5*5-1]), .o_out_fmap(xor_out[120*24*24*bW:121*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[125*5*5:126*5*5-1]), .o_out_fmap(xor_out[125*24*24*bW:126*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[130*5*5:131*5*5-1]), .o_out_fmap(xor_out[130*24*24*bW:131*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[135*5*5:136*5*5-1]), .o_out_fmap(xor_out[135*24*24*bW:136*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[140*5*5:141*5*5-1]), .o_out_fmap(xor_out[140*24*24*bW:141*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[145*5*5:146*5*5-1]), .o_out_fmap(xor_out[145*24*24*bW:146*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[150*5*5:151*5*5-1]), .o_out_fmap(xor_out[150*24*24*bW:151*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[155*5*5:156*5*5-1]), .o_out_fmap(xor_out[155*24*24*bW:156*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[160*5*5:161*5*5-1]), .o_out_fmap(xor_out[160*24*24*bW:161*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[165*5*5:166*5*5-1]), .o_out_fmap(xor_out[165*24*24*bW:166*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[170*5*5:171*5*5-1]), .o_out_fmap(xor_out[170*24*24*bW:171*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[175*5*5:176*5*5-1]), .o_out_fmap(xor_out[175*24*24*bW:176*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[180*5*5:181*5*5-1]), .o_out_fmap(xor_out[180*24*24*bW:181*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[185*5*5:186*5*5-1]), .o_out_fmap(xor_out[185*24*24*bW:186*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[190*5*5:191*5*5-1]), .o_out_fmap(xor_out[190*24*24*bW:191*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[195*5*5:196*5*5-1]), .o_out_fmap(xor_out[195*24*24*bW:196*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[200*5*5:201*5*5-1]), .o_out_fmap(xor_out[200*24*24*bW:201*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[205*5*5:206*5*5-1]), .o_out_fmap(xor_out[205*24*24*bW:206*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[210*5*5:211*5*5-1]), .o_out_fmap(xor_out[210*24*24*bW:211*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[215*5*5:216*5*5-1]), .o_out_fmap(xor_out[215*24*24*bW:216*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[220*5*5:221*5*5-1]), .o_out_fmap(xor_out[220*24*24*bW:221*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[225*5*5:226*5*5-1]), .o_out_fmap(xor_out[225*24*24*bW:226*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[230*5*5:231*5*5-1]), .o_out_fmap(xor_out[230*24*24*bW:231*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[235*5*5:236*5*5-1]), .o_out_fmap(xor_out[235*24*24*bW:236*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[240*5*5:241*5*5-1]), .o_out_fmap(xor_out[240*24*24*bW:241*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[245*5*5:246*5*5-1]), .o_out_fmap(xor_out[245*24*24*bW:246*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[250*5*5:251*5*5-1]), .o_out_fmap(xor_out[250*24*24*bW:251*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[255*5*5:256*5*5-1]), .o_out_fmap(xor_out[255*24*24*bW:256*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[260*5*5:261*5*5-1]), .o_out_fmap(xor_out[260*24*24*bW:261*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[265*5*5:266*5*5-1]), .o_out_fmap(xor_out[265*24*24*bW:266*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[270*5*5:271*5*5-1]), .o_out_fmap(xor_out[270*24*24*bW:271*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[275*5*5:276*5*5-1]), .o_out_fmap(xor_out[275*24*24*bW:276*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[280*5*5:281*5*5-1]), .o_out_fmap(xor_out[280*24*24*bW:281*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[285*5*5:286*5*5-1]), .o_out_fmap(xor_out[285*24*24*bW:286*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[290*5*5:291*5*5-1]), .o_out_fmap(xor_out[290*24*24*bW:291*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[5*12*12:6*12*12-1]), .i_kernel(kernels[295*5*5:296*5*5-1]), .o_out_fmap(xor_out[295*24*24*bW:296*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[6*5*5:7*5*5-1]), .o_out_fmap(xor_out[6*24*24*bW:7*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[12*5*5:13*5*5-1]), .o_out_fmap(xor_out[12*24*24*bW:13*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[18*5*5:19*5*5-1]), .o_out_fmap(xor_out[18*24*24*bW:19*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[24*5*5:25*5*5-1]), .o_out_fmap(xor_out[24*24*24*bW:25*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[30*5*5:31*5*5-1]), .o_out_fmap(xor_out[30*24*24*bW:31*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[36*5*5:37*5*5-1]), .o_out_fmap(xor_out[36*24*24*bW:37*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[42*5*5:43*5*5-1]), .o_out_fmap(xor_out[42*24*24*bW:43*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[48*5*5:49*5*5-1]), .o_out_fmap(xor_out[48*24*24*bW:49*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[54*5*5:55*5*5-1]), .o_out_fmap(xor_out[54*24*24*bW:55*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[60*5*5:61*5*5-1]), .o_out_fmap(xor_out[60*24*24*bW:61*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[66*5*5:67*5*5-1]), .o_out_fmap(xor_out[66*24*24*bW:67*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[72*5*5:73*5*5-1]), .o_out_fmap(xor_out[72*24*24*bW:73*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[78*5*5:79*5*5-1]), .o_out_fmap(xor_out[78*24*24*bW:79*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[84*5*5:85*5*5-1]), .o_out_fmap(xor_out[84*24*24*bW:85*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[90*5*5:91*5*5-1]), .o_out_fmap(xor_out[90*24*24*bW:91*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[96*5*5:97*5*5-1]), .o_out_fmap(xor_out[96*24*24*bW:97*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[102*5*5:103*5*5-1]), .o_out_fmap(xor_out[102*24*24*bW:103*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[108*5*5:109*5*5-1]), .o_out_fmap(xor_out[108*24*24*bW:109*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[114*5*5:115*5*5-1]), .o_out_fmap(xor_out[114*24*24*bW:115*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[120*5*5:121*5*5-1]), .o_out_fmap(xor_out[120*24*24*bW:121*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[126*5*5:127*5*5-1]), .o_out_fmap(xor_out[126*24*24*bW:127*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[132*5*5:133*5*5-1]), .o_out_fmap(xor_out[132*24*24*bW:133*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[138*5*5:139*5*5-1]), .o_out_fmap(xor_out[138*24*24*bW:139*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[144*5*5:145*5*5-1]), .o_out_fmap(xor_out[144*24*24*bW:145*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[150*5*5:151*5*5-1]), .o_out_fmap(xor_out[150*24*24*bW:151*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[156*5*5:157*5*5-1]), .o_out_fmap(xor_out[156*24*24*bW:157*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[162*5*5:163*5*5-1]), .o_out_fmap(xor_out[162*24*24*bW:163*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[168*5*5:169*5*5-1]), .o_out_fmap(xor_out[168*24*24*bW:169*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[174*5*5:175*5*5-1]), .o_out_fmap(xor_out[174*24*24*bW:175*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[180*5*5:181*5*5-1]), .o_out_fmap(xor_out[180*24*24*bW:181*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[186*5*5:187*5*5-1]), .o_out_fmap(xor_out[186*24*24*bW:187*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[192*5*5:193*5*5-1]), .o_out_fmap(xor_out[192*24*24*bW:193*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[198*5*5:199*5*5-1]), .o_out_fmap(xor_out[198*24*24*bW:199*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[204*5*5:205*5*5-1]), .o_out_fmap(xor_out[204*24*24*bW:205*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[210*5*5:211*5*5-1]), .o_out_fmap(xor_out[210*24*24*bW:211*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[216*5*5:217*5*5-1]), .o_out_fmap(xor_out[216*24*24*bW:217*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[222*5*5:223*5*5-1]), .o_out_fmap(xor_out[222*24*24*bW:223*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[228*5*5:229*5*5-1]), .o_out_fmap(xor_out[228*24*24*bW:229*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[234*5*5:235*5*5-1]), .o_out_fmap(xor_out[234*24*24*bW:235*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[240*5*5:241*5*5-1]), .o_out_fmap(xor_out[240*24*24*bW:241*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[246*5*5:247*5*5-1]), .o_out_fmap(xor_out[246*24*24*bW:247*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[252*5*5:253*5*5-1]), .o_out_fmap(xor_out[252*24*24*bW:253*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[258*5*5:259*5*5-1]), .o_out_fmap(xor_out[258*24*24*bW:259*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[264*5*5:265*5*5-1]), .o_out_fmap(xor_out[264*24*24*bW:265*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[270*5*5:271*5*5-1]), .o_out_fmap(xor_out[270*24*24*bW:271*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[276*5*5:277*5*5-1]), .o_out_fmap(xor_out[276*24*24*bW:277*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[282*5*5:283*5*5-1]), .o_out_fmap(xor_out[282*24*24*bW:283*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[288*5*5:289*5*5-1]), .o_out_fmap(xor_out[288*24*24*bW:289*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[294*5*5:295*5*5-1]), .o_out_fmap(xor_out[294*24*24*bW:295*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[300*5*5:301*5*5-1]), .o_out_fmap(xor_out[300*24*24*bW:301*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[306*5*5:307*5*5-1]), .o_out_fmap(xor_out[306*24*24*bW:307*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[312*5*5:313*5*5-1]), .o_out_fmap(xor_out[312*24*24*bW:313*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[318*5*5:319*5*5-1]), .o_out_fmap(xor_out[318*24*24*bW:319*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[324*5*5:325*5*5-1]), .o_out_fmap(xor_out[324*24*24*bW:325*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[330*5*5:331*5*5-1]), .o_out_fmap(xor_out[330*24*24*bW:331*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[336*5*5:337*5*5-1]), .o_out_fmap(xor_out[336*24*24*bW:337*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[342*5*5:343*5*5-1]), .o_out_fmap(xor_out[342*24*24*bW:343*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[348*5*5:349*5*5-1]), .o_out_fmap(xor_out[348*24*24*bW:349*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[6*12*12:7*12*12-1]), .i_kernel(kernels[354*5*5:355*5*5-1]), .o_out_fmap(xor_out[354*24*24*bW:355*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[7*5*5:8*5*5-1]), .o_out_fmap(xor_out[7*24*24*bW:8*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[14*5*5:15*5*5-1]), .o_out_fmap(xor_out[14*24*24*bW:15*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[21*5*5:22*5*5-1]), .o_out_fmap(xor_out[21*24*24*bW:22*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[28*5*5:29*5*5-1]), .o_out_fmap(xor_out[28*24*24*bW:29*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[35*5*5:36*5*5-1]), .o_out_fmap(xor_out[35*24*24*bW:36*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[42*5*5:43*5*5-1]), .o_out_fmap(xor_out[42*24*24*bW:43*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[49*5*5:50*5*5-1]), .o_out_fmap(xor_out[49*24*24*bW:50*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[56*5*5:57*5*5-1]), .o_out_fmap(xor_out[56*24*24*bW:57*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[63*5*5:64*5*5-1]), .o_out_fmap(xor_out[63*24*24*bW:64*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[70*5*5:71*5*5-1]), .o_out_fmap(xor_out[70*24*24*bW:71*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[77*5*5:78*5*5-1]), .o_out_fmap(xor_out[77*24*24*bW:78*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[84*5*5:85*5*5-1]), .o_out_fmap(xor_out[84*24*24*bW:85*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[91*5*5:92*5*5-1]), .o_out_fmap(xor_out[91*24*24*bW:92*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[98*5*5:99*5*5-1]), .o_out_fmap(xor_out[98*24*24*bW:99*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[105*5*5:106*5*5-1]), .o_out_fmap(xor_out[105*24*24*bW:106*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[112*5*5:113*5*5-1]), .o_out_fmap(xor_out[112*24*24*bW:113*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[119*5*5:120*5*5-1]), .o_out_fmap(xor_out[119*24*24*bW:120*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[126*5*5:127*5*5-1]), .o_out_fmap(xor_out[126*24*24*bW:127*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[133*5*5:134*5*5-1]), .o_out_fmap(xor_out[133*24*24*bW:134*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[140*5*5:141*5*5-1]), .o_out_fmap(xor_out[140*24*24*bW:141*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[147*5*5:148*5*5-1]), .o_out_fmap(xor_out[147*24*24*bW:148*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[154*5*5:155*5*5-1]), .o_out_fmap(xor_out[154*24*24*bW:155*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[161*5*5:162*5*5-1]), .o_out_fmap(xor_out[161*24*24*bW:162*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[168*5*5:169*5*5-1]), .o_out_fmap(xor_out[168*24*24*bW:169*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[175*5*5:176*5*5-1]), .o_out_fmap(xor_out[175*24*24*bW:176*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[182*5*5:183*5*5-1]), .o_out_fmap(xor_out[182*24*24*bW:183*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[189*5*5:190*5*5-1]), .o_out_fmap(xor_out[189*24*24*bW:190*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[196*5*5:197*5*5-1]), .o_out_fmap(xor_out[196*24*24*bW:197*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[203*5*5:204*5*5-1]), .o_out_fmap(xor_out[203*24*24*bW:204*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[210*5*5:211*5*5-1]), .o_out_fmap(xor_out[210*24*24*bW:211*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[217*5*5:218*5*5-1]), .o_out_fmap(xor_out[217*24*24*bW:218*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[224*5*5:225*5*5-1]), .o_out_fmap(xor_out[224*24*24*bW:225*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[231*5*5:232*5*5-1]), .o_out_fmap(xor_out[231*24*24*bW:232*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[238*5*5:239*5*5-1]), .o_out_fmap(xor_out[238*24*24*bW:239*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[245*5*5:246*5*5-1]), .o_out_fmap(xor_out[245*24*24*bW:246*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[252*5*5:253*5*5-1]), .o_out_fmap(xor_out[252*24*24*bW:253*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[259*5*5:260*5*5-1]), .o_out_fmap(xor_out[259*24*24*bW:260*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[266*5*5:267*5*5-1]), .o_out_fmap(xor_out[266*24*24*bW:267*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[273*5*5:274*5*5-1]), .o_out_fmap(xor_out[273*24*24*bW:274*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[280*5*5:281*5*5-1]), .o_out_fmap(xor_out[280*24*24*bW:281*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[287*5*5:288*5*5-1]), .o_out_fmap(xor_out[287*24*24*bW:288*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[294*5*5:295*5*5-1]), .o_out_fmap(xor_out[294*24*24*bW:295*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[301*5*5:302*5*5-1]), .o_out_fmap(xor_out[301*24*24*bW:302*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[308*5*5:309*5*5-1]), .o_out_fmap(xor_out[308*24*24*bW:309*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[315*5*5:316*5*5-1]), .o_out_fmap(xor_out[315*24*24*bW:316*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[322*5*5:323*5*5-1]), .o_out_fmap(xor_out[322*24*24*bW:323*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[329*5*5:330*5*5-1]), .o_out_fmap(xor_out[329*24*24*bW:330*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[336*5*5:337*5*5-1]), .o_out_fmap(xor_out[336*24*24*bW:337*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[343*5*5:344*5*5-1]), .o_out_fmap(xor_out[343*24*24*bW:344*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[350*5*5:351*5*5-1]), .o_out_fmap(xor_out[350*24*24*bW:351*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[357*5*5:358*5*5-1]), .o_out_fmap(xor_out[357*24*24*bW:358*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[364*5*5:365*5*5-1]), .o_out_fmap(xor_out[364*24*24*bW:365*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[371*5*5:372*5*5-1]), .o_out_fmap(xor_out[371*24*24*bW:372*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[378*5*5:379*5*5-1]), .o_out_fmap(xor_out[378*24*24*bW:379*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[385*5*5:386*5*5-1]), .o_out_fmap(xor_out[385*24*24*bW:386*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[392*5*5:393*5*5-1]), .o_out_fmap(xor_out[392*24*24*bW:393*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[399*5*5:400*5*5-1]), .o_out_fmap(xor_out[399*24*24*bW:400*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[406*5*5:407*5*5-1]), .o_out_fmap(xor_out[406*24*24*bW:407*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[7*12*12:8*12*12-1]), .i_kernel(kernels[413*5*5:414*5*5-1]), .o_out_fmap(xor_out[413*24*24*bW:414*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[8*5*5:9*5*5-1]), .o_out_fmap(xor_out[8*24*24*bW:9*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[16*5*5:17*5*5-1]), .o_out_fmap(xor_out[16*24*24*bW:17*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[24*5*5:25*5*5-1]), .o_out_fmap(xor_out[24*24*24*bW:25*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[32*5*5:33*5*5-1]), .o_out_fmap(xor_out[32*24*24*bW:33*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[40*5*5:41*5*5-1]), .o_out_fmap(xor_out[40*24*24*bW:41*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[48*5*5:49*5*5-1]), .o_out_fmap(xor_out[48*24*24*bW:49*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[56*5*5:57*5*5-1]), .o_out_fmap(xor_out[56*24*24*bW:57*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[64*5*5:65*5*5-1]), .o_out_fmap(xor_out[64*24*24*bW:65*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[72*5*5:73*5*5-1]), .o_out_fmap(xor_out[72*24*24*bW:73*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[80*5*5:81*5*5-1]), .o_out_fmap(xor_out[80*24*24*bW:81*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[88*5*5:89*5*5-1]), .o_out_fmap(xor_out[88*24*24*bW:89*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[96*5*5:97*5*5-1]), .o_out_fmap(xor_out[96*24*24*bW:97*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[104*5*5:105*5*5-1]), .o_out_fmap(xor_out[104*24*24*bW:105*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[112*5*5:113*5*5-1]), .o_out_fmap(xor_out[112*24*24*bW:113*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[120*5*5:121*5*5-1]), .o_out_fmap(xor_out[120*24*24*bW:121*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[128*5*5:129*5*5-1]), .o_out_fmap(xor_out[128*24*24*bW:129*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[136*5*5:137*5*5-1]), .o_out_fmap(xor_out[136*24*24*bW:137*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[144*5*5:145*5*5-1]), .o_out_fmap(xor_out[144*24*24*bW:145*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[152*5*5:153*5*5-1]), .o_out_fmap(xor_out[152*24*24*bW:153*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[160*5*5:161*5*5-1]), .o_out_fmap(xor_out[160*24*24*bW:161*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[168*5*5:169*5*5-1]), .o_out_fmap(xor_out[168*24*24*bW:169*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[176*5*5:177*5*5-1]), .o_out_fmap(xor_out[176*24*24*bW:177*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[184*5*5:185*5*5-1]), .o_out_fmap(xor_out[184*24*24*bW:185*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[192*5*5:193*5*5-1]), .o_out_fmap(xor_out[192*24*24*bW:193*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[200*5*5:201*5*5-1]), .o_out_fmap(xor_out[200*24*24*bW:201*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[208*5*5:209*5*5-1]), .o_out_fmap(xor_out[208*24*24*bW:209*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[216*5*5:217*5*5-1]), .o_out_fmap(xor_out[216*24*24*bW:217*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[224*5*5:225*5*5-1]), .o_out_fmap(xor_out[224*24*24*bW:225*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[232*5*5:233*5*5-1]), .o_out_fmap(xor_out[232*24*24*bW:233*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[240*5*5:241*5*5-1]), .o_out_fmap(xor_out[240*24*24*bW:241*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[248*5*5:249*5*5-1]), .o_out_fmap(xor_out[248*24*24*bW:249*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[256*5*5:257*5*5-1]), .o_out_fmap(xor_out[256*24*24*bW:257*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[264*5*5:265*5*5-1]), .o_out_fmap(xor_out[264*24*24*bW:265*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[272*5*5:273*5*5-1]), .o_out_fmap(xor_out[272*24*24*bW:273*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[280*5*5:281*5*5-1]), .o_out_fmap(xor_out[280*24*24*bW:281*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[288*5*5:289*5*5-1]), .o_out_fmap(xor_out[288*24*24*bW:289*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[296*5*5:297*5*5-1]), .o_out_fmap(xor_out[296*24*24*bW:297*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[304*5*5:305*5*5-1]), .o_out_fmap(xor_out[304*24*24*bW:305*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[312*5*5:313*5*5-1]), .o_out_fmap(xor_out[312*24*24*bW:313*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[320*5*5:321*5*5-1]), .o_out_fmap(xor_out[320*24*24*bW:321*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[328*5*5:329*5*5-1]), .o_out_fmap(xor_out[328*24*24*bW:329*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[336*5*5:337*5*5-1]), .o_out_fmap(xor_out[336*24*24*bW:337*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[344*5*5:345*5*5-1]), .o_out_fmap(xor_out[344*24*24*bW:345*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[352*5*5:353*5*5-1]), .o_out_fmap(xor_out[352*24*24*bW:353*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[360*5*5:361*5*5-1]), .o_out_fmap(xor_out[360*24*24*bW:361*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[368*5*5:369*5*5-1]), .o_out_fmap(xor_out[368*24*24*bW:369*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[376*5*5:377*5*5-1]), .o_out_fmap(xor_out[376*24*24*bW:377*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[384*5*5:385*5*5-1]), .o_out_fmap(xor_out[384*24*24*bW:385*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[392*5*5:393*5*5-1]), .o_out_fmap(xor_out[392*24*24*bW:393*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[400*5*5:401*5*5-1]), .o_out_fmap(xor_out[400*24*24*bW:401*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[408*5*5:409*5*5-1]), .o_out_fmap(xor_out[408*24*24*bW:409*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[416*5*5:417*5*5-1]), .o_out_fmap(xor_out[416*24*24*bW:417*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[424*5*5:425*5*5-1]), .o_out_fmap(xor_out[424*24*24*bW:425*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[432*5*5:433*5*5-1]), .o_out_fmap(xor_out[432*24*24*bW:433*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[440*5*5:441*5*5-1]), .o_out_fmap(xor_out[440*24*24*bW:441*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[448*5*5:449*5*5-1]), .o_out_fmap(xor_out[448*24*24*bW:449*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[456*5*5:457*5*5-1]), .o_out_fmap(xor_out[456*24*24*bW:457*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[464*5*5:465*5*5-1]), .o_out_fmap(xor_out[464*24*24*bW:465*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[8*12*12:9*12*12-1]), .i_kernel(kernels[472*5*5:473*5*5-1]), .o_out_fmap(xor_out[472*24*24*bW:473*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[9*5*5:10*5*5-1]), .o_out_fmap(xor_out[9*24*24*bW:10*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[18*5*5:19*5*5-1]), .o_out_fmap(xor_out[18*24*24*bW:19*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[27*5*5:28*5*5-1]), .o_out_fmap(xor_out[27*24*24*bW:28*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[36*5*5:37*5*5-1]), .o_out_fmap(xor_out[36*24*24*bW:37*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[45*5*5:46*5*5-1]), .o_out_fmap(xor_out[45*24*24*bW:46*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[54*5*5:55*5*5-1]), .o_out_fmap(xor_out[54*24*24*bW:55*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[63*5*5:64*5*5-1]), .o_out_fmap(xor_out[63*24*24*bW:64*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[72*5*5:73*5*5-1]), .o_out_fmap(xor_out[72*24*24*bW:73*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[81*5*5:82*5*5-1]), .o_out_fmap(xor_out[81*24*24*bW:82*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[90*5*5:91*5*5-1]), .o_out_fmap(xor_out[90*24*24*bW:91*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[99*5*5:100*5*5-1]), .o_out_fmap(xor_out[99*24*24*bW:100*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[108*5*5:109*5*5-1]), .o_out_fmap(xor_out[108*24*24*bW:109*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[117*5*5:118*5*5-1]), .o_out_fmap(xor_out[117*24*24*bW:118*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[126*5*5:127*5*5-1]), .o_out_fmap(xor_out[126*24*24*bW:127*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[135*5*5:136*5*5-1]), .o_out_fmap(xor_out[135*24*24*bW:136*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[144*5*5:145*5*5-1]), .o_out_fmap(xor_out[144*24*24*bW:145*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[153*5*5:154*5*5-1]), .o_out_fmap(xor_out[153*24*24*bW:154*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[162*5*5:163*5*5-1]), .o_out_fmap(xor_out[162*24*24*bW:163*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[171*5*5:172*5*5-1]), .o_out_fmap(xor_out[171*24*24*bW:172*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[180*5*5:181*5*5-1]), .o_out_fmap(xor_out[180*24*24*bW:181*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[189*5*5:190*5*5-1]), .o_out_fmap(xor_out[189*24*24*bW:190*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[198*5*5:199*5*5-1]), .o_out_fmap(xor_out[198*24*24*bW:199*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[207*5*5:208*5*5-1]), .o_out_fmap(xor_out[207*24*24*bW:208*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[216*5*5:217*5*5-1]), .o_out_fmap(xor_out[216*24*24*bW:217*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[225*5*5:226*5*5-1]), .o_out_fmap(xor_out[225*24*24*bW:226*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[234*5*5:235*5*5-1]), .o_out_fmap(xor_out[234*24*24*bW:235*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[243*5*5:244*5*5-1]), .o_out_fmap(xor_out[243*24*24*bW:244*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[252*5*5:253*5*5-1]), .o_out_fmap(xor_out[252*24*24*bW:253*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[261*5*5:262*5*5-1]), .o_out_fmap(xor_out[261*24*24*bW:262*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[270*5*5:271*5*5-1]), .o_out_fmap(xor_out[270*24*24*bW:271*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[279*5*5:280*5*5-1]), .o_out_fmap(xor_out[279*24*24*bW:280*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[288*5*5:289*5*5-1]), .o_out_fmap(xor_out[288*24*24*bW:289*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[297*5*5:298*5*5-1]), .o_out_fmap(xor_out[297*24*24*bW:298*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[306*5*5:307*5*5-1]), .o_out_fmap(xor_out[306*24*24*bW:307*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[315*5*5:316*5*5-1]), .o_out_fmap(xor_out[315*24*24*bW:316*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[324*5*5:325*5*5-1]), .o_out_fmap(xor_out[324*24*24*bW:325*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[333*5*5:334*5*5-1]), .o_out_fmap(xor_out[333*24*24*bW:334*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[342*5*5:343*5*5-1]), .o_out_fmap(xor_out[342*24*24*bW:343*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[351*5*5:352*5*5-1]), .o_out_fmap(xor_out[351*24*24*bW:352*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[360*5*5:361*5*5-1]), .o_out_fmap(xor_out[360*24*24*bW:361*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[369*5*5:370*5*5-1]), .o_out_fmap(xor_out[369*24*24*bW:370*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[378*5*5:379*5*5-1]), .o_out_fmap(xor_out[378*24*24*bW:379*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[387*5*5:388*5*5-1]), .o_out_fmap(xor_out[387*24*24*bW:388*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[396*5*5:397*5*5-1]), .o_out_fmap(xor_out[396*24*24*bW:397*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[405*5*5:406*5*5-1]), .o_out_fmap(xor_out[405*24*24*bW:406*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[414*5*5:415*5*5-1]), .o_out_fmap(xor_out[414*24*24*bW:415*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[423*5*5:424*5*5-1]), .o_out_fmap(xor_out[423*24*24*bW:424*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[432*5*5:433*5*5-1]), .o_out_fmap(xor_out[432*24*24*bW:433*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[441*5*5:442*5*5-1]), .o_out_fmap(xor_out[441*24*24*bW:442*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[450*5*5:451*5*5-1]), .o_out_fmap(xor_out[450*24*24*bW:451*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[459*5*5:460*5*5-1]), .o_out_fmap(xor_out[459*24*24*bW:460*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[468*5*5:469*5*5-1]), .o_out_fmap(xor_out[468*24*24*bW:469*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[477*5*5:478*5*5-1]), .o_out_fmap(xor_out[477*24*24*bW:478*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[486*5*5:487*5*5-1]), .o_out_fmap(xor_out[486*24*24*bW:487*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[495*5*5:496*5*5-1]), .o_out_fmap(xor_out[495*24*24*bW:496*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[504*5*5:505*5*5-1]), .o_out_fmap(xor_out[504*24*24*bW:505*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[513*5*5:514*5*5-1]), .o_out_fmap(xor_out[513*24*24*bW:514*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[522*5*5:523*5*5-1]), .o_out_fmap(xor_out[522*24*24*bW:523*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[9*12*12:10*12*12-1]), .i_kernel(kernels[531*5*5:532*5*5-1]), .o_out_fmap(xor_out[531*24*24*bW:532*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[10*5*5:11*5*5-1]), .o_out_fmap(xor_out[10*24*24*bW:11*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[20*5*5:21*5*5-1]), .o_out_fmap(xor_out[20*24*24*bW:21*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[30*5*5:31*5*5-1]), .o_out_fmap(xor_out[30*24*24*bW:31*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[40*5*5:41*5*5-1]), .o_out_fmap(xor_out[40*24*24*bW:41*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[50*5*5:51*5*5-1]), .o_out_fmap(xor_out[50*24*24*bW:51*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[60*5*5:61*5*5-1]), .o_out_fmap(xor_out[60*24*24*bW:61*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[70*5*5:71*5*5-1]), .o_out_fmap(xor_out[70*24*24*bW:71*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[80*5*5:81*5*5-1]), .o_out_fmap(xor_out[80*24*24*bW:81*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[90*5*5:91*5*5-1]), .o_out_fmap(xor_out[90*24*24*bW:91*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[100*5*5:101*5*5-1]), .o_out_fmap(xor_out[100*24*24*bW:101*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[110*5*5:111*5*5-1]), .o_out_fmap(xor_out[110*24*24*bW:111*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[120*5*5:121*5*5-1]), .o_out_fmap(xor_out[120*24*24*bW:121*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[130*5*5:131*5*5-1]), .o_out_fmap(xor_out[130*24*24*bW:131*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[140*5*5:141*5*5-1]), .o_out_fmap(xor_out[140*24*24*bW:141*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[150*5*5:151*5*5-1]), .o_out_fmap(xor_out[150*24*24*bW:151*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[160*5*5:161*5*5-1]), .o_out_fmap(xor_out[160*24*24*bW:161*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[170*5*5:171*5*5-1]), .o_out_fmap(xor_out[170*24*24*bW:171*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[180*5*5:181*5*5-1]), .o_out_fmap(xor_out[180*24*24*bW:181*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[190*5*5:191*5*5-1]), .o_out_fmap(xor_out[190*24*24*bW:191*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[200*5*5:201*5*5-1]), .o_out_fmap(xor_out[200*24*24*bW:201*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[210*5*5:211*5*5-1]), .o_out_fmap(xor_out[210*24*24*bW:211*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[220*5*5:221*5*5-1]), .o_out_fmap(xor_out[220*24*24*bW:221*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[230*5*5:231*5*5-1]), .o_out_fmap(xor_out[230*24*24*bW:231*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[240*5*5:241*5*5-1]), .o_out_fmap(xor_out[240*24*24*bW:241*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[250*5*5:251*5*5-1]), .o_out_fmap(xor_out[250*24*24*bW:251*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[260*5*5:261*5*5-1]), .o_out_fmap(xor_out[260*24*24*bW:261*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[270*5*5:271*5*5-1]), .o_out_fmap(xor_out[270*24*24*bW:271*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[280*5*5:281*5*5-1]), .o_out_fmap(xor_out[280*24*24*bW:281*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[290*5*5:291*5*5-1]), .o_out_fmap(xor_out[290*24*24*bW:291*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[300*5*5:301*5*5-1]), .o_out_fmap(xor_out[300*24*24*bW:301*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[310*5*5:311*5*5-1]), .o_out_fmap(xor_out[310*24*24*bW:311*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[320*5*5:321*5*5-1]), .o_out_fmap(xor_out[320*24*24*bW:321*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[330*5*5:331*5*5-1]), .o_out_fmap(xor_out[330*24*24*bW:331*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[340*5*5:341*5*5-1]), .o_out_fmap(xor_out[340*24*24*bW:341*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[350*5*5:351*5*5-1]), .o_out_fmap(xor_out[350*24*24*bW:351*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[360*5*5:361*5*5-1]), .o_out_fmap(xor_out[360*24*24*bW:361*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[370*5*5:371*5*5-1]), .o_out_fmap(xor_out[370*24*24*bW:371*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[380*5*5:381*5*5-1]), .o_out_fmap(xor_out[380*24*24*bW:381*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[390*5*5:391*5*5-1]), .o_out_fmap(xor_out[390*24*24*bW:391*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[400*5*5:401*5*5-1]), .o_out_fmap(xor_out[400*24*24*bW:401*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[410*5*5:411*5*5-1]), .o_out_fmap(xor_out[410*24*24*bW:411*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[420*5*5:421*5*5-1]), .o_out_fmap(xor_out[420*24*24*bW:421*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[430*5*5:431*5*5-1]), .o_out_fmap(xor_out[430*24*24*bW:431*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[440*5*5:441*5*5-1]), .o_out_fmap(xor_out[440*24*24*bW:441*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[450*5*5:451*5*5-1]), .o_out_fmap(xor_out[450*24*24*bW:451*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[460*5*5:461*5*5-1]), .o_out_fmap(xor_out[460*24*24*bW:461*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[470*5*5:471*5*5-1]), .o_out_fmap(xor_out[470*24*24*bW:471*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[480*5*5:481*5*5-1]), .o_out_fmap(xor_out[480*24*24*bW:481*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[490*5*5:491*5*5-1]), .o_out_fmap(xor_out[490*24*24*bW:491*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[500*5*5:501*5*5-1]), .o_out_fmap(xor_out[500*24*24*bW:501*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[510*5*5:511*5*5-1]), .o_out_fmap(xor_out[510*24*24*bW:511*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[520*5*5:521*5*5-1]), .o_out_fmap(xor_out[520*24*24*bW:521*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[530*5*5:531*5*5-1]), .o_out_fmap(xor_out[530*24*24*bW:531*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[540*5*5:541*5*5-1]), .o_out_fmap(xor_out[540*24*24*bW:541*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[550*5*5:551*5*5-1]), .o_out_fmap(xor_out[550*24*24*bW:551*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[560*5*5:561*5*5-1]), .o_out_fmap(xor_out[560*24*24*bW:561*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[570*5*5:571*5*5-1]), .o_out_fmap(xor_out[570*24*24*bW:571*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[580*5*5:581*5*5-1]), .o_out_fmap(xor_out[580*24*24*bW:581*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[10*12*12:11*12*12-1]), .i_kernel(kernels[590*5*5:591*5*5-1]), .o_out_fmap(xor_out[590*24*24*bW:591*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[11*5*5:12*5*5-1]), .o_out_fmap(xor_out[11*24*24*bW:12*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[22*5*5:23*5*5-1]), .o_out_fmap(xor_out[22*24*24*bW:23*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[33*5*5:34*5*5-1]), .o_out_fmap(xor_out[33*24*24*bW:34*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[44*5*5:45*5*5-1]), .o_out_fmap(xor_out[44*24*24*bW:45*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[55*5*5:56*5*5-1]), .o_out_fmap(xor_out[55*24*24*bW:56*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[66*5*5:67*5*5-1]), .o_out_fmap(xor_out[66*24*24*bW:67*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[77*5*5:78*5*5-1]), .o_out_fmap(xor_out[77*24*24*bW:78*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[88*5*5:89*5*5-1]), .o_out_fmap(xor_out[88*24*24*bW:89*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[99*5*5:100*5*5-1]), .o_out_fmap(xor_out[99*24*24*bW:100*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[110*5*5:111*5*5-1]), .o_out_fmap(xor_out[110*24*24*bW:111*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[121*5*5:122*5*5-1]), .o_out_fmap(xor_out[121*24*24*bW:122*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[132*5*5:133*5*5-1]), .o_out_fmap(xor_out[132*24*24*bW:133*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[143*5*5:144*5*5-1]), .o_out_fmap(xor_out[143*24*24*bW:144*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[154*5*5:155*5*5-1]), .o_out_fmap(xor_out[154*24*24*bW:155*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[165*5*5:166*5*5-1]), .o_out_fmap(xor_out[165*24*24*bW:166*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[176*5*5:177*5*5-1]), .o_out_fmap(xor_out[176*24*24*bW:177*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[187*5*5:188*5*5-1]), .o_out_fmap(xor_out[187*24*24*bW:188*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[198*5*5:199*5*5-1]), .o_out_fmap(xor_out[198*24*24*bW:199*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[209*5*5:210*5*5-1]), .o_out_fmap(xor_out[209*24*24*bW:210*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[220*5*5:221*5*5-1]), .o_out_fmap(xor_out[220*24*24*bW:221*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[231*5*5:232*5*5-1]), .o_out_fmap(xor_out[231*24*24*bW:232*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[242*5*5:243*5*5-1]), .o_out_fmap(xor_out[242*24*24*bW:243*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[253*5*5:254*5*5-1]), .o_out_fmap(xor_out[253*24*24*bW:254*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[264*5*5:265*5*5-1]), .o_out_fmap(xor_out[264*24*24*bW:265*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[275*5*5:276*5*5-1]), .o_out_fmap(xor_out[275*24*24*bW:276*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[286*5*5:287*5*5-1]), .o_out_fmap(xor_out[286*24*24*bW:287*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[297*5*5:298*5*5-1]), .o_out_fmap(xor_out[297*24*24*bW:298*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[308*5*5:309*5*5-1]), .o_out_fmap(xor_out[308*24*24*bW:309*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[319*5*5:320*5*5-1]), .o_out_fmap(xor_out[319*24*24*bW:320*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[330*5*5:331*5*5-1]), .o_out_fmap(xor_out[330*24*24*bW:331*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[341*5*5:342*5*5-1]), .o_out_fmap(xor_out[341*24*24*bW:342*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[352*5*5:353*5*5-1]), .o_out_fmap(xor_out[352*24*24*bW:353*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[363*5*5:364*5*5-1]), .o_out_fmap(xor_out[363*24*24*bW:364*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[374*5*5:375*5*5-1]), .o_out_fmap(xor_out[374*24*24*bW:375*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[385*5*5:386*5*5-1]), .o_out_fmap(xor_out[385*24*24*bW:386*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[396*5*5:397*5*5-1]), .o_out_fmap(xor_out[396*24*24*bW:397*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[407*5*5:408*5*5-1]), .o_out_fmap(xor_out[407*24*24*bW:408*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[418*5*5:419*5*5-1]), .o_out_fmap(xor_out[418*24*24*bW:419*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[429*5*5:430*5*5-1]), .o_out_fmap(xor_out[429*24*24*bW:430*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[440*5*5:441*5*5-1]), .o_out_fmap(xor_out[440*24*24*bW:441*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[451*5*5:452*5*5-1]), .o_out_fmap(xor_out[451*24*24*bW:452*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[462*5*5:463*5*5-1]), .o_out_fmap(xor_out[462*24*24*bW:463*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[473*5*5:474*5*5-1]), .o_out_fmap(xor_out[473*24*24*bW:474*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[484*5*5:485*5*5-1]), .o_out_fmap(xor_out[484*24*24*bW:485*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[495*5*5:496*5*5-1]), .o_out_fmap(xor_out[495*24*24*bW:496*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[506*5*5:507*5*5-1]), .o_out_fmap(xor_out[506*24*24*bW:507*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[517*5*5:518*5*5-1]), .o_out_fmap(xor_out[517*24*24*bW:518*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[528*5*5:529*5*5-1]), .o_out_fmap(xor_out[528*24*24*bW:529*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[539*5*5:540*5*5-1]), .o_out_fmap(xor_out[539*24*24*bW:540*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[550*5*5:551*5*5-1]), .o_out_fmap(xor_out[550*24*24*bW:551*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[561*5*5:562*5*5-1]), .o_out_fmap(xor_out[561*24*24*bW:562*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[572*5*5:573*5*5-1]), .o_out_fmap(xor_out[572*24*24*bW:573*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[583*5*5:584*5*5-1]), .o_out_fmap(xor_out[583*24*24*bW:584*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[594*5*5:595*5*5-1]), .o_out_fmap(xor_out[594*24*24*bW:595*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[605*5*5:606*5*5-1]), .o_out_fmap(xor_out[605*24*24*bW:606*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[616*5*5:617*5*5-1]), .o_out_fmap(xor_out[616*24*24*bW:617*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[627*5*5:628*5*5-1]), .o_out_fmap(xor_out[627*24*24*bW:628*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[638*5*5:639*5*5-1]), .o_out_fmap(xor_out[638*24*24*bW:639*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[11*12*12:12*12*12-1]), .i_kernel(kernels[649*5*5:650*5*5-1]), .o_out_fmap(xor_out[649*24*24*bW:650*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[12*5*5:13*5*5-1]), .o_out_fmap(xor_out[12*24*24*bW:13*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[24*5*5:25*5*5-1]), .o_out_fmap(xor_out[24*24*24*bW:25*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[36*5*5:37*5*5-1]), .o_out_fmap(xor_out[36*24*24*bW:37*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[48*5*5:49*5*5-1]), .o_out_fmap(xor_out[48*24*24*bW:49*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[60*5*5:61*5*5-1]), .o_out_fmap(xor_out[60*24*24*bW:61*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[72*5*5:73*5*5-1]), .o_out_fmap(xor_out[72*24*24*bW:73*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[84*5*5:85*5*5-1]), .o_out_fmap(xor_out[84*24*24*bW:85*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[96*5*5:97*5*5-1]), .o_out_fmap(xor_out[96*24*24*bW:97*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[108*5*5:109*5*5-1]), .o_out_fmap(xor_out[108*24*24*bW:109*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[120*5*5:121*5*5-1]), .o_out_fmap(xor_out[120*24*24*bW:121*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[132*5*5:133*5*5-1]), .o_out_fmap(xor_out[132*24*24*bW:133*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[144*5*5:145*5*5-1]), .o_out_fmap(xor_out[144*24*24*bW:145*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[156*5*5:157*5*5-1]), .o_out_fmap(xor_out[156*24*24*bW:157*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[168*5*5:169*5*5-1]), .o_out_fmap(xor_out[168*24*24*bW:169*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[180*5*5:181*5*5-1]), .o_out_fmap(xor_out[180*24*24*bW:181*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[192*5*5:193*5*5-1]), .o_out_fmap(xor_out[192*24*24*bW:193*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[204*5*5:205*5*5-1]), .o_out_fmap(xor_out[204*24*24*bW:205*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[216*5*5:217*5*5-1]), .o_out_fmap(xor_out[216*24*24*bW:217*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[228*5*5:229*5*5-1]), .o_out_fmap(xor_out[228*24*24*bW:229*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[240*5*5:241*5*5-1]), .o_out_fmap(xor_out[240*24*24*bW:241*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[252*5*5:253*5*5-1]), .o_out_fmap(xor_out[252*24*24*bW:253*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[264*5*5:265*5*5-1]), .o_out_fmap(xor_out[264*24*24*bW:265*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[276*5*5:277*5*5-1]), .o_out_fmap(xor_out[276*24*24*bW:277*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[288*5*5:289*5*5-1]), .o_out_fmap(xor_out[288*24*24*bW:289*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[300*5*5:301*5*5-1]), .o_out_fmap(xor_out[300*24*24*bW:301*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[312*5*5:313*5*5-1]), .o_out_fmap(xor_out[312*24*24*bW:313*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[324*5*5:325*5*5-1]), .o_out_fmap(xor_out[324*24*24*bW:325*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[336*5*5:337*5*5-1]), .o_out_fmap(xor_out[336*24*24*bW:337*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[348*5*5:349*5*5-1]), .o_out_fmap(xor_out[348*24*24*bW:349*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[360*5*5:361*5*5-1]), .o_out_fmap(xor_out[360*24*24*bW:361*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[372*5*5:373*5*5-1]), .o_out_fmap(xor_out[372*24*24*bW:373*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[384*5*5:385*5*5-1]), .o_out_fmap(xor_out[384*24*24*bW:385*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[396*5*5:397*5*5-1]), .o_out_fmap(xor_out[396*24*24*bW:397*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[408*5*5:409*5*5-1]), .o_out_fmap(xor_out[408*24*24*bW:409*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[420*5*5:421*5*5-1]), .o_out_fmap(xor_out[420*24*24*bW:421*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[432*5*5:433*5*5-1]), .o_out_fmap(xor_out[432*24*24*bW:433*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[444*5*5:445*5*5-1]), .o_out_fmap(xor_out[444*24*24*bW:445*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[456*5*5:457*5*5-1]), .o_out_fmap(xor_out[456*24*24*bW:457*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[468*5*5:469*5*5-1]), .o_out_fmap(xor_out[468*24*24*bW:469*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[480*5*5:481*5*5-1]), .o_out_fmap(xor_out[480*24*24*bW:481*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[492*5*5:493*5*5-1]), .o_out_fmap(xor_out[492*24*24*bW:493*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[504*5*5:505*5*5-1]), .o_out_fmap(xor_out[504*24*24*bW:505*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[516*5*5:517*5*5-1]), .o_out_fmap(xor_out[516*24*24*bW:517*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[528*5*5:529*5*5-1]), .o_out_fmap(xor_out[528*24*24*bW:529*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[540*5*5:541*5*5-1]), .o_out_fmap(xor_out[540*24*24*bW:541*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[552*5*5:553*5*5-1]), .o_out_fmap(xor_out[552*24*24*bW:553*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[564*5*5:565*5*5-1]), .o_out_fmap(xor_out[564*24*24*bW:565*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[576*5*5:577*5*5-1]), .o_out_fmap(xor_out[576*24*24*bW:577*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[588*5*5:589*5*5-1]), .o_out_fmap(xor_out[588*24*24*bW:589*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[600*5*5:601*5*5-1]), .o_out_fmap(xor_out[600*24*24*bW:601*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[612*5*5:613*5*5-1]), .o_out_fmap(xor_out[612*24*24*bW:613*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[624*5*5:625*5*5-1]), .o_out_fmap(xor_out[624*24*24*bW:625*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[636*5*5:637*5*5-1]), .o_out_fmap(xor_out[636*24*24*bW:637*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[648*5*5:649*5*5-1]), .o_out_fmap(xor_out[648*24*24*bW:649*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[660*5*5:661*5*5-1]), .o_out_fmap(xor_out[660*24*24*bW:661*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[672*5*5:673*5*5-1]), .o_out_fmap(xor_out[672*24*24*bW:673*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[684*5*5:685*5*5-1]), .o_out_fmap(xor_out[684*24*24*bW:685*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[696*5*5:697*5*5-1]), .o_out_fmap(xor_out[696*24*24*bW:697*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[12*12*12:13*12*12-1]), .i_kernel(kernels[708*5*5:709*5*5-1]), .o_out_fmap(xor_out[708*24*24*bW:709*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[13*5*5:14*5*5-1]), .o_out_fmap(xor_out[13*24*24*bW:14*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[26*5*5:27*5*5-1]), .o_out_fmap(xor_out[26*24*24*bW:27*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[39*5*5:40*5*5-1]), .o_out_fmap(xor_out[39*24*24*bW:40*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[52*5*5:53*5*5-1]), .o_out_fmap(xor_out[52*24*24*bW:53*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[65*5*5:66*5*5-1]), .o_out_fmap(xor_out[65*24*24*bW:66*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[78*5*5:79*5*5-1]), .o_out_fmap(xor_out[78*24*24*bW:79*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[91*5*5:92*5*5-1]), .o_out_fmap(xor_out[91*24*24*bW:92*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[104*5*5:105*5*5-1]), .o_out_fmap(xor_out[104*24*24*bW:105*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[117*5*5:118*5*5-1]), .o_out_fmap(xor_out[117*24*24*bW:118*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[130*5*5:131*5*5-1]), .o_out_fmap(xor_out[130*24*24*bW:131*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[143*5*5:144*5*5-1]), .o_out_fmap(xor_out[143*24*24*bW:144*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[156*5*5:157*5*5-1]), .o_out_fmap(xor_out[156*24*24*bW:157*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[169*5*5:170*5*5-1]), .o_out_fmap(xor_out[169*24*24*bW:170*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[182*5*5:183*5*5-1]), .o_out_fmap(xor_out[182*24*24*bW:183*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[195*5*5:196*5*5-1]), .o_out_fmap(xor_out[195*24*24*bW:196*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[208*5*5:209*5*5-1]), .o_out_fmap(xor_out[208*24*24*bW:209*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[221*5*5:222*5*5-1]), .o_out_fmap(xor_out[221*24*24*bW:222*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[234*5*5:235*5*5-1]), .o_out_fmap(xor_out[234*24*24*bW:235*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[247*5*5:248*5*5-1]), .o_out_fmap(xor_out[247*24*24*bW:248*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[260*5*5:261*5*5-1]), .o_out_fmap(xor_out[260*24*24*bW:261*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[273*5*5:274*5*5-1]), .o_out_fmap(xor_out[273*24*24*bW:274*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[286*5*5:287*5*5-1]), .o_out_fmap(xor_out[286*24*24*bW:287*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[299*5*5:300*5*5-1]), .o_out_fmap(xor_out[299*24*24*bW:300*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[312*5*5:313*5*5-1]), .o_out_fmap(xor_out[312*24*24*bW:313*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[325*5*5:326*5*5-1]), .o_out_fmap(xor_out[325*24*24*bW:326*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[338*5*5:339*5*5-1]), .o_out_fmap(xor_out[338*24*24*bW:339*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[351*5*5:352*5*5-1]), .o_out_fmap(xor_out[351*24*24*bW:352*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[364*5*5:365*5*5-1]), .o_out_fmap(xor_out[364*24*24*bW:365*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[377*5*5:378*5*5-1]), .o_out_fmap(xor_out[377*24*24*bW:378*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[390*5*5:391*5*5-1]), .o_out_fmap(xor_out[390*24*24*bW:391*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[403*5*5:404*5*5-1]), .o_out_fmap(xor_out[403*24*24*bW:404*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[416*5*5:417*5*5-1]), .o_out_fmap(xor_out[416*24*24*bW:417*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[429*5*5:430*5*5-1]), .o_out_fmap(xor_out[429*24*24*bW:430*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[442*5*5:443*5*5-1]), .o_out_fmap(xor_out[442*24*24*bW:443*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[455*5*5:456*5*5-1]), .o_out_fmap(xor_out[455*24*24*bW:456*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[468*5*5:469*5*5-1]), .o_out_fmap(xor_out[468*24*24*bW:469*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[481*5*5:482*5*5-1]), .o_out_fmap(xor_out[481*24*24*bW:482*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[494*5*5:495*5*5-1]), .o_out_fmap(xor_out[494*24*24*bW:495*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[507*5*5:508*5*5-1]), .o_out_fmap(xor_out[507*24*24*bW:508*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[520*5*5:521*5*5-1]), .o_out_fmap(xor_out[520*24*24*bW:521*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[533*5*5:534*5*5-1]), .o_out_fmap(xor_out[533*24*24*bW:534*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[546*5*5:547*5*5-1]), .o_out_fmap(xor_out[546*24*24*bW:547*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[559*5*5:560*5*5-1]), .o_out_fmap(xor_out[559*24*24*bW:560*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[572*5*5:573*5*5-1]), .o_out_fmap(xor_out[572*24*24*bW:573*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[585*5*5:586*5*5-1]), .o_out_fmap(xor_out[585*24*24*bW:586*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[598*5*5:599*5*5-1]), .o_out_fmap(xor_out[598*24*24*bW:599*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[611*5*5:612*5*5-1]), .o_out_fmap(xor_out[611*24*24*bW:612*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[624*5*5:625*5*5-1]), .o_out_fmap(xor_out[624*24*24*bW:625*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[637*5*5:638*5*5-1]), .o_out_fmap(xor_out[637*24*24*bW:638*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[650*5*5:651*5*5-1]), .o_out_fmap(xor_out[650*24*24*bW:651*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[663*5*5:664*5*5-1]), .o_out_fmap(xor_out[663*24*24*bW:664*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[676*5*5:677*5*5-1]), .o_out_fmap(xor_out[676*24*24*bW:677*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[689*5*5:690*5*5-1]), .o_out_fmap(xor_out[689*24*24*bW:690*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[702*5*5:703*5*5-1]), .o_out_fmap(xor_out[702*24*24*bW:703*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[715*5*5:716*5*5-1]), .o_out_fmap(xor_out[715*24*24*bW:716*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[728*5*5:729*5*5-1]), .o_out_fmap(xor_out[728*24*24*bW:729*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[741*5*5:742*5*5-1]), .o_out_fmap(xor_out[741*24*24*bW:742*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[754*5*5:755*5*5-1]), .o_out_fmap(xor_out[754*24*24*bW:755*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[13*12*12:14*12*12-1]), .i_kernel(kernels[767*5*5:768*5*5-1]), .o_out_fmap(xor_out[767*24*24*bW:768*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[14*5*5:15*5*5-1]), .o_out_fmap(xor_out[14*24*24*bW:15*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[28*5*5:29*5*5-1]), .o_out_fmap(xor_out[28*24*24*bW:29*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[42*5*5:43*5*5-1]), .o_out_fmap(xor_out[42*24*24*bW:43*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[56*5*5:57*5*5-1]), .o_out_fmap(xor_out[56*24*24*bW:57*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[70*5*5:71*5*5-1]), .o_out_fmap(xor_out[70*24*24*bW:71*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[84*5*5:85*5*5-1]), .o_out_fmap(xor_out[84*24*24*bW:85*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[98*5*5:99*5*5-1]), .o_out_fmap(xor_out[98*24*24*bW:99*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[112*5*5:113*5*5-1]), .o_out_fmap(xor_out[112*24*24*bW:113*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[126*5*5:127*5*5-1]), .o_out_fmap(xor_out[126*24*24*bW:127*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[140*5*5:141*5*5-1]), .o_out_fmap(xor_out[140*24*24*bW:141*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[154*5*5:155*5*5-1]), .o_out_fmap(xor_out[154*24*24*bW:155*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[168*5*5:169*5*5-1]), .o_out_fmap(xor_out[168*24*24*bW:169*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[182*5*5:183*5*5-1]), .o_out_fmap(xor_out[182*24*24*bW:183*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[196*5*5:197*5*5-1]), .o_out_fmap(xor_out[196*24*24*bW:197*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[210*5*5:211*5*5-1]), .o_out_fmap(xor_out[210*24*24*bW:211*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[224*5*5:225*5*5-1]), .o_out_fmap(xor_out[224*24*24*bW:225*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[238*5*5:239*5*5-1]), .o_out_fmap(xor_out[238*24*24*bW:239*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[252*5*5:253*5*5-1]), .o_out_fmap(xor_out[252*24*24*bW:253*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[266*5*5:267*5*5-1]), .o_out_fmap(xor_out[266*24*24*bW:267*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[280*5*5:281*5*5-1]), .o_out_fmap(xor_out[280*24*24*bW:281*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[294*5*5:295*5*5-1]), .o_out_fmap(xor_out[294*24*24*bW:295*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[308*5*5:309*5*5-1]), .o_out_fmap(xor_out[308*24*24*bW:309*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[322*5*5:323*5*5-1]), .o_out_fmap(xor_out[322*24*24*bW:323*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[336*5*5:337*5*5-1]), .o_out_fmap(xor_out[336*24*24*bW:337*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[350*5*5:351*5*5-1]), .o_out_fmap(xor_out[350*24*24*bW:351*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[364*5*5:365*5*5-1]), .o_out_fmap(xor_out[364*24*24*bW:365*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[378*5*5:379*5*5-1]), .o_out_fmap(xor_out[378*24*24*bW:379*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[392*5*5:393*5*5-1]), .o_out_fmap(xor_out[392*24*24*bW:393*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[406*5*5:407*5*5-1]), .o_out_fmap(xor_out[406*24*24*bW:407*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[420*5*5:421*5*5-1]), .o_out_fmap(xor_out[420*24*24*bW:421*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[434*5*5:435*5*5-1]), .o_out_fmap(xor_out[434*24*24*bW:435*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[448*5*5:449*5*5-1]), .o_out_fmap(xor_out[448*24*24*bW:449*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[462*5*5:463*5*5-1]), .o_out_fmap(xor_out[462*24*24*bW:463*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[476*5*5:477*5*5-1]), .o_out_fmap(xor_out[476*24*24*bW:477*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[490*5*5:491*5*5-1]), .o_out_fmap(xor_out[490*24*24*bW:491*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[504*5*5:505*5*5-1]), .o_out_fmap(xor_out[504*24*24*bW:505*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[518*5*5:519*5*5-1]), .o_out_fmap(xor_out[518*24*24*bW:519*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[532*5*5:533*5*5-1]), .o_out_fmap(xor_out[532*24*24*bW:533*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[546*5*5:547*5*5-1]), .o_out_fmap(xor_out[546*24*24*bW:547*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[560*5*5:561*5*5-1]), .o_out_fmap(xor_out[560*24*24*bW:561*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[574*5*5:575*5*5-1]), .o_out_fmap(xor_out[574*24*24*bW:575*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[588*5*5:589*5*5-1]), .o_out_fmap(xor_out[588*24*24*bW:589*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[602*5*5:603*5*5-1]), .o_out_fmap(xor_out[602*24*24*bW:603*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[616*5*5:617*5*5-1]), .o_out_fmap(xor_out[616*24*24*bW:617*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[630*5*5:631*5*5-1]), .o_out_fmap(xor_out[630*24*24*bW:631*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[644*5*5:645*5*5-1]), .o_out_fmap(xor_out[644*24*24*bW:645*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[658*5*5:659*5*5-1]), .o_out_fmap(xor_out[658*24*24*bW:659*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[672*5*5:673*5*5-1]), .o_out_fmap(xor_out[672*24*24*bW:673*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[686*5*5:687*5*5-1]), .o_out_fmap(xor_out[686*24*24*bW:687*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[700*5*5:701*5*5-1]), .o_out_fmap(xor_out[700*24*24*bW:701*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[714*5*5:715*5*5-1]), .o_out_fmap(xor_out[714*24*24*bW:715*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[728*5*5:729*5*5-1]), .o_out_fmap(xor_out[728*24*24*bW:729*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[742*5*5:743*5*5-1]), .o_out_fmap(xor_out[742*24*24*bW:743*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[756*5*5:757*5*5-1]), .o_out_fmap(xor_out[756*24*24*bW:757*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[770*5*5:771*5*5-1]), .o_out_fmap(xor_out[770*24*24*bW:771*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[784*5*5:785*5*5-1]), .o_out_fmap(xor_out[784*24*24*bW:785*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[798*5*5:799*5*5-1]), .o_out_fmap(xor_out[798*24*24*bW:799*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[812*5*5:813*5*5-1]), .o_out_fmap(xor_out[812*24*24*bW:813*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[14*12*12:15*12*12-1]), .i_kernel(kernels[826*5*5:827*5*5-1]), .o_out_fmap(xor_out[826*24*24*bW:827*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[15*5*5:16*5*5-1]), .o_out_fmap(xor_out[15*24*24*bW:16*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[30*5*5:31*5*5-1]), .o_out_fmap(xor_out[30*24*24*bW:31*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[45*5*5:46*5*5-1]), .o_out_fmap(xor_out[45*24*24*bW:46*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[60*5*5:61*5*5-1]), .o_out_fmap(xor_out[60*24*24*bW:61*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[75*5*5:76*5*5-1]), .o_out_fmap(xor_out[75*24*24*bW:76*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[90*5*5:91*5*5-1]), .o_out_fmap(xor_out[90*24*24*bW:91*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[105*5*5:106*5*5-1]), .o_out_fmap(xor_out[105*24*24*bW:106*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[120*5*5:121*5*5-1]), .o_out_fmap(xor_out[120*24*24*bW:121*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[135*5*5:136*5*5-1]), .o_out_fmap(xor_out[135*24*24*bW:136*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[150*5*5:151*5*5-1]), .o_out_fmap(xor_out[150*24*24*bW:151*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[165*5*5:166*5*5-1]), .o_out_fmap(xor_out[165*24*24*bW:166*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[180*5*5:181*5*5-1]), .o_out_fmap(xor_out[180*24*24*bW:181*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[195*5*5:196*5*5-1]), .o_out_fmap(xor_out[195*24*24*bW:196*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[210*5*5:211*5*5-1]), .o_out_fmap(xor_out[210*24*24*bW:211*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[225*5*5:226*5*5-1]), .o_out_fmap(xor_out[225*24*24*bW:226*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[240*5*5:241*5*5-1]), .o_out_fmap(xor_out[240*24*24*bW:241*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[255*5*5:256*5*5-1]), .o_out_fmap(xor_out[255*24*24*bW:256*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[270*5*5:271*5*5-1]), .o_out_fmap(xor_out[270*24*24*bW:271*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[285*5*5:286*5*5-1]), .o_out_fmap(xor_out[285*24*24*bW:286*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[300*5*5:301*5*5-1]), .o_out_fmap(xor_out[300*24*24*bW:301*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[315*5*5:316*5*5-1]), .o_out_fmap(xor_out[315*24*24*bW:316*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[330*5*5:331*5*5-1]), .o_out_fmap(xor_out[330*24*24*bW:331*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[345*5*5:346*5*5-1]), .o_out_fmap(xor_out[345*24*24*bW:346*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[360*5*5:361*5*5-1]), .o_out_fmap(xor_out[360*24*24*bW:361*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[375*5*5:376*5*5-1]), .o_out_fmap(xor_out[375*24*24*bW:376*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[390*5*5:391*5*5-1]), .o_out_fmap(xor_out[390*24*24*bW:391*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[405*5*5:406*5*5-1]), .o_out_fmap(xor_out[405*24*24*bW:406*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[420*5*5:421*5*5-1]), .o_out_fmap(xor_out[420*24*24*bW:421*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[435*5*5:436*5*5-1]), .o_out_fmap(xor_out[435*24*24*bW:436*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[450*5*5:451*5*5-1]), .o_out_fmap(xor_out[450*24*24*bW:451*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[465*5*5:466*5*5-1]), .o_out_fmap(xor_out[465*24*24*bW:466*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[480*5*5:481*5*5-1]), .o_out_fmap(xor_out[480*24*24*bW:481*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[495*5*5:496*5*5-1]), .o_out_fmap(xor_out[495*24*24*bW:496*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[510*5*5:511*5*5-1]), .o_out_fmap(xor_out[510*24*24*bW:511*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[525*5*5:526*5*5-1]), .o_out_fmap(xor_out[525*24*24*bW:526*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[540*5*5:541*5*5-1]), .o_out_fmap(xor_out[540*24*24*bW:541*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[555*5*5:556*5*5-1]), .o_out_fmap(xor_out[555*24*24*bW:556*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[570*5*5:571*5*5-1]), .o_out_fmap(xor_out[570*24*24*bW:571*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[585*5*5:586*5*5-1]), .o_out_fmap(xor_out[585*24*24*bW:586*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[600*5*5:601*5*5-1]), .o_out_fmap(xor_out[600*24*24*bW:601*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[615*5*5:616*5*5-1]), .o_out_fmap(xor_out[615*24*24*bW:616*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[630*5*5:631*5*5-1]), .o_out_fmap(xor_out[630*24*24*bW:631*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[645*5*5:646*5*5-1]), .o_out_fmap(xor_out[645*24*24*bW:646*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[660*5*5:661*5*5-1]), .o_out_fmap(xor_out[660*24*24*bW:661*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[675*5*5:676*5*5-1]), .o_out_fmap(xor_out[675*24*24*bW:676*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[690*5*5:691*5*5-1]), .o_out_fmap(xor_out[690*24*24*bW:691*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[705*5*5:706*5*5-1]), .o_out_fmap(xor_out[705*24*24*bW:706*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[720*5*5:721*5*5-1]), .o_out_fmap(xor_out[720*24*24*bW:721*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[735*5*5:736*5*5-1]), .o_out_fmap(xor_out[735*24*24*bW:736*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[750*5*5:751*5*5-1]), .o_out_fmap(xor_out[750*24*24*bW:751*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[765*5*5:766*5*5-1]), .o_out_fmap(xor_out[765*24*24*bW:766*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[780*5*5:781*5*5-1]), .o_out_fmap(xor_out[780*24*24*bW:781*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[795*5*5:796*5*5-1]), .o_out_fmap(xor_out[795*24*24*bW:796*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[810*5*5:811*5*5-1]), .o_out_fmap(xor_out[810*24*24*bW:811*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[825*5*5:826*5*5-1]), .o_out_fmap(xor_out[825*24*24*bW:826*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[840*5*5:841*5*5-1]), .o_out_fmap(xor_out[840*24*24*bW:841*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[855*5*5:856*5*5-1]), .o_out_fmap(xor_out[855*24*24*bW:856*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[870*5*5:871*5*5-1]), .o_out_fmap(xor_out[870*24*24*bW:871*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[15*12*12:16*12*12-1]), .i_kernel(kernels[885*5*5:886*5*5-1]), .o_out_fmap(xor_out[885*24*24*bW:886*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[16*5*5:17*5*5-1]), .o_out_fmap(xor_out[16*24*24*bW:17*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[32*5*5:33*5*5-1]), .o_out_fmap(xor_out[32*24*24*bW:33*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[48*5*5:49*5*5-1]), .o_out_fmap(xor_out[48*24*24*bW:49*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[64*5*5:65*5*5-1]), .o_out_fmap(xor_out[64*24*24*bW:65*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[80*5*5:81*5*5-1]), .o_out_fmap(xor_out[80*24*24*bW:81*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[96*5*5:97*5*5-1]), .o_out_fmap(xor_out[96*24*24*bW:97*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[112*5*5:113*5*5-1]), .o_out_fmap(xor_out[112*24*24*bW:113*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[128*5*5:129*5*5-1]), .o_out_fmap(xor_out[128*24*24*bW:129*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[144*5*5:145*5*5-1]), .o_out_fmap(xor_out[144*24*24*bW:145*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[160*5*5:161*5*5-1]), .o_out_fmap(xor_out[160*24*24*bW:161*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[176*5*5:177*5*5-1]), .o_out_fmap(xor_out[176*24*24*bW:177*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[192*5*5:193*5*5-1]), .o_out_fmap(xor_out[192*24*24*bW:193*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[208*5*5:209*5*5-1]), .o_out_fmap(xor_out[208*24*24*bW:209*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[224*5*5:225*5*5-1]), .o_out_fmap(xor_out[224*24*24*bW:225*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[240*5*5:241*5*5-1]), .o_out_fmap(xor_out[240*24*24*bW:241*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[256*5*5:257*5*5-1]), .o_out_fmap(xor_out[256*24*24*bW:257*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[272*5*5:273*5*5-1]), .o_out_fmap(xor_out[272*24*24*bW:273*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[288*5*5:289*5*5-1]), .o_out_fmap(xor_out[288*24*24*bW:289*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[304*5*5:305*5*5-1]), .o_out_fmap(xor_out[304*24*24*bW:305*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[320*5*5:321*5*5-1]), .o_out_fmap(xor_out[320*24*24*bW:321*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[336*5*5:337*5*5-1]), .o_out_fmap(xor_out[336*24*24*bW:337*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[352*5*5:353*5*5-1]), .o_out_fmap(xor_out[352*24*24*bW:353*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[368*5*5:369*5*5-1]), .o_out_fmap(xor_out[368*24*24*bW:369*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[384*5*5:385*5*5-1]), .o_out_fmap(xor_out[384*24*24*bW:385*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[400*5*5:401*5*5-1]), .o_out_fmap(xor_out[400*24*24*bW:401*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[416*5*5:417*5*5-1]), .o_out_fmap(xor_out[416*24*24*bW:417*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[432*5*5:433*5*5-1]), .o_out_fmap(xor_out[432*24*24*bW:433*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[448*5*5:449*5*5-1]), .o_out_fmap(xor_out[448*24*24*bW:449*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[464*5*5:465*5*5-1]), .o_out_fmap(xor_out[464*24*24*bW:465*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[480*5*5:481*5*5-1]), .o_out_fmap(xor_out[480*24*24*bW:481*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[496*5*5:497*5*5-1]), .o_out_fmap(xor_out[496*24*24*bW:497*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[512*5*5:513*5*5-1]), .o_out_fmap(xor_out[512*24*24*bW:513*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[528*5*5:529*5*5-1]), .o_out_fmap(xor_out[528*24*24*bW:529*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[544*5*5:545*5*5-1]), .o_out_fmap(xor_out[544*24*24*bW:545*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[560*5*5:561*5*5-1]), .o_out_fmap(xor_out[560*24*24*bW:561*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[576*5*5:577*5*5-1]), .o_out_fmap(xor_out[576*24*24*bW:577*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[592*5*5:593*5*5-1]), .o_out_fmap(xor_out[592*24*24*bW:593*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[608*5*5:609*5*5-1]), .o_out_fmap(xor_out[608*24*24*bW:609*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[624*5*5:625*5*5-1]), .o_out_fmap(xor_out[624*24*24*bW:625*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[640*5*5:641*5*5-1]), .o_out_fmap(xor_out[640*24*24*bW:641*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[656*5*5:657*5*5-1]), .o_out_fmap(xor_out[656*24*24*bW:657*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[672*5*5:673*5*5-1]), .o_out_fmap(xor_out[672*24*24*bW:673*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[688*5*5:689*5*5-1]), .o_out_fmap(xor_out[688*24*24*bW:689*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[704*5*5:705*5*5-1]), .o_out_fmap(xor_out[704*24*24*bW:705*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[720*5*5:721*5*5-1]), .o_out_fmap(xor_out[720*24*24*bW:721*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[736*5*5:737*5*5-1]), .o_out_fmap(xor_out[736*24*24*bW:737*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[752*5*5:753*5*5-1]), .o_out_fmap(xor_out[752*24*24*bW:753*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[768*5*5:769*5*5-1]), .o_out_fmap(xor_out[768*24*24*bW:769*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[784*5*5:785*5*5-1]), .o_out_fmap(xor_out[784*24*24*bW:785*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[800*5*5:801*5*5-1]), .o_out_fmap(xor_out[800*24*24*bW:801*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[816*5*5:817*5*5-1]), .o_out_fmap(xor_out[816*24*24*bW:817*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[832*5*5:833*5*5-1]), .o_out_fmap(xor_out[832*24*24*bW:833*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[848*5*5:849*5*5-1]), .o_out_fmap(xor_out[848*24*24*bW:849*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[864*5*5:865*5*5-1]), .o_out_fmap(xor_out[864*24*24*bW:865*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[880*5*5:881*5*5-1]), .o_out_fmap(xor_out[880*24*24*bW:881*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[896*5*5:897*5*5-1]), .o_out_fmap(xor_out[896*24*24*bW:897*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[912*5*5:913*5*5-1]), .o_out_fmap(xor_out[912*24*24*bW:913*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[928*5*5:929*5*5-1]), .o_out_fmap(xor_out[928*24*24*bW:929*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[16*12*12:17*12*12-1]), .i_kernel(kernels[944*5*5:945*5*5-1]), .o_out_fmap(xor_out[944*24*24*bW:945*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[17*5*5:18*5*5-1]), .o_out_fmap(xor_out[17*24*24*bW:18*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[34*5*5:35*5*5-1]), .o_out_fmap(xor_out[34*24*24*bW:35*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[51*5*5:52*5*5-1]), .o_out_fmap(xor_out[51*24*24*bW:52*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[68*5*5:69*5*5-1]), .o_out_fmap(xor_out[68*24*24*bW:69*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[85*5*5:86*5*5-1]), .o_out_fmap(xor_out[85*24*24*bW:86*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[102*5*5:103*5*5-1]), .o_out_fmap(xor_out[102*24*24*bW:103*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[119*5*5:120*5*5-1]), .o_out_fmap(xor_out[119*24*24*bW:120*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[136*5*5:137*5*5-1]), .o_out_fmap(xor_out[136*24*24*bW:137*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[153*5*5:154*5*5-1]), .o_out_fmap(xor_out[153*24*24*bW:154*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[170*5*5:171*5*5-1]), .o_out_fmap(xor_out[170*24*24*bW:171*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[187*5*5:188*5*5-1]), .o_out_fmap(xor_out[187*24*24*bW:188*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[204*5*5:205*5*5-1]), .o_out_fmap(xor_out[204*24*24*bW:205*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[221*5*5:222*5*5-1]), .o_out_fmap(xor_out[221*24*24*bW:222*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[238*5*5:239*5*5-1]), .o_out_fmap(xor_out[238*24*24*bW:239*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[255*5*5:256*5*5-1]), .o_out_fmap(xor_out[255*24*24*bW:256*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[272*5*5:273*5*5-1]), .o_out_fmap(xor_out[272*24*24*bW:273*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[289*5*5:290*5*5-1]), .o_out_fmap(xor_out[289*24*24*bW:290*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[306*5*5:307*5*5-1]), .o_out_fmap(xor_out[306*24*24*bW:307*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[323*5*5:324*5*5-1]), .o_out_fmap(xor_out[323*24*24*bW:324*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[340*5*5:341*5*5-1]), .o_out_fmap(xor_out[340*24*24*bW:341*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[357*5*5:358*5*5-1]), .o_out_fmap(xor_out[357*24*24*bW:358*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[374*5*5:375*5*5-1]), .o_out_fmap(xor_out[374*24*24*bW:375*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[391*5*5:392*5*5-1]), .o_out_fmap(xor_out[391*24*24*bW:392*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[408*5*5:409*5*5-1]), .o_out_fmap(xor_out[408*24*24*bW:409*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[425*5*5:426*5*5-1]), .o_out_fmap(xor_out[425*24*24*bW:426*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[442*5*5:443*5*5-1]), .o_out_fmap(xor_out[442*24*24*bW:443*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[459*5*5:460*5*5-1]), .o_out_fmap(xor_out[459*24*24*bW:460*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[476*5*5:477*5*5-1]), .o_out_fmap(xor_out[476*24*24*bW:477*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[493*5*5:494*5*5-1]), .o_out_fmap(xor_out[493*24*24*bW:494*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[510*5*5:511*5*5-1]), .o_out_fmap(xor_out[510*24*24*bW:511*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[527*5*5:528*5*5-1]), .o_out_fmap(xor_out[527*24*24*bW:528*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[544*5*5:545*5*5-1]), .o_out_fmap(xor_out[544*24*24*bW:545*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[561*5*5:562*5*5-1]), .o_out_fmap(xor_out[561*24*24*bW:562*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[578*5*5:579*5*5-1]), .o_out_fmap(xor_out[578*24*24*bW:579*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[595*5*5:596*5*5-1]), .o_out_fmap(xor_out[595*24*24*bW:596*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[612*5*5:613*5*5-1]), .o_out_fmap(xor_out[612*24*24*bW:613*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[629*5*5:630*5*5-1]), .o_out_fmap(xor_out[629*24*24*bW:630*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[646*5*5:647*5*5-1]), .o_out_fmap(xor_out[646*24*24*bW:647*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[663*5*5:664*5*5-1]), .o_out_fmap(xor_out[663*24*24*bW:664*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[680*5*5:681*5*5-1]), .o_out_fmap(xor_out[680*24*24*bW:681*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[697*5*5:698*5*5-1]), .o_out_fmap(xor_out[697*24*24*bW:698*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[714*5*5:715*5*5-1]), .o_out_fmap(xor_out[714*24*24*bW:715*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[731*5*5:732*5*5-1]), .o_out_fmap(xor_out[731*24*24*bW:732*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[748*5*5:749*5*5-1]), .o_out_fmap(xor_out[748*24*24*bW:749*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[765*5*5:766*5*5-1]), .o_out_fmap(xor_out[765*24*24*bW:766*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[782*5*5:783*5*5-1]), .o_out_fmap(xor_out[782*24*24*bW:783*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[799*5*5:800*5*5-1]), .o_out_fmap(xor_out[799*24*24*bW:800*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[816*5*5:817*5*5-1]), .o_out_fmap(xor_out[816*24*24*bW:817*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[833*5*5:834*5*5-1]), .o_out_fmap(xor_out[833*24*24*bW:834*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[850*5*5:851*5*5-1]), .o_out_fmap(xor_out[850*24*24*bW:851*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[867*5*5:868*5*5-1]), .o_out_fmap(xor_out[867*24*24*bW:868*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[884*5*5:885*5*5-1]), .o_out_fmap(xor_out[884*24*24*bW:885*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[901*5*5:902*5*5-1]), .o_out_fmap(xor_out[901*24*24*bW:902*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[918*5*5:919*5*5-1]), .o_out_fmap(xor_out[918*24*24*bW:919*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[935*5*5:936*5*5-1]), .o_out_fmap(xor_out[935*24*24*bW:936*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[952*5*5:953*5*5-1]), .o_out_fmap(xor_out[952*24*24*bW:953*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[969*5*5:970*5*5-1]), .o_out_fmap(xor_out[969*24*24*bW:970*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[986*5*5:987*5*5-1]), .o_out_fmap(xor_out[986*24*24*bW:987*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[17*12*12:18*12*12-1]), .i_kernel(kernels[1003*5*5:1004*5*5-1]), .o_out_fmap(xor_out[1003*24*24*bW:1004*24*24*bW-1]));

endmodule