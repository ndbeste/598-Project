module conv2
    #( parameter bW = 8 )
    (
    input  logic [0:18*12*12 -1] image         ,
    input  logic [0:18*60*5*5-1] kernels       ,
    input  logic [0:60*bW    -1] kernel_offset ,
    output logic [0:60*8*8   -1] conv_one_out 
    );

logic [0:18*60*24*24*bW-1] xor_out;

convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*24*24*bW:1*24*24*bW-1]));
convchan2 c_2_1 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[1*5*5:2*5*5-1]), .o_out_fmap(xor_out[1*24*24*bW:2*24*24*bW-1]));
convchan2 c_2_2 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[2*5*5:3*5*5-1]), .o_out_fmap(xor_out[2*24*24*bW:3*24*24*bW-1]));
convchan2 c_2_3 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[3*5*5:4*5*5-1]), .o_out_fmap(xor_out[3*24*24*bW:4*24*24*bW-1]));
convchan2 c_2_4 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[4*5*5:5*5*5-1]), .o_out_fmap(xor_out[4*24*24*bW:5*24*24*bW-1]));
convchan2 c_2_5 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[5*5*5:6*5*5-1]), .o_out_fmap(xor_out[5*24*24*bW:6*24*24*bW-1]));
convchan2 c_2_6 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[6*5*5:7*5*5-1]), .o_out_fmap(xor_out[6*24*24*bW:7*24*24*bW-1]));
convchan2 c_2_7 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[7*5*5:8*5*5-1]), .o_out_fmap(xor_out[7*24*24*bW:8*24*24*bW-1]));
convchan2 c_2_8 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[8*5*5:9*5*5-1]), .o_out_fmap(xor_out[8*24*24*bW:9*24*24*bW-1]));
convchan2 c_2_9 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[9*5*5:10*5*5-1]), .o_out_fmap(xor_out[9*24*24*bW:10*24*24*bW-1]));
convchan2 c_2_10 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[10*5*5:11*5*5-1]), .o_out_fmap(xor_out[10*24*24*bW:11*24*24*bW-1]));
convchan2 c_2_11 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[11*5*5:12*5*5-1]), .o_out_fmap(xor_out[11*24*24*bW:12*24*24*bW-1]));
convchan2 c_2_12 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[12*5*5:13*5*5-1]), .o_out_fmap(xor_out[12*24*24*bW:13*24*24*bW-1]));
convchan2 c_2_13 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[13*5*5:14*5*5-1]), .o_out_fmap(xor_out[13*24*24*bW:14*24*24*bW-1]));
convchan2 c_2_14 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[14*5*5:15*5*5-1]), .o_out_fmap(xor_out[14*24*24*bW:15*24*24*bW-1]));
convchan2 c_2_15 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[15*5*5:16*5*5-1]), .o_out_fmap(xor_out[15*24*24*bW:16*24*24*bW-1]));
convchan2 c_2_16 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[16*5*5:17*5*5-1]), .o_out_fmap(xor_out[16*24*24*bW:17*24*24*bW-1]));
convchan2 c_2_17 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[17*5*5:18*5*5-1]), .o_out_fmap(xor_out[17*24*24*bW:18*24*24*bW-1]));
convchan2 c_2_18 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[18*5*5:19*5*5-1]), .o_out_fmap(xor_out[18*24*24*bW:19*24*24*bW-1]));
convchan2 c_2_19 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[19*5*5:20*5*5-1]), .o_out_fmap(xor_out[19*24*24*bW:20*24*24*bW-1]));
convchan2 c_2_20 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[20*5*5:21*5*5-1]), .o_out_fmap(xor_out[20*24*24*bW:21*24*24*bW-1]));
convchan2 c_2_21 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[21*5*5:22*5*5-1]), .o_out_fmap(xor_out[21*24*24*bW:22*24*24*bW-1]));
convchan2 c_2_22 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[22*5*5:23*5*5-1]), .o_out_fmap(xor_out[22*24*24*bW:23*24*24*bW-1]));
convchan2 c_2_23 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[23*5*5:24*5*5-1]), .o_out_fmap(xor_out[23*24*24*bW:24*24*24*bW-1]));
convchan2 c_2_24 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[24*5*5:25*5*5-1]), .o_out_fmap(xor_out[24*24*24*bW:25*24*24*bW-1]));
convchan2 c_2_25 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[25*5*5:26*5*5-1]), .o_out_fmap(xor_out[25*24*24*bW:26*24*24*bW-1]));
convchan2 c_2_26 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[26*5*5:27*5*5-1]), .o_out_fmap(xor_out[26*24*24*bW:27*24*24*bW-1]));
convchan2 c_2_27 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[27*5*5:28*5*5-1]), .o_out_fmap(xor_out[27*24*24*bW:28*24*24*bW-1]));
convchan2 c_2_28 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[28*5*5:29*5*5-1]), .o_out_fmap(xor_out[28*24*24*bW:29*24*24*bW-1]));
convchan2 c_2_29 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[29*5*5:30*5*5-1]), .o_out_fmap(xor_out[29*24*24*bW:30*24*24*bW-1]));
convchan2 c_2_30 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[30*5*5:31*5*5-1]), .o_out_fmap(xor_out[30*24*24*bW:31*24*24*bW-1]));
convchan2 c_2_31 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[31*5*5:32*5*5-1]), .o_out_fmap(xor_out[31*24*24*bW:32*24*24*bW-1]));
convchan2 c_2_32 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[32*5*5:33*5*5-1]), .o_out_fmap(xor_out[32*24*24*bW:33*24*24*bW-1]));
convchan2 c_2_33 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[33*5*5:34*5*5-1]), .o_out_fmap(xor_out[33*24*24*bW:34*24*24*bW-1]));
convchan2 c_2_34 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[34*5*5:35*5*5-1]), .o_out_fmap(xor_out[34*24*24*bW:35*24*24*bW-1]));
convchan2 c_2_35 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[35*5*5:36*5*5-1]), .o_out_fmap(xor_out[35*24*24*bW:36*24*24*bW-1]));
convchan2 c_2_36 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[36*5*5:37*5*5-1]), .o_out_fmap(xor_out[36*24*24*bW:37*24*24*bW-1]));
convchan2 c_2_37 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[37*5*5:38*5*5-1]), .o_out_fmap(xor_out[37*24*24*bW:38*24*24*bW-1]));
convchan2 c_2_38 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[38*5*5:39*5*5-1]), .o_out_fmap(xor_out[38*24*24*bW:39*24*24*bW-1]));
convchan2 c_2_39 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[39*5*5:40*5*5-1]), .o_out_fmap(xor_out[39*24*24*bW:40*24*24*bW-1]));
convchan2 c_2_40 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[40*5*5:41*5*5-1]), .o_out_fmap(xor_out[40*24*24*bW:41*24*24*bW-1]));
convchan2 c_2_41 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[41*5*5:42*5*5-1]), .o_out_fmap(xor_out[41*24*24*bW:42*24*24*bW-1]));
convchan2 c_2_42 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[42*5*5:43*5*5-1]), .o_out_fmap(xor_out[42*24*24*bW:43*24*24*bW-1]));
convchan2 c_2_43 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[43*5*5:44*5*5-1]), .o_out_fmap(xor_out[43*24*24*bW:44*24*24*bW-1]));
convchan2 c_2_44 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[44*5*5:45*5*5-1]), .o_out_fmap(xor_out[44*24*24*bW:45*24*24*bW-1]));
convchan2 c_2_45 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[45*5*5:46*5*5-1]), .o_out_fmap(xor_out[45*24*24*bW:46*24*24*bW-1]));
convchan2 c_2_46 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[46*5*5:47*5*5-1]), .o_out_fmap(xor_out[46*24*24*bW:47*24*24*bW-1]));
convchan2 c_2_47 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[47*5*5:48*5*5-1]), .o_out_fmap(xor_out[47*24*24*bW:48*24*24*bW-1]));
convchan2 c_2_48 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[48*5*5:49*5*5-1]), .o_out_fmap(xor_out[48*24*24*bW:49*24*24*bW-1]));
convchan2 c_2_49 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[49*5*5:50*5*5-1]), .o_out_fmap(xor_out[49*24*24*bW:50*24*24*bW-1]));
convchan2 c_2_50 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[50*5*5:51*5*5-1]), .o_out_fmap(xor_out[50*24*24*bW:51*24*24*bW-1]));
convchan2 c_2_51 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[51*5*5:52*5*5-1]), .o_out_fmap(xor_out[51*24*24*bW:52*24*24*bW-1]));
convchan2 c_2_52 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[52*5*5:53*5*5-1]), .o_out_fmap(xor_out[52*24*24*bW:53*24*24*bW-1]));
convchan2 c_2_53 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[53*5*5:54*5*5-1]), .o_out_fmap(xor_out[53*24*24*bW:54*24*24*bW-1]));
convchan2 c_2_54 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[54*5*5:55*5*5-1]), .o_out_fmap(xor_out[54*24*24*bW:55*24*24*bW-1]));
convchan2 c_2_55 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[55*5*5:56*5*5-1]), .o_out_fmap(xor_out[55*24*24*bW:56*24*24*bW-1]));
convchan2 c_2_56 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[56*5*5:57*5*5-1]), .o_out_fmap(xor_out[56*24*24*bW:57*24*24*bW-1]));
convchan2 c_2_57 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[57*5*5:58*5*5-1]), .o_out_fmap(xor_out[57*24*24*bW:58*24*24*bW-1]));
convchan2 c_2_58 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[58*5*5:59*5*5-1]), .o_out_fmap(xor_out[58*24*24*bW:59*24*24*bW-1]));
convchan2 c_2_59 (.i_image(image[0*12*12:1*12*12*+1]), .i_kernel(kernels[59*5*5:60*5*5-1]), .o_out_fmap(xor_out[59*24*24*bW:60*24*24*bW-1]));
convchan2 c_2_60 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[60*5*5:61*5*5-1]), .o_out_fmap(xor_out[60*24*24*bW:61*24*24*bW-1]));
convchan2 c_2_61 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[61*5*5:62*5*5-1]), .o_out_fmap(xor_out[61*24*24*bW:62*24*24*bW-1]));
convchan2 c_2_62 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[62*5*5:63*5*5-1]), .o_out_fmap(xor_out[62*24*24*bW:63*24*24*bW-1]));
convchan2 c_2_63 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[63*5*5:64*5*5-1]), .o_out_fmap(xor_out[63*24*24*bW:64*24*24*bW-1]));
convchan2 c_2_64 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[64*5*5:65*5*5-1]), .o_out_fmap(xor_out[64*24*24*bW:65*24*24*bW-1]));
convchan2 c_2_65 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[65*5*5:66*5*5-1]), .o_out_fmap(xor_out[65*24*24*bW:66*24*24*bW-1]));
convchan2 c_2_66 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[66*5*5:67*5*5-1]), .o_out_fmap(xor_out[66*24*24*bW:67*24*24*bW-1]));
convchan2 c_2_67 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[67*5*5:68*5*5-1]), .o_out_fmap(xor_out[67*24*24*bW:68*24*24*bW-1]));
convchan2 c_2_68 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[68*5*5:69*5*5-1]), .o_out_fmap(xor_out[68*24*24*bW:69*24*24*bW-1]));
convchan2 c_2_69 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[69*5*5:70*5*5-1]), .o_out_fmap(xor_out[69*24*24*bW:70*24*24*bW-1]));
convchan2 c_2_70 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[70*5*5:71*5*5-1]), .o_out_fmap(xor_out[70*24*24*bW:71*24*24*bW-1]));
convchan2 c_2_71 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[71*5*5:72*5*5-1]), .o_out_fmap(xor_out[71*24*24*bW:72*24*24*bW-1]));
convchan2 c_2_72 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[72*5*5:73*5*5-1]), .o_out_fmap(xor_out[72*24*24*bW:73*24*24*bW-1]));
convchan2 c_2_73 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[73*5*5:74*5*5-1]), .o_out_fmap(xor_out[73*24*24*bW:74*24*24*bW-1]));
convchan2 c_2_74 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[74*5*5:75*5*5-1]), .o_out_fmap(xor_out[74*24*24*bW:75*24*24*bW-1]));
convchan2 c_2_75 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[75*5*5:76*5*5-1]), .o_out_fmap(xor_out[75*24*24*bW:76*24*24*bW-1]));
convchan2 c_2_76 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[76*5*5:77*5*5-1]), .o_out_fmap(xor_out[76*24*24*bW:77*24*24*bW-1]));
convchan2 c_2_77 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[77*5*5:78*5*5-1]), .o_out_fmap(xor_out[77*24*24*bW:78*24*24*bW-1]));
convchan2 c_2_78 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[78*5*5:79*5*5-1]), .o_out_fmap(xor_out[78*24*24*bW:79*24*24*bW-1]));
convchan2 c_2_79 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[79*5*5:80*5*5-1]), .o_out_fmap(xor_out[79*24*24*bW:80*24*24*bW-1]));
convchan2 c_2_80 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[80*5*5:81*5*5-1]), .o_out_fmap(xor_out[80*24*24*bW:81*24*24*bW-1]));
convchan2 c_2_81 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[81*5*5:82*5*5-1]), .o_out_fmap(xor_out[81*24*24*bW:82*24*24*bW-1]));
convchan2 c_2_82 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[82*5*5:83*5*5-1]), .o_out_fmap(xor_out[82*24*24*bW:83*24*24*bW-1]));
convchan2 c_2_83 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[83*5*5:84*5*5-1]), .o_out_fmap(xor_out[83*24*24*bW:84*24*24*bW-1]));
convchan2 c_2_84 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[84*5*5:85*5*5-1]), .o_out_fmap(xor_out[84*24*24*bW:85*24*24*bW-1]));
convchan2 c_2_85 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[85*5*5:86*5*5-1]), .o_out_fmap(xor_out[85*24*24*bW:86*24*24*bW-1]));
convchan2 c_2_86 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[86*5*5:87*5*5-1]), .o_out_fmap(xor_out[86*24*24*bW:87*24*24*bW-1]));
convchan2 c_2_87 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[87*5*5:88*5*5-1]), .o_out_fmap(xor_out[87*24*24*bW:88*24*24*bW-1]));
convchan2 c_2_88 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[88*5*5:89*5*5-1]), .o_out_fmap(xor_out[88*24*24*bW:89*24*24*bW-1]));
convchan2 c_2_89 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[89*5*5:90*5*5-1]), .o_out_fmap(xor_out[89*24*24*bW:90*24*24*bW-1]));
convchan2 c_2_90 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[90*5*5:91*5*5-1]), .o_out_fmap(xor_out[90*24*24*bW:91*24*24*bW-1]));
convchan2 c_2_91 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[91*5*5:92*5*5-1]), .o_out_fmap(xor_out[91*24*24*bW:92*24*24*bW-1]));
convchan2 c_2_92 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[92*5*5:93*5*5-1]), .o_out_fmap(xor_out[92*24*24*bW:93*24*24*bW-1]));
convchan2 c_2_93 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[93*5*5:94*5*5-1]), .o_out_fmap(xor_out[93*24*24*bW:94*24*24*bW-1]));
convchan2 c_2_94 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[94*5*5:95*5*5-1]), .o_out_fmap(xor_out[94*24*24*bW:95*24*24*bW-1]));
convchan2 c_2_95 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[95*5*5:96*5*5-1]), .o_out_fmap(xor_out[95*24*24*bW:96*24*24*bW-1]));
convchan2 c_2_96 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[96*5*5:97*5*5-1]), .o_out_fmap(xor_out[96*24*24*bW:97*24*24*bW-1]));
convchan2 c_2_97 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[97*5*5:98*5*5-1]), .o_out_fmap(xor_out[97*24*24*bW:98*24*24*bW-1]));
convchan2 c_2_98 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[98*5*5:99*5*5-1]), .o_out_fmap(xor_out[98*24*24*bW:99*24*24*bW-1]));
convchan2 c_2_99 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[99*5*5:100*5*5-1]), .o_out_fmap(xor_out[99*24*24*bW:100*24*24*bW-1]));
convchan2 c_2_100 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[100*5*5:101*5*5-1]), .o_out_fmap(xor_out[100*24*24*bW:101*24*24*bW-1]));
convchan2 c_2_101 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[101*5*5:102*5*5-1]), .o_out_fmap(xor_out[101*24*24*bW:102*24*24*bW-1]));
convchan2 c_2_102 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[102*5*5:103*5*5-1]), .o_out_fmap(xor_out[102*24*24*bW:103*24*24*bW-1]));
convchan2 c_2_103 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[103*5*5:104*5*5-1]), .o_out_fmap(xor_out[103*24*24*bW:104*24*24*bW-1]));
convchan2 c_2_104 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[104*5*5:105*5*5-1]), .o_out_fmap(xor_out[104*24*24*bW:105*24*24*bW-1]));
convchan2 c_2_105 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[105*5*5:106*5*5-1]), .o_out_fmap(xor_out[105*24*24*bW:106*24*24*bW-1]));
convchan2 c_2_106 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[106*5*5:107*5*5-1]), .o_out_fmap(xor_out[106*24*24*bW:107*24*24*bW-1]));
convchan2 c_2_107 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[107*5*5:108*5*5-1]), .o_out_fmap(xor_out[107*24*24*bW:108*24*24*bW-1]));
convchan2 c_2_108 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[108*5*5:109*5*5-1]), .o_out_fmap(xor_out[108*24*24*bW:109*24*24*bW-1]));
convchan2 c_2_109 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[109*5*5:110*5*5-1]), .o_out_fmap(xor_out[109*24*24*bW:110*24*24*bW-1]));
convchan2 c_2_110 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[110*5*5:111*5*5-1]), .o_out_fmap(xor_out[110*24*24*bW:111*24*24*bW-1]));
convchan2 c_2_111 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[111*5*5:112*5*5-1]), .o_out_fmap(xor_out[111*24*24*bW:112*24*24*bW-1]));
convchan2 c_2_112 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[112*5*5:113*5*5-1]), .o_out_fmap(xor_out[112*24*24*bW:113*24*24*bW-1]));
convchan2 c_2_113 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[113*5*5:114*5*5-1]), .o_out_fmap(xor_out[113*24*24*bW:114*24*24*bW-1]));
convchan2 c_2_114 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[114*5*5:115*5*5-1]), .o_out_fmap(xor_out[114*24*24*bW:115*24*24*bW-1]));
convchan2 c_2_115 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[115*5*5:116*5*5-1]), .o_out_fmap(xor_out[115*24*24*bW:116*24*24*bW-1]));
convchan2 c_2_116 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[116*5*5:117*5*5-1]), .o_out_fmap(xor_out[116*24*24*bW:117*24*24*bW-1]));
convchan2 c_2_117 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[117*5*5:118*5*5-1]), .o_out_fmap(xor_out[117*24*24*bW:118*24*24*bW-1]));
convchan2 c_2_118 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[118*5*5:119*5*5-1]), .o_out_fmap(xor_out[118*24*24*bW:119*24*24*bW-1]));
convchan2 c_2_119 (.i_image(image[1*12*12:2*12*12*+1]), .i_kernel(kernels[119*5*5:120*5*5-1]), .o_out_fmap(xor_out[119*24*24*bW:120*24*24*bW-1]));
convchan2 c_2_120 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[120*5*5:121*5*5-1]), .o_out_fmap(xor_out[120*24*24*bW:121*24*24*bW-1]));
convchan2 c_2_121 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[121*5*5:122*5*5-1]), .o_out_fmap(xor_out[121*24*24*bW:122*24*24*bW-1]));
convchan2 c_2_122 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[122*5*5:123*5*5-1]), .o_out_fmap(xor_out[122*24*24*bW:123*24*24*bW-1]));
convchan2 c_2_123 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[123*5*5:124*5*5-1]), .o_out_fmap(xor_out[123*24*24*bW:124*24*24*bW-1]));
convchan2 c_2_124 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[124*5*5:125*5*5-1]), .o_out_fmap(xor_out[124*24*24*bW:125*24*24*bW-1]));
convchan2 c_2_125 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[125*5*5:126*5*5-1]), .o_out_fmap(xor_out[125*24*24*bW:126*24*24*bW-1]));
convchan2 c_2_126 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[126*5*5:127*5*5-1]), .o_out_fmap(xor_out[126*24*24*bW:127*24*24*bW-1]));
convchan2 c_2_127 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[127*5*5:128*5*5-1]), .o_out_fmap(xor_out[127*24*24*bW:128*24*24*bW-1]));
convchan2 c_2_128 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[128*5*5:129*5*5-1]), .o_out_fmap(xor_out[128*24*24*bW:129*24*24*bW-1]));
convchan2 c_2_129 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[129*5*5:130*5*5-1]), .o_out_fmap(xor_out[129*24*24*bW:130*24*24*bW-1]));
convchan2 c_2_130 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[130*5*5:131*5*5-1]), .o_out_fmap(xor_out[130*24*24*bW:131*24*24*bW-1]));
convchan2 c_2_131 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[131*5*5:132*5*5-1]), .o_out_fmap(xor_out[131*24*24*bW:132*24*24*bW-1]));
convchan2 c_2_132 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[132*5*5:133*5*5-1]), .o_out_fmap(xor_out[132*24*24*bW:133*24*24*bW-1]));
convchan2 c_2_133 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[133*5*5:134*5*5-1]), .o_out_fmap(xor_out[133*24*24*bW:134*24*24*bW-1]));
convchan2 c_2_134 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[134*5*5:135*5*5-1]), .o_out_fmap(xor_out[134*24*24*bW:135*24*24*bW-1]));
convchan2 c_2_135 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[135*5*5:136*5*5-1]), .o_out_fmap(xor_out[135*24*24*bW:136*24*24*bW-1]));
convchan2 c_2_136 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[136*5*5:137*5*5-1]), .o_out_fmap(xor_out[136*24*24*bW:137*24*24*bW-1]));
convchan2 c_2_137 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[137*5*5:138*5*5-1]), .o_out_fmap(xor_out[137*24*24*bW:138*24*24*bW-1]));
convchan2 c_2_138 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[138*5*5:139*5*5-1]), .o_out_fmap(xor_out[138*24*24*bW:139*24*24*bW-1]));
convchan2 c_2_139 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[139*5*5:140*5*5-1]), .o_out_fmap(xor_out[139*24*24*bW:140*24*24*bW-1]));
convchan2 c_2_140 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[140*5*5:141*5*5-1]), .o_out_fmap(xor_out[140*24*24*bW:141*24*24*bW-1]));
convchan2 c_2_141 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[141*5*5:142*5*5-1]), .o_out_fmap(xor_out[141*24*24*bW:142*24*24*bW-1]));
convchan2 c_2_142 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[142*5*5:143*5*5-1]), .o_out_fmap(xor_out[142*24*24*bW:143*24*24*bW-1]));
convchan2 c_2_143 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[143*5*5:144*5*5-1]), .o_out_fmap(xor_out[143*24*24*bW:144*24*24*bW-1]));
convchan2 c_2_144 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[144*5*5:145*5*5-1]), .o_out_fmap(xor_out[144*24*24*bW:145*24*24*bW-1]));
convchan2 c_2_145 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[145*5*5:146*5*5-1]), .o_out_fmap(xor_out[145*24*24*bW:146*24*24*bW-1]));
convchan2 c_2_146 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[146*5*5:147*5*5-1]), .o_out_fmap(xor_out[146*24*24*bW:147*24*24*bW-1]));
convchan2 c_2_147 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[147*5*5:148*5*5-1]), .o_out_fmap(xor_out[147*24*24*bW:148*24*24*bW-1]));
convchan2 c_2_148 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[148*5*5:149*5*5-1]), .o_out_fmap(xor_out[148*24*24*bW:149*24*24*bW-1]));
convchan2 c_2_149 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[149*5*5:150*5*5-1]), .o_out_fmap(xor_out[149*24*24*bW:150*24*24*bW-1]));
convchan2 c_2_150 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[150*5*5:151*5*5-1]), .o_out_fmap(xor_out[150*24*24*bW:151*24*24*bW-1]));
convchan2 c_2_151 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[151*5*5:152*5*5-1]), .o_out_fmap(xor_out[151*24*24*bW:152*24*24*bW-1]));
convchan2 c_2_152 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[152*5*5:153*5*5-1]), .o_out_fmap(xor_out[152*24*24*bW:153*24*24*bW-1]));
convchan2 c_2_153 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[153*5*5:154*5*5-1]), .o_out_fmap(xor_out[153*24*24*bW:154*24*24*bW-1]));
convchan2 c_2_154 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[154*5*5:155*5*5-1]), .o_out_fmap(xor_out[154*24*24*bW:155*24*24*bW-1]));
convchan2 c_2_155 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[155*5*5:156*5*5-1]), .o_out_fmap(xor_out[155*24*24*bW:156*24*24*bW-1]));
convchan2 c_2_156 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[156*5*5:157*5*5-1]), .o_out_fmap(xor_out[156*24*24*bW:157*24*24*bW-1]));
convchan2 c_2_157 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[157*5*5:158*5*5-1]), .o_out_fmap(xor_out[157*24*24*bW:158*24*24*bW-1]));
convchan2 c_2_158 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[158*5*5:159*5*5-1]), .o_out_fmap(xor_out[158*24*24*bW:159*24*24*bW-1]));
convchan2 c_2_159 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[159*5*5:160*5*5-1]), .o_out_fmap(xor_out[159*24*24*bW:160*24*24*bW-1]));
convchan2 c_2_160 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[160*5*5:161*5*5-1]), .o_out_fmap(xor_out[160*24*24*bW:161*24*24*bW-1]));
convchan2 c_2_161 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[161*5*5:162*5*5-1]), .o_out_fmap(xor_out[161*24*24*bW:162*24*24*bW-1]));
convchan2 c_2_162 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[162*5*5:163*5*5-1]), .o_out_fmap(xor_out[162*24*24*bW:163*24*24*bW-1]));
convchan2 c_2_163 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[163*5*5:164*5*5-1]), .o_out_fmap(xor_out[163*24*24*bW:164*24*24*bW-1]));
convchan2 c_2_164 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[164*5*5:165*5*5-1]), .o_out_fmap(xor_out[164*24*24*bW:165*24*24*bW-1]));
convchan2 c_2_165 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[165*5*5:166*5*5-1]), .o_out_fmap(xor_out[165*24*24*bW:166*24*24*bW-1]));
convchan2 c_2_166 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[166*5*5:167*5*5-1]), .o_out_fmap(xor_out[166*24*24*bW:167*24*24*bW-1]));
convchan2 c_2_167 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[167*5*5:168*5*5-1]), .o_out_fmap(xor_out[167*24*24*bW:168*24*24*bW-1]));
convchan2 c_2_168 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[168*5*5:169*5*5-1]), .o_out_fmap(xor_out[168*24*24*bW:169*24*24*bW-1]));
convchan2 c_2_169 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[169*5*5:170*5*5-1]), .o_out_fmap(xor_out[169*24*24*bW:170*24*24*bW-1]));
convchan2 c_2_170 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[170*5*5:171*5*5-1]), .o_out_fmap(xor_out[170*24*24*bW:171*24*24*bW-1]));
convchan2 c_2_171 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[171*5*5:172*5*5-1]), .o_out_fmap(xor_out[171*24*24*bW:172*24*24*bW-1]));
convchan2 c_2_172 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[172*5*5:173*5*5-1]), .o_out_fmap(xor_out[172*24*24*bW:173*24*24*bW-1]));
convchan2 c_2_173 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[173*5*5:174*5*5-1]), .o_out_fmap(xor_out[173*24*24*bW:174*24*24*bW-1]));
convchan2 c_2_174 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[174*5*5:175*5*5-1]), .o_out_fmap(xor_out[174*24*24*bW:175*24*24*bW-1]));
convchan2 c_2_175 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[175*5*5:176*5*5-1]), .o_out_fmap(xor_out[175*24*24*bW:176*24*24*bW-1]));
convchan2 c_2_176 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[176*5*5:177*5*5-1]), .o_out_fmap(xor_out[176*24*24*bW:177*24*24*bW-1]));
convchan2 c_2_177 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[177*5*5:178*5*5-1]), .o_out_fmap(xor_out[177*24*24*bW:178*24*24*bW-1]));
convchan2 c_2_178 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[178*5*5:179*5*5-1]), .o_out_fmap(xor_out[178*24*24*bW:179*24*24*bW-1]));
convchan2 c_2_179 (.i_image(image[2*12*12:3*12*12*+1]), .i_kernel(kernels[179*5*5:180*5*5-1]), .o_out_fmap(xor_out[179*24*24*bW:180*24*24*bW-1]));
convchan2 c_2_180 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[180*5*5:181*5*5-1]), .o_out_fmap(xor_out[180*24*24*bW:181*24*24*bW-1]));
convchan2 c_2_181 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[181*5*5:182*5*5-1]), .o_out_fmap(xor_out[181*24*24*bW:182*24*24*bW-1]));
convchan2 c_2_182 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[182*5*5:183*5*5-1]), .o_out_fmap(xor_out[182*24*24*bW:183*24*24*bW-1]));
convchan2 c_2_183 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[183*5*5:184*5*5-1]), .o_out_fmap(xor_out[183*24*24*bW:184*24*24*bW-1]));
convchan2 c_2_184 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[184*5*5:185*5*5-1]), .o_out_fmap(xor_out[184*24*24*bW:185*24*24*bW-1]));
convchan2 c_2_185 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[185*5*5:186*5*5-1]), .o_out_fmap(xor_out[185*24*24*bW:186*24*24*bW-1]));
convchan2 c_2_186 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[186*5*5:187*5*5-1]), .o_out_fmap(xor_out[186*24*24*bW:187*24*24*bW-1]));
convchan2 c_2_187 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[187*5*5:188*5*5-1]), .o_out_fmap(xor_out[187*24*24*bW:188*24*24*bW-1]));
convchan2 c_2_188 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[188*5*5:189*5*5-1]), .o_out_fmap(xor_out[188*24*24*bW:189*24*24*bW-1]));
convchan2 c_2_189 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[189*5*5:190*5*5-1]), .o_out_fmap(xor_out[189*24*24*bW:190*24*24*bW-1]));
convchan2 c_2_190 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[190*5*5:191*5*5-1]), .o_out_fmap(xor_out[190*24*24*bW:191*24*24*bW-1]));
convchan2 c_2_191 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[191*5*5:192*5*5-1]), .o_out_fmap(xor_out[191*24*24*bW:192*24*24*bW-1]));
convchan2 c_2_192 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[192*5*5:193*5*5-1]), .o_out_fmap(xor_out[192*24*24*bW:193*24*24*bW-1]));
convchan2 c_2_193 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[193*5*5:194*5*5-1]), .o_out_fmap(xor_out[193*24*24*bW:194*24*24*bW-1]));
convchan2 c_2_194 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[194*5*5:195*5*5-1]), .o_out_fmap(xor_out[194*24*24*bW:195*24*24*bW-1]));
convchan2 c_2_195 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[195*5*5:196*5*5-1]), .o_out_fmap(xor_out[195*24*24*bW:196*24*24*bW-1]));
convchan2 c_2_196 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[196*5*5:197*5*5-1]), .o_out_fmap(xor_out[196*24*24*bW:197*24*24*bW-1]));
convchan2 c_2_197 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[197*5*5:198*5*5-1]), .o_out_fmap(xor_out[197*24*24*bW:198*24*24*bW-1]));
convchan2 c_2_198 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[198*5*5:199*5*5-1]), .o_out_fmap(xor_out[198*24*24*bW:199*24*24*bW-1]));
convchan2 c_2_199 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[199*5*5:200*5*5-1]), .o_out_fmap(xor_out[199*24*24*bW:200*24*24*bW-1]));
convchan2 c_2_200 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[200*5*5:201*5*5-1]), .o_out_fmap(xor_out[200*24*24*bW:201*24*24*bW-1]));
convchan2 c_2_201 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[201*5*5:202*5*5-1]), .o_out_fmap(xor_out[201*24*24*bW:202*24*24*bW-1]));
convchan2 c_2_202 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[202*5*5:203*5*5-1]), .o_out_fmap(xor_out[202*24*24*bW:203*24*24*bW-1]));
convchan2 c_2_203 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[203*5*5:204*5*5-1]), .o_out_fmap(xor_out[203*24*24*bW:204*24*24*bW-1]));
convchan2 c_2_204 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[204*5*5:205*5*5-1]), .o_out_fmap(xor_out[204*24*24*bW:205*24*24*bW-1]));
convchan2 c_2_205 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[205*5*5:206*5*5-1]), .o_out_fmap(xor_out[205*24*24*bW:206*24*24*bW-1]));
convchan2 c_2_206 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[206*5*5:207*5*5-1]), .o_out_fmap(xor_out[206*24*24*bW:207*24*24*bW-1]));
convchan2 c_2_207 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[207*5*5:208*5*5-1]), .o_out_fmap(xor_out[207*24*24*bW:208*24*24*bW-1]));
convchan2 c_2_208 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[208*5*5:209*5*5-1]), .o_out_fmap(xor_out[208*24*24*bW:209*24*24*bW-1]));
convchan2 c_2_209 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[209*5*5:210*5*5-1]), .o_out_fmap(xor_out[209*24*24*bW:210*24*24*bW-1]));
convchan2 c_2_210 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[210*5*5:211*5*5-1]), .o_out_fmap(xor_out[210*24*24*bW:211*24*24*bW-1]));
convchan2 c_2_211 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[211*5*5:212*5*5-1]), .o_out_fmap(xor_out[211*24*24*bW:212*24*24*bW-1]));
convchan2 c_2_212 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[212*5*5:213*5*5-1]), .o_out_fmap(xor_out[212*24*24*bW:213*24*24*bW-1]));
convchan2 c_2_213 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[213*5*5:214*5*5-1]), .o_out_fmap(xor_out[213*24*24*bW:214*24*24*bW-1]));
convchan2 c_2_214 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[214*5*5:215*5*5-1]), .o_out_fmap(xor_out[214*24*24*bW:215*24*24*bW-1]));
convchan2 c_2_215 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[215*5*5:216*5*5-1]), .o_out_fmap(xor_out[215*24*24*bW:216*24*24*bW-1]));
convchan2 c_2_216 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[216*5*5:217*5*5-1]), .o_out_fmap(xor_out[216*24*24*bW:217*24*24*bW-1]));
convchan2 c_2_217 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[217*5*5:218*5*5-1]), .o_out_fmap(xor_out[217*24*24*bW:218*24*24*bW-1]));
convchan2 c_2_218 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[218*5*5:219*5*5-1]), .o_out_fmap(xor_out[218*24*24*bW:219*24*24*bW-1]));
convchan2 c_2_219 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[219*5*5:220*5*5-1]), .o_out_fmap(xor_out[219*24*24*bW:220*24*24*bW-1]));
convchan2 c_2_220 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[220*5*5:221*5*5-1]), .o_out_fmap(xor_out[220*24*24*bW:221*24*24*bW-1]));
convchan2 c_2_221 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[221*5*5:222*5*5-1]), .o_out_fmap(xor_out[221*24*24*bW:222*24*24*bW-1]));
convchan2 c_2_222 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[222*5*5:223*5*5-1]), .o_out_fmap(xor_out[222*24*24*bW:223*24*24*bW-1]));
convchan2 c_2_223 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[223*5*5:224*5*5-1]), .o_out_fmap(xor_out[223*24*24*bW:224*24*24*bW-1]));
convchan2 c_2_224 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[224*5*5:225*5*5-1]), .o_out_fmap(xor_out[224*24*24*bW:225*24*24*bW-1]));
convchan2 c_2_225 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[225*5*5:226*5*5-1]), .o_out_fmap(xor_out[225*24*24*bW:226*24*24*bW-1]));
convchan2 c_2_226 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[226*5*5:227*5*5-1]), .o_out_fmap(xor_out[226*24*24*bW:227*24*24*bW-1]));
convchan2 c_2_227 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[227*5*5:228*5*5-1]), .o_out_fmap(xor_out[227*24*24*bW:228*24*24*bW-1]));
convchan2 c_2_228 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[228*5*5:229*5*5-1]), .o_out_fmap(xor_out[228*24*24*bW:229*24*24*bW-1]));
convchan2 c_2_229 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[229*5*5:230*5*5-1]), .o_out_fmap(xor_out[229*24*24*bW:230*24*24*bW-1]));
convchan2 c_2_230 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[230*5*5:231*5*5-1]), .o_out_fmap(xor_out[230*24*24*bW:231*24*24*bW-1]));
convchan2 c_2_231 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[231*5*5:232*5*5-1]), .o_out_fmap(xor_out[231*24*24*bW:232*24*24*bW-1]));
convchan2 c_2_232 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[232*5*5:233*5*5-1]), .o_out_fmap(xor_out[232*24*24*bW:233*24*24*bW-1]));
convchan2 c_2_233 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[233*5*5:234*5*5-1]), .o_out_fmap(xor_out[233*24*24*bW:234*24*24*bW-1]));
convchan2 c_2_234 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[234*5*5:235*5*5-1]), .o_out_fmap(xor_out[234*24*24*bW:235*24*24*bW-1]));
convchan2 c_2_235 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[235*5*5:236*5*5-1]), .o_out_fmap(xor_out[235*24*24*bW:236*24*24*bW-1]));
convchan2 c_2_236 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[236*5*5:237*5*5-1]), .o_out_fmap(xor_out[236*24*24*bW:237*24*24*bW-1]));
convchan2 c_2_237 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[237*5*5:238*5*5-1]), .o_out_fmap(xor_out[237*24*24*bW:238*24*24*bW-1]));
convchan2 c_2_238 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[238*5*5:239*5*5-1]), .o_out_fmap(xor_out[238*24*24*bW:239*24*24*bW-1]));
convchan2 c_2_239 (.i_image(image[3*12*12:4*12*12*+1]), .i_kernel(kernels[239*5*5:240*5*5-1]), .o_out_fmap(xor_out[239*24*24*bW:240*24*24*bW-1]));
convchan2 c_2_240 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[240*5*5:241*5*5-1]), .o_out_fmap(xor_out[240*24*24*bW:241*24*24*bW-1]));
convchan2 c_2_241 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[241*5*5:242*5*5-1]), .o_out_fmap(xor_out[241*24*24*bW:242*24*24*bW-1]));
convchan2 c_2_242 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[242*5*5:243*5*5-1]), .o_out_fmap(xor_out[242*24*24*bW:243*24*24*bW-1]));
convchan2 c_2_243 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[243*5*5:244*5*5-1]), .o_out_fmap(xor_out[243*24*24*bW:244*24*24*bW-1]));
convchan2 c_2_244 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[244*5*5:245*5*5-1]), .o_out_fmap(xor_out[244*24*24*bW:245*24*24*bW-1]));
convchan2 c_2_245 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[245*5*5:246*5*5-1]), .o_out_fmap(xor_out[245*24*24*bW:246*24*24*bW-1]));
convchan2 c_2_246 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[246*5*5:247*5*5-1]), .o_out_fmap(xor_out[246*24*24*bW:247*24*24*bW-1]));
convchan2 c_2_247 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[247*5*5:248*5*5-1]), .o_out_fmap(xor_out[247*24*24*bW:248*24*24*bW-1]));
convchan2 c_2_248 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[248*5*5:249*5*5-1]), .o_out_fmap(xor_out[248*24*24*bW:249*24*24*bW-1]));
convchan2 c_2_249 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[249*5*5:250*5*5-1]), .o_out_fmap(xor_out[249*24*24*bW:250*24*24*bW-1]));
convchan2 c_2_250 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[250*5*5:251*5*5-1]), .o_out_fmap(xor_out[250*24*24*bW:251*24*24*bW-1]));
convchan2 c_2_251 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[251*5*5:252*5*5-1]), .o_out_fmap(xor_out[251*24*24*bW:252*24*24*bW-1]));
convchan2 c_2_252 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[252*5*5:253*5*5-1]), .o_out_fmap(xor_out[252*24*24*bW:253*24*24*bW-1]));
convchan2 c_2_253 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[253*5*5:254*5*5-1]), .o_out_fmap(xor_out[253*24*24*bW:254*24*24*bW-1]));
convchan2 c_2_254 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[254*5*5:255*5*5-1]), .o_out_fmap(xor_out[254*24*24*bW:255*24*24*bW-1]));
convchan2 c_2_255 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[255*5*5:256*5*5-1]), .o_out_fmap(xor_out[255*24*24*bW:256*24*24*bW-1]));
convchan2 c_2_256 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[256*5*5:257*5*5-1]), .o_out_fmap(xor_out[256*24*24*bW:257*24*24*bW-1]));
convchan2 c_2_257 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[257*5*5:258*5*5-1]), .o_out_fmap(xor_out[257*24*24*bW:258*24*24*bW-1]));
convchan2 c_2_258 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[258*5*5:259*5*5-1]), .o_out_fmap(xor_out[258*24*24*bW:259*24*24*bW-1]));
convchan2 c_2_259 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[259*5*5:260*5*5-1]), .o_out_fmap(xor_out[259*24*24*bW:260*24*24*bW-1]));
convchan2 c_2_260 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[260*5*5:261*5*5-1]), .o_out_fmap(xor_out[260*24*24*bW:261*24*24*bW-1]));
convchan2 c_2_261 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[261*5*5:262*5*5-1]), .o_out_fmap(xor_out[261*24*24*bW:262*24*24*bW-1]));
convchan2 c_2_262 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[262*5*5:263*5*5-1]), .o_out_fmap(xor_out[262*24*24*bW:263*24*24*bW-1]));
convchan2 c_2_263 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[263*5*5:264*5*5-1]), .o_out_fmap(xor_out[263*24*24*bW:264*24*24*bW-1]));
convchan2 c_2_264 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[264*5*5:265*5*5-1]), .o_out_fmap(xor_out[264*24*24*bW:265*24*24*bW-1]));
convchan2 c_2_265 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[265*5*5:266*5*5-1]), .o_out_fmap(xor_out[265*24*24*bW:266*24*24*bW-1]));
convchan2 c_2_266 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[266*5*5:267*5*5-1]), .o_out_fmap(xor_out[266*24*24*bW:267*24*24*bW-1]));
convchan2 c_2_267 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[267*5*5:268*5*5-1]), .o_out_fmap(xor_out[267*24*24*bW:268*24*24*bW-1]));
convchan2 c_2_268 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[268*5*5:269*5*5-1]), .o_out_fmap(xor_out[268*24*24*bW:269*24*24*bW-1]));
convchan2 c_2_269 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[269*5*5:270*5*5-1]), .o_out_fmap(xor_out[269*24*24*bW:270*24*24*bW-1]));
convchan2 c_2_270 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[270*5*5:271*5*5-1]), .o_out_fmap(xor_out[270*24*24*bW:271*24*24*bW-1]));
convchan2 c_2_271 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[271*5*5:272*5*5-1]), .o_out_fmap(xor_out[271*24*24*bW:272*24*24*bW-1]));
convchan2 c_2_272 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[272*5*5:273*5*5-1]), .o_out_fmap(xor_out[272*24*24*bW:273*24*24*bW-1]));
convchan2 c_2_273 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[273*5*5:274*5*5-1]), .o_out_fmap(xor_out[273*24*24*bW:274*24*24*bW-1]));
convchan2 c_2_274 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[274*5*5:275*5*5-1]), .o_out_fmap(xor_out[274*24*24*bW:275*24*24*bW-1]));
convchan2 c_2_275 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[275*5*5:276*5*5-1]), .o_out_fmap(xor_out[275*24*24*bW:276*24*24*bW-1]));
convchan2 c_2_276 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[276*5*5:277*5*5-1]), .o_out_fmap(xor_out[276*24*24*bW:277*24*24*bW-1]));
convchan2 c_2_277 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[277*5*5:278*5*5-1]), .o_out_fmap(xor_out[277*24*24*bW:278*24*24*bW-1]));
convchan2 c_2_278 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[278*5*5:279*5*5-1]), .o_out_fmap(xor_out[278*24*24*bW:279*24*24*bW-1]));
convchan2 c_2_279 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[279*5*5:280*5*5-1]), .o_out_fmap(xor_out[279*24*24*bW:280*24*24*bW-1]));
convchan2 c_2_280 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[280*5*5:281*5*5-1]), .o_out_fmap(xor_out[280*24*24*bW:281*24*24*bW-1]));
convchan2 c_2_281 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[281*5*5:282*5*5-1]), .o_out_fmap(xor_out[281*24*24*bW:282*24*24*bW-1]));
convchan2 c_2_282 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[282*5*5:283*5*5-1]), .o_out_fmap(xor_out[282*24*24*bW:283*24*24*bW-1]));
convchan2 c_2_283 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[283*5*5:284*5*5-1]), .o_out_fmap(xor_out[283*24*24*bW:284*24*24*bW-1]));
convchan2 c_2_284 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[284*5*5:285*5*5-1]), .o_out_fmap(xor_out[284*24*24*bW:285*24*24*bW-1]));
convchan2 c_2_285 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[285*5*5:286*5*5-1]), .o_out_fmap(xor_out[285*24*24*bW:286*24*24*bW-1]));
convchan2 c_2_286 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[286*5*5:287*5*5-1]), .o_out_fmap(xor_out[286*24*24*bW:287*24*24*bW-1]));
convchan2 c_2_287 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[287*5*5:288*5*5-1]), .o_out_fmap(xor_out[287*24*24*bW:288*24*24*bW-1]));
convchan2 c_2_288 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[288*5*5:289*5*5-1]), .o_out_fmap(xor_out[288*24*24*bW:289*24*24*bW-1]));
convchan2 c_2_289 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[289*5*5:290*5*5-1]), .o_out_fmap(xor_out[289*24*24*bW:290*24*24*bW-1]));
convchan2 c_2_290 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[290*5*5:291*5*5-1]), .o_out_fmap(xor_out[290*24*24*bW:291*24*24*bW-1]));
convchan2 c_2_291 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[291*5*5:292*5*5-1]), .o_out_fmap(xor_out[291*24*24*bW:292*24*24*bW-1]));
convchan2 c_2_292 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[292*5*5:293*5*5-1]), .o_out_fmap(xor_out[292*24*24*bW:293*24*24*bW-1]));
convchan2 c_2_293 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[293*5*5:294*5*5-1]), .o_out_fmap(xor_out[293*24*24*bW:294*24*24*bW-1]));
convchan2 c_2_294 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[294*5*5:295*5*5-1]), .o_out_fmap(xor_out[294*24*24*bW:295*24*24*bW-1]));
convchan2 c_2_295 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[295*5*5:296*5*5-1]), .o_out_fmap(xor_out[295*24*24*bW:296*24*24*bW-1]));
convchan2 c_2_296 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[296*5*5:297*5*5-1]), .o_out_fmap(xor_out[296*24*24*bW:297*24*24*bW-1]));
convchan2 c_2_297 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[297*5*5:298*5*5-1]), .o_out_fmap(xor_out[297*24*24*bW:298*24*24*bW-1]));
convchan2 c_2_298 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[298*5*5:299*5*5-1]), .o_out_fmap(xor_out[298*24*24*bW:299*24*24*bW-1]));
convchan2 c_2_299 (.i_image(image[4*12*12:5*12*12*+1]), .i_kernel(kernels[299*5*5:300*5*5-1]), .o_out_fmap(xor_out[299*24*24*bW:300*24*24*bW-1]));
convchan2 c_2_300 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[300*5*5:301*5*5-1]), .o_out_fmap(xor_out[300*24*24*bW:301*24*24*bW-1]));
convchan2 c_2_301 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[301*5*5:302*5*5-1]), .o_out_fmap(xor_out[301*24*24*bW:302*24*24*bW-1]));
convchan2 c_2_302 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[302*5*5:303*5*5-1]), .o_out_fmap(xor_out[302*24*24*bW:303*24*24*bW-1]));
convchan2 c_2_303 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[303*5*5:304*5*5-1]), .o_out_fmap(xor_out[303*24*24*bW:304*24*24*bW-1]));
convchan2 c_2_304 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[304*5*5:305*5*5-1]), .o_out_fmap(xor_out[304*24*24*bW:305*24*24*bW-1]));
convchan2 c_2_305 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[305*5*5:306*5*5-1]), .o_out_fmap(xor_out[305*24*24*bW:306*24*24*bW-1]));
convchan2 c_2_306 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[306*5*5:307*5*5-1]), .o_out_fmap(xor_out[306*24*24*bW:307*24*24*bW-1]));
convchan2 c_2_307 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[307*5*5:308*5*5-1]), .o_out_fmap(xor_out[307*24*24*bW:308*24*24*bW-1]));
convchan2 c_2_308 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[308*5*5:309*5*5-1]), .o_out_fmap(xor_out[308*24*24*bW:309*24*24*bW-1]));
convchan2 c_2_309 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[309*5*5:310*5*5-1]), .o_out_fmap(xor_out[309*24*24*bW:310*24*24*bW-1]));
convchan2 c_2_310 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[310*5*5:311*5*5-1]), .o_out_fmap(xor_out[310*24*24*bW:311*24*24*bW-1]));
convchan2 c_2_311 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[311*5*5:312*5*5-1]), .o_out_fmap(xor_out[311*24*24*bW:312*24*24*bW-1]));
convchan2 c_2_312 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[312*5*5:313*5*5-1]), .o_out_fmap(xor_out[312*24*24*bW:313*24*24*bW-1]));
convchan2 c_2_313 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[313*5*5:314*5*5-1]), .o_out_fmap(xor_out[313*24*24*bW:314*24*24*bW-1]));
convchan2 c_2_314 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[314*5*5:315*5*5-1]), .o_out_fmap(xor_out[314*24*24*bW:315*24*24*bW-1]));
convchan2 c_2_315 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[315*5*5:316*5*5-1]), .o_out_fmap(xor_out[315*24*24*bW:316*24*24*bW-1]));
convchan2 c_2_316 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[316*5*5:317*5*5-1]), .o_out_fmap(xor_out[316*24*24*bW:317*24*24*bW-1]));
convchan2 c_2_317 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[317*5*5:318*5*5-1]), .o_out_fmap(xor_out[317*24*24*bW:318*24*24*bW-1]));
convchan2 c_2_318 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[318*5*5:319*5*5-1]), .o_out_fmap(xor_out[318*24*24*bW:319*24*24*bW-1]));
convchan2 c_2_319 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[319*5*5:320*5*5-1]), .o_out_fmap(xor_out[319*24*24*bW:320*24*24*bW-1]));
convchan2 c_2_320 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[320*5*5:321*5*5-1]), .o_out_fmap(xor_out[320*24*24*bW:321*24*24*bW-1]));
convchan2 c_2_321 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[321*5*5:322*5*5-1]), .o_out_fmap(xor_out[321*24*24*bW:322*24*24*bW-1]));
convchan2 c_2_322 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[322*5*5:323*5*5-1]), .o_out_fmap(xor_out[322*24*24*bW:323*24*24*bW-1]));
convchan2 c_2_323 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[323*5*5:324*5*5-1]), .o_out_fmap(xor_out[323*24*24*bW:324*24*24*bW-1]));
convchan2 c_2_324 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[324*5*5:325*5*5-1]), .o_out_fmap(xor_out[324*24*24*bW:325*24*24*bW-1]));
convchan2 c_2_325 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[325*5*5:326*5*5-1]), .o_out_fmap(xor_out[325*24*24*bW:326*24*24*bW-1]));
convchan2 c_2_326 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[326*5*5:327*5*5-1]), .o_out_fmap(xor_out[326*24*24*bW:327*24*24*bW-1]));
convchan2 c_2_327 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[327*5*5:328*5*5-1]), .o_out_fmap(xor_out[327*24*24*bW:328*24*24*bW-1]));
convchan2 c_2_328 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[328*5*5:329*5*5-1]), .o_out_fmap(xor_out[328*24*24*bW:329*24*24*bW-1]));
convchan2 c_2_329 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[329*5*5:330*5*5-1]), .o_out_fmap(xor_out[329*24*24*bW:330*24*24*bW-1]));
convchan2 c_2_330 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[330*5*5:331*5*5-1]), .o_out_fmap(xor_out[330*24*24*bW:331*24*24*bW-1]));
convchan2 c_2_331 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[331*5*5:332*5*5-1]), .o_out_fmap(xor_out[331*24*24*bW:332*24*24*bW-1]));
convchan2 c_2_332 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[332*5*5:333*5*5-1]), .o_out_fmap(xor_out[332*24*24*bW:333*24*24*bW-1]));
convchan2 c_2_333 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[333*5*5:334*5*5-1]), .o_out_fmap(xor_out[333*24*24*bW:334*24*24*bW-1]));
convchan2 c_2_334 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[334*5*5:335*5*5-1]), .o_out_fmap(xor_out[334*24*24*bW:335*24*24*bW-1]));
convchan2 c_2_335 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[335*5*5:336*5*5-1]), .o_out_fmap(xor_out[335*24*24*bW:336*24*24*bW-1]));
convchan2 c_2_336 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[336*5*5:337*5*5-1]), .o_out_fmap(xor_out[336*24*24*bW:337*24*24*bW-1]));
convchan2 c_2_337 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[337*5*5:338*5*5-1]), .o_out_fmap(xor_out[337*24*24*bW:338*24*24*bW-1]));
convchan2 c_2_338 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[338*5*5:339*5*5-1]), .o_out_fmap(xor_out[338*24*24*bW:339*24*24*bW-1]));
convchan2 c_2_339 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[339*5*5:340*5*5-1]), .o_out_fmap(xor_out[339*24*24*bW:340*24*24*bW-1]));
convchan2 c_2_340 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[340*5*5:341*5*5-1]), .o_out_fmap(xor_out[340*24*24*bW:341*24*24*bW-1]));
convchan2 c_2_341 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[341*5*5:342*5*5-1]), .o_out_fmap(xor_out[341*24*24*bW:342*24*24*bW-1]));
convchan2 c_2_342 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[342*5*5:343*5*5-1]), .o_out_fmap(xor_out[342*24*24*bW:343*24*24*bW-1]));
convchan2 c_2_343 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[343*5*5:344*5*5-1]), .o_out_fmap(xor_out[343*24*24*bW:344*24*24*bW-1]));
convchan2 c_2_344 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[344*5*5:345*5*5-1]), .o_out_fmap(xor_out[344*24*24*bW:345*24*24*bW-1]));
convchan2 c_2_345 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[345*5*5:346*5*5-1]), .o_out_fmap(xor_out[345*24*24*bW:346*24*24*bW-1]));
convchan2 c_2_346 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[346*5*5:347*5*5-1]), .o_out_fmap(xor_out[346*24*24*bW:347*24*24*bW-1]));
convchan2 c_2_347 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[347*5*5:348*5*5-1]), .o_out_fmap(xor_out[347*24*24*bW:348*24*24*bW-1]));
convchan2 c_2_348 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[348*5*5:349*5*5-1]), .o_out_fmap(xor_out[348*24*24*bW:349*24*24*bW-1]));
convchan2 c_2_349 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[349*5*5:350*5*5-1]), .o_out_fmap(xor_out[349*24*24*bW:350*24*24*bW-1]));
convchan2 c_2_350 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[350*5*5:351*5*5-1]), .o_out_fmap(xor_out[350*24*24*bW:351*24*24*bW-1]));
convchan2 c_2_351 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[351*5*5:352*5*5-1]), .o_out_fmap(xor_out[351*24*24*bW:352*24*24*bW-1]));
convchan2 c_2_352 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[352*5*5:353*5*5-1]), .o_out_fmap(xor_out[352*24*24*bW:353*24*24*bW-1]));
convchan2 c_2_353 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[353*5*5:354*5*5-1]), .o_out_fmap(xor_out[353*24*24*bW:354*24*24*bW-1]));
convchan2 c_2_354 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[354*5*5:355*5*5-1]), .o_out_fmap(xor_out[354*24*24*bW:355*24*24*bW-1]));
convchan2 c_2_355 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[355*5*5:356*5*5-1]), .o_out_fmap(xor_out[355*24*24*bW:356*24*24*bW-1]));
convchan2 c_2_356 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[356*5*5:357*5*5-1]), .o_out_fmap(xor_out[356*24*24*bW:357*24*24*bW-1]));
convchan2 c_2_357 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[357*5*5:358*5*5-1]), .o_out_fmap(xor_out[357*24*24*bW:358*24*24*bW-1]));
convchan2 c_2_358 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[358*5*5:359*5*5-1]), .o_out_fmap(xor_out[358*24*24*bW:359*24*24*bW-1]));
convchan2 c_2_359 (.i_image(image[5*12*12:6*12*12*+1]), .i_kernel(kernels[359*5*5:360*5*5-1]), .o_out_fmap(xor_out[359*24*24*bW:360*24*24*bW-1]));
convchan2 c_2_360 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[360*5*5:361*5*5-1]), .o_out_fmap(xor_out[360*24*24*bW:361*24*24*bW-1]));
convchan2 c_2_361 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[361*5*5:362*5*5-1]), .o_out_fmap(xor_out[361*24*24*bW:362*24*24*bW-1]));
convchan2 c_2_362 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[362*5*5:363*5*5-1]), .o_out_fmap(xor_out[362*24*24*bW:363*24*24*bW-1]));
convchan2 c_2_363 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[363*5*5:364*5*5-1]), .o_out_fmap(xor_out[363*24*24*bW:364*24*24*bW-1]));
convchan2 c_2_364 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[364*5*5:365*5*5-1]), .o_out_fmap(xor_out[364*24*24*bW:365*24*24*bW-1]));
convchan2 c_2_365 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[365*5*5:366*5*5-1]), .o_out_fmap(xor_out[365*24*24*bW:366*24*24*bW-1]));
convchan2 c_2_366 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[366*5*5:367*5*5-1]), .o_out_fmap(xor_out[366*24*24*bW:367*24*24*bW-1]));
convchan2 c_2_367 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[367*5*5:368*5*5-1]), .o_out_fmap(xor_out[367*24*24*bW:368*24*24*bW-1]));
convchan2 c_2_368 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[368*5*5:369*5*5-1]), .o_out_fmap(xor_out[368*24*24*bW:369*24*24*bW-1]));
convchan2 c_2_369 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[369*5*5:370*5*5-1]), .o_out_fmap(xor_out[369*24*24*bW:370*24*24*bW-1]));
convchan2 c_2_370 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[370*5*5:371*5*5-1]), .o_out_fmap(xor_out[370*24*24*bW:371*24*24*bW-1]));
convchan2 c_2_371 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[371*5*5:372*5*5-1]), .o_out_fmap(xor_out[371*24*24*bW:372*24*24*bW-1]));
convchan2 c_2_372 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[372*5*5:373*5*5-1]), .o_out_fmap(xor_out[372*24*24*bW:373*24*24*bW-1]));
convchan2 c_2_373 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[373*5*5:374*5*5-1]), .o_out_fmap(xor_out[373*24*24*bW:374*24*24*bW-1]));
convchan2 c_2_374 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[374*5*5:375*5*5-1]), .o_out_fmap(xor_out[374*24*24*bW:375*24*24*bW-1]));
convchan2 c_2_375 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[375*5*5:376*5*5-1]), .o_out_fmap(xor_out[375*24*24*bW:376*24*24*bW-1]));
convchan2 c_2_376 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[376*5*5:377*5*5-1]), .o_out_fmap(xor_out[376*24*24*bW:377*24*24*bW-1]));
convchan2 c_2_377 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[377*5*5:378*5*5-1]), .o_out_fmap(xor_out[377*24*24*bW:378*24*24*bW-1]));
convchan2 c_2_378 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[378*5*5:379*5*5-1]), .o_out_fmap(xor_out[378*24*24*bW:379*24*24*bW-1]));
convchan2 c_2_379 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[379*5*5:380*5*5-1]), .o_out_fmap(xor_out[379*24*24*bW:380*24*24*bW-1]));
convchan2 c_2_380 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[380*5*5:381*5*5-1]), .o_out_fmap(xor_out[380*24*24*bW:381*24*24*bW-1]));
convchan2 c_2_381 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[381*5*5:382*5*5-1]), .o_out_fmap(xor_out[381*24*24*bW:382*24*24*bW-1]));
convchan2 c_2_382 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[382*5*5:383*5*5-1]), .o_out_fmap(xor_out[382*24*24*bW:383*24*24*bW-1]));
convchan2 c_2_383 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[383*5*5:384*5*5-1]), .o_out_fmap(xor_out[383*24*24*bW:384*24*24*bW-1]));
convchan2 c_2_384 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[384*5*5:385*5*5-1]), .o_out_fmap(xor_out[384*24*24*bW:385*24*24*bW-1]));
convchan2 c_2_385 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[385*5*5:386*5*5-1]), .o_out_fmap(xor_out[385*24*24*bW:386*24*24*bW-1]));
convchan2 c_2_386 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[386*5*5:387*5*5-1]), .o_out_fmap(xor_out[386*24*24*bW:387*24*24*bW-1]));
convchan2 c_2_387 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[387*5*5:388*5*5-1]), .o_out_fmap(xor_out[387*24*24*bW:388*24*24*bW-1]));
convchan2 c_2_388 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[388*5*5:389*5*5-1]), .o_out_fmap(xor_out[388*24*24*bW:389*24*24*bW-1]));
convchan2 c_2_389 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[389*5*5:390*5*5-1]), .o_out_fmap(xor_out[389*24*24*bW:390*24*24*bW-1]));
convchan2 c_2_390 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[390*5*5:391*5*5-1]), .o_out_fmap(xor_out[390*24*24*bW:391*24*24*bW-1]));
convchan2 c_2_391 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[391*5*5:392*5*5-1]), .o_out_fmap(xor_out[391*24*24*bW:392*24*24*bW-1]));
convchan2 c_2_392 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[392*5*5:393*5*5-1]), .o_out_fmap(xor_out[392*24*24*bW:393*24*24*bW-1]));
convchan2 c_2_393 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[393*5*5:394*5*5-1]), .o_out_fmap(xor_out[393*24*24*bW:394*24*24*bW-1]));
convchan2 c_2_394 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[394*5*5:395*5*5-1]), .o_out_fmap(xor_out[394*24*24*bW:395*24*24*bW-1]));
convchan2 c_2_395 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[395*5*5:396*5*5-1]), .o_out_fmap(xor_out[395*24*24*bW:396*24*24*bW-1]));
convchan2 c_2_396 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[396*5*5:397*5*5-1]), .o_out_fmap(xor_out[396*24*24*bW:397*24*24*bW-1]));
convchan2 c_2_397 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[397*5*5:398*5*5-1]), .o_out_fmap(xor_out[397*24*24*bW:398*24*24*bW-1]));
convchan2 c_2_398 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[398*5*5:399*5*5-1]), .o_out_fmap(xor_out[398*24*24*bW:399*24*24*bW-1]));
convchan2 c_2_399 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[399*5*5:400*5*5-1]), .o_out_fmap(xor_out[399*24*24*bW:400*24*24*bW-1]));
convchan2 c_2_400 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[400*5*5:401*5*5-1]), .o_out_fmap(xor_out[400*24*24*bW:401*24*24*bW-1]));
convchan2 c_2_401 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[401*5*5:402*5*5-1]), .o_out_fmap(xor_out[401*24*24*bW:402*24*24*bW-1]));
convchan2 c_2_402 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[402*5*5:403*5*5-1]), .o_out_fmap(xor_out[402*24*24*bW:403*24*24*bW-1]));
convchan2 c_2_403 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[403*5*5:404*5*5-1]), .o_out_fmap(xor_out[403*24*24*bW:404*24*24*bW-1]));
convchan2 c_2_404 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[404*5*5:405*5*5-1]), .o_out_fmap(xor_out[404*24*24*bW:405*24*24*bW-1]));
convchan2 c_2_405 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[405*5*5:406*5*5-1]), .o_out_fmap(xor_out[405*24*24*bW:406*24*24*bW-1]));
convchan2 c_2_406 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[406*5*5:407*5*5-1]), .o_out_fmap(xor_out[406*24*24*bW:407*24*24*bW-1]));
convchan2 c_2_407 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[407*5*5:408*5*5-1]), .o_out_fmap(xor_out[407*24*24*bW:408*24*24*bW-1]));
convchan2 c_2_408 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[408*5*5:409*5*5-1]), .o_out_fmap(xor_out[408*24*24*bW:409*24*24*bW-1]));
convchan2 c_2_409 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[409*5*5:410*5*5-1]), .o_out_fmap(xor_out[409*24*24*bW:410*24*24*bW-1]));
convchan2 c_2_410 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[410*5*5:411*5*5-1]), .o_out_fmap(xor_out[410*24*24*bW:411*24*24*bW-1]));
convchan2 c_2_411 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[411*5*5:412*5*5-1]), .o_out_fmap(xor_out[411*24*24*bW:412*24*24*bW-1]));
convchan2 c_2_412 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[412*5*5:413*5*5-1]), .o_out_fmap(xor_out[412*24*24*bW:413*24*24*bW-1]));
convchan2 c_2_413 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[413*5*5:414*5*5-1]), .o_out_fmap(xor_out[413*24*24*bW:414*24*24*bW-1]));
convchan2 c_2_414 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[414*5*5:415*5*5-1]), .o_out_fmap(xor_out[414*24*24*bW:415*24*24*bW-1]));
convchan2 c_2_415 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[415*5*5:416*5*5-1]), .o_out_fmap(xor_out[415*24*24*bW:416*24*24*bW-1]));
convchan2 c_2_416 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[416*5*5:417*5*5-1]), .o_out_fmap(xor_out[416*24*24*bW:417*24*24*bW-1]));
convchan2 c_2_417 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[417*5*5:418*5*5-1]), .o_out_fmap(xor_out[417*24*24*bW:418*24*24*bW-1]));
convchan2 c_2_418 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[418*5*5:419*5*5-1]), .o_out_fmap(xor_out[418*24*24*bW:419*24*24*bW-1]));
convchan2 c_2_419 (.i_image(image[6*12*12:7*12*12*+1]), .i_kernel(kernels[419*5*5:420*5*5-1]), .o_out_fmap(xor_out[419*24*24*bW:420*24*24*bW-1]));
convchan2 c_2_420 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[420*5*5:421*5*5-1]), .o_out_fmap(xor_out[420*24*24*bW:421*24*24*bW-1]));
convchan2 c_2_421 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[421*5*5:422*5*5-1]), .o_out_fmap(xor_out[421*24*24*bW:422*24*24*bW-1]));
convchan2 c_2_422 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[422*5*5:423*5*5-1]), .o_out_fmap(xor_out[422*24*24*bW:423*24*24*bW-1]));
convchan2 c_2_423 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[423*5*5:424*5*5-1]), .o_out_fmap(xor_out[423*24*24*bW:424*24*24*bW-1]));
convchan2 c_2_424 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[424*5*5:425*5*5-1]), .o_out_fmap(xor_out[424*24*24*bW:425*24*24*bW-1]));
convchan2 c_2_425 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[425*5*5:426*5*5-1]), .o_out_fmap(xor_out[425*24*24*bW:426*24*24*bW-1]));
convchan2 c_2_426 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[426*5*5:427*5*5-1]), .o_out_fmap(xor_out[426*24*24*bW:427*24*24*bW-1]));
convchan2 c_2_427 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[427*5*5:428*5*5-1]), .o_out_fmap(xor_out[427*24*24*bW:428*24*24*bW-1]));
convchan2 c_2_428 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[428*5*5:429*5*5-1]), .o_out_fmap(xor_out[428*24*24*bW:429*24*24*bW-1]));
convchan2 c_2_429 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[429*5*5:430*5*5-1]), .o_out_fmap(xor_out[429*24*24*bW:430*24*24*bW-1]));
convchan2 c_2_430 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[430*5*5:431*5*5-1]), .o_out_fmap(xor_out[430*24*24*bW:431*24*24*bW-1]));
convchan2 c_2_431 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[431*5*5:432*5*5-1]), .o_out_fmap(xor_out[431*24*24*bW:432*24*24*bW-1]));
convchan2 c_2_432 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[432*5*5:433*5*5-1]), .o_out_fmap(xor_out[432*24*24*bW:433*24*24*bW-1]));
convchan2 c_2_433 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[433*5*5:434*5*5-1]), .o_out_fmap(xor_out[433*24*24*bW:434*24*24*bW-1]));
convchan2 c_2_434 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[434*5*5:435*5*5-1]), .o_out_fmap(xor_out[434*24*24*bW:435*24*24*bW-1]));
convchan2 c_2_435 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[435*5*5:436*5*5-1]), .o_out_fmap(xor_out[435*24*24*bW:436*24*24*bW-1]));
convchan2 c_2_436 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[436*5*5:437*5*5-1]), .o_out_fmap(xor_out[436*24*24*bW:437*24*24*bW-1]));
convchan2 c_2_437 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[437*5*5:438*5*5-1]), .o_out_fmap(xor_out[437*24*24*bW:438*24*24*bW-1]));
convchan2 c_2_438 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[438*5*5:439*5*5-1]), .o_out_fmap(xor_out[438*24*24*bW:439*24*24*bW-1]));
convchan2 c_2_439 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[439*5*5:440*5*5-1]), .o_out_fmap(xor_out[439*24*24*bW:440*24*24*bW-1]));
convchan2 c_2_440 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[440*5*5:441*5*5-1]), .o_out_fmap(xor_out[440*24*24*bW:441*24*24*bW-1]));
convchan2 c_2_441 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[441*5*5:442*5*5-1]), .o_out_fmap(xor_out[441*24*24*bW:442*24*24*bW-1]));
convchan2 c_2_442 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[442*5*5:443*5*5-1]), .o_out_fmap(xor_out[442*24*24*bW:443*24*24*bW-1]));
convchan2 c_2_443 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[443*5*5:444*5*5-1]), .o_out_fmap(xor_out[443*24*24*bW:444*24*24*bW-1]));
convchan2 c_2_444 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[444*5*5:445*5*5-1]), .o_out_fmap(xor_out[444*24*24*bW:445*24*24*bW-1]));
convchan2 c_2_445 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[445*5*5:446*5*5-1]), .o_out_fmap(xor_out[445*24*24*bW:446*24*24*bW-1]));
convchan2 c_2_446 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[446*5*5:447*5*5-1]), .o_out_fmap(xor_out[446*24*24*bW:447*24*24*bW-1]));
convchan2 c_2_447 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[447*5*5:448*5*5-1]), .o_out_fmap(xor_out[447*24*24*bW:448*24*24*bW-1]));
convchan2 c_2_448 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[448*5*5:449*5*5-1]), .o_out_fmap(xor_out[448*24*24*bW:449*24*24*bW-1]));
convchan2 c_2_449 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[449*5*5:450*5*5-1]), .o_out_fmap(xor_out[449*24*24*bW:450*24*24*bW-1]));
convchan2 c_2_450 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[450*5*5:451*5*5-1]), .o_out_fmap(xor_out[450*24*24*bW:451*24*24*bW-1]));
convchan2 c_2_451 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[451*5*5:452*5*5-1]), .o_out_fmap(xor_out[451*24*24*bW:452*24*24*bW-1]));
convchan2 c_2_452 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[452*5*5:453*5*5-1]), .o_out_fmap(xor_out[452*24*24*bW:453*24*24*bW-1]));
convchan2 c_2_453 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[453*5*5:454*5*5-1]), .o_out_fmap(xor_out[453*24*24*bW:454*24*24*bW-1]));
convchan2 c_2_454 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[454*5*5:455*5*5-1]), .o_out_fmap(xor_out[454*24*24*bW:455*24*24*bW-1]));
convchan2 c_2_455 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[455*5*5:456*5*5-1]), .o_out_fmap(xor_out[455*24*24*bW:456*24*24*bW-1]));
convchan2 c_2_456 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[456*5*5:457*5*5-1]), .o_out_fmap(xor_out[456*24*24*bW:457*24*24*bW-1]));
convchan2 c_2_457 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[457*5*5:458*5*5-1]), .o_out_fmap(xor_out[457*24*24*bW:458*24*24*bW-1]));
convchan2 c_2_458 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[458*5*5:459*5*5-1]), .o_out_fmap(xor_out[458*24*24*bW:459*24*24*bW-1]));
convchan2 c_2_459 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[459*5*5:460*5*5-1]), .o_out_fmap(xor_out[459*24*24*bW:460*24*24*bW-1]));
convchan2 c_2_460 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[460*5*5:461*5*5-1]), .o_out_fmap(xor_out[460*24*24*bW:461*24*24*bW-1]));
convchan2 c_2_461 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[461*5*5:462*5*5-1]), .o_out_fmap(xor_out[461*24*24*bW:462*24*24*bW-1]));
convchan2 c_2_462 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[462*5*5:463*5*5-1]), .o_out_fmap(xor_out[462*24*24*bW:463*24*24*bW-1]));
convchan2 c_2_463 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[463*5*5:464*5*5-1]), .o_out_fmap(xor_out[463*24*24*bW:464*24*24*bW-1]));
convchan2 c_2_464 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[464*5*5:465*5*5-1]), .o_out_fmap(xor_out[464*24*24*bW:465*24*24*bW-1]));
convchan2 c_2_465 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[465*5*5:466*5*5-1]), .o_out_fmap(xor_out[465*24*24*bW:466*24*24*bW-1]));
convchan2 c_2_466 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[466*5*5:467*5*5-1]), .o_out_fmap(xor_out[466*24*24*bW:467*24*24*bW-1]));
convchan2 c_2_467 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[467*5*5:468*5*5-1]), .o_out_fmap(xor_out[467*24*24*bW:468*24*24*bW-1]));
convchan2 c_2_468 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[468*5*5:469*5*5-1]), .o_out_fmap(xor_out[468*24*24*bW:469*24*24*bW-1]));
convchan2 c_2_469 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[469*5*5:470*5*5-1]), .o_out_fmap(xor_out[469*24*24*bW:470*24*24*bW-1]));
convchan2 c_2_470 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[470*5*5:471*5*5-1]), .o_out_fmap(xor_out[470*24*24*bW:471*24*24*bW-1]));
convchan2 c_2_471 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[471*5*5:472*5*5-1]), .o_out_fmap(xor_out[471*24*24*bW:472*24*24*bW-1]));
convchan2 c_2_472 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[472*5*5:473*5*5-1]), .o_out_fmap(xor_out[472*24*24*bW:473*24*24*bW-1]));
convchan2 c_2_473 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[473*5*5:474*5*5-1]), .o_out_fmap(xor_out[473*24*24*bW:474*24*24*bW-1]));
convchan2 c_2_474 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[474*5*5:475*5*5-1]), .o_out_fmap(xor_out[474*24*24*bW:475*24*24*bW-1]));
convchan2 c_2_475 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[475*5*5:476*5*5-1]), .o_out_fmap(xor_out[475*24*24*bW:476*24*24*bW-1]));
convchan2 c_2_476 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[476*5*5:477*5*5-1]), .o_out_fmap(xor_out[476*24*24*bW:477*24*24*bW-1]));
convchan2 c_2_477 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[477*5*5:478*5*5-1]), .o_out_fmap(xor_out[477*24*24*bW:478*24*24*bW-1]));
convchan2 c_2_478 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[478*5*5:479*5*5-1]), .o_out_fmap(xor_out[478*24*24*bW:479*24*24*bW-1]));
convchan2 c_2_479 (.i_image(image[7*12*12:8*12*12*+1]), .i_kernel(kernels[479*5*5:480*5*5-1]), .o_out_fmap(xor_out[479*24*24*bW:480*24*24*bW-1]));
convchan2 c_2_480 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[480*5*5:481*5*5-1]), .o_out_fmap(xor_out[480*24*24*bW:481*24*24*bW-1]));
convchan2 c_2_481 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[481*5*5:482*5*5-1]), .o_out_fmap(xor_out[481*24*24*bW:482*24*24*bW-1]));
convchan2 c_2_482 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[482*5*5:483*5*5-1]), .o_out_fmap(xor_out[482*24*24*bW:483*24*24*bW-1]));
convchan2 c_2_483 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[483*5*5:484*5*5-1]), .o_out_fmap(xor_out[483*24*24*bW:484*24*24*bW-1]));
convchan2 c_2_484 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[484*5*5:485*5*5-1]), .o_out_fmap(xor_out[484*24*24*bW:485*24*24*bW-1]));
convchan2 c_2_485 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[485*5*5:486*5*5-1]), .o_out_fmap(xor_out[485*24*24*bW:486*24*24*bW-1]));
convchan2 c_2_486 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[486*5*5:487*5*5-1]), .o_out_fmap(xor_out[486*24*24*bW:487*24*24*bW-1]));
convchan2 c_2_487 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[487*5*5:488*5*5-1]), .o_out_fmap(xor_out[487*24*24*bW:488*24*24*bW-1]));
convchan2 c_2_488 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[488*5*5:489*5*5-1]), .o_out_fmap(xor_out[488*24*24*bW:489*24*24*bW-1]));
convchan2 c_2_489 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[489*5*5:490*5*5-1]), .o_out_fmap(xor_out[489*24*24*bW:490*24*24*bW-1]));
convchan2 c_2_490 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[490*5*5:491*5*5-1]), .o_out_fmap(xor_out[490*24*24*bW:491*24*24*bW-1]));
convchan2 c_2_491 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[491*5*5:492*5*5-1]), .o_out_fmap(xor_out[491*24*24*bW:492*24*24*bW-1]));
convchan2 c_2_492 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[492*5*5:493*5*5-1]), .o_out_fmap(xor_out[492*24*24*bW:493*24*24*bW-1]));
convchan2 c_2_493 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[493*5*5:494*5*5-1]), .o_out_fmap(xor_out[493*24*24*bW:494*24*24*bW-1]));
convchan2 c_2_494 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[494*5*5:495*5*5-1]), .o_out_fmap(xor_out[494*24*24*bW:495*24*24*bW-1]));
convchan2 c_2_495 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[495*5*5:496*5*5-1]), .o_out_fmap(xor_out[495*24*24*bW:496*24*24*bW-1]));
convchan2 c_2_496 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[496*5*5:497*5*5-1]), .o_out_fmap(xor_out[496*24*24*bW:497*24*24*bW-1]));
convchan2 c_2_497 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[497*5*5:498*5*5-1]), .o_out_fmap(xor_out[497*24*24*bW:498*24*24*bW-1]));
convchan2 c_2_498 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[498*5*5:499*5*5-1]), .o_out_fmap(xor_out[498*24*24*bW:499*24*24*bW-1]));
convchan2 c_2_499 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[499*5*5:500*5*5-1]), .o_out_fmap(xor_out[499*24*24*bW:500*24*24*bW-1]));
convchan2 c_2_500 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[500*5*5:501*5*5-1]), .o_out_fmap(xor_out[500*24*24*bW:501*24*24*bW-1]));
convchan2 c_2_501 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[501*5*5:502*5*5-1]), .o_out_fmap(xor_out[501*24*24*bW:502*24*24*bW-1]));
convchan2 c_2_502 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[502*5*5:503*5*5-1]), .o_out_fmap(xor_out[502*24*24*bW:503*24*24*bW-1]));
convchan2 c_2_503 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[503*5*5:504*5*5-1]), .o_out_fmap(xor_out[503*24*24*bW:504*24*24*bW-1]));
convchan2 c_2_504 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[504*5*5:505*5*5-1]), .o_out_fmap(xor_out[504*24*24*bW:505*24*24*bW-1]));
convchan2 c_2_505 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[505*5*5:506*5*5-1]), .o_out_fmap(xor_out[505*24*24*bW:506*24*24*bW-1]));
convchan2 c_2_506 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[506*5*5:507*5*5-1]), .o_out_fmap(xor_out[506*24*24*bW:507*24*24*bW-1]));
convchan2 c_2_507 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[507*5*5:508*5*5-1]), .o_out_fmap(xor_out[507*24*24*bW:508*24*24*bW-1]));
convchan2 c_2_508 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[508*5*5:509*5*5-1]), .o_out_fmap(xor_out[508*24*24*bW:509*24*24*bW-1]));
convchan2 c_2_509 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[509*5*5:510*5*5-1]), .o_out_fmap(xor_out[509*24*24*bW:510*24*24*bW-1]));
convchan2 c_2_510 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[510*5*5:511*5*5-1]), .o_out_fmap(xor_out[510*24*24*bW:511*24*24*bW-1]));
convchan2 c_2_511 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[511*5*5:512*5*5-1]), .o_out_fmap(xor_out[511*24*24*bW:512*24*24*bW-1]));
convchan2 c_2_512 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[512*5*5:513*5*5-1]), .o_out_fmap(xor_out[512*24*24*bW:513*24*24*bW-1]));
convchan2 c_2_513 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[513*5*5:514*5*5-1]), .o_out_fmap(xor_out[513*24*24*bW:514*24*24*bW-1]));
convchan2 c_2_514 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[514*5*5:515*5*5-1]), .o_out_fmap(xor_out[514*24*24*bW:515*24*24*bW-1]));
convchan2 c_2_515 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[515*5*5:516*5*5-1]), .o_out_fmap(xor_out[515*24*24*bW:516*24*24*bW-1]));
convchan2 c_2_516 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[516*5*5:517*5*5-1]), .o_out_fmap(xor_out[516*24*24*bW:517*24*24*bW-1]));
convchan2 c_2_517 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[517*5*5:518*5*5-1]), .o_out_fmap(xor_out[517*24*24*bW:518*24*24*bW-1]));
convchan2 c_2_518 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[518*5*5:519*5*5-1]), .o_out_fmap(xor_out[518*24*24*bW:519*24*24*bW-1]));
convchan2 c_2_519 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[519*5*5:520*5*5-1]), .o_out_fmap(xor_out[519*24*24*bW:520*24*24*bW-1]));
convchan2 c_2_520 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[520*5*5:521*5*5-1]), .o_out_fmap(xor_out[520*24*24*bW:521*24*24*bW-1]));
convchan2 c_2_521 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[521*5*5:522*5*5-1]), .o_out_fmap(xor_out[521*24*24*bW:522*24*24*bW-1]));
convchan2 c_2_522 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[522*5*5:523*5*5-1]), .o_out_fmap(xor_out[522*24*24*bW:523*24*24*bW-1]));
convchan2 c_2_523 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[523*5*5:524*5*5-1]), .o_out_fmap(xor_out[523*24*24*bW:524*24*24*bW-1]));
convchan2 c_2_524 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[524*5*5:525*5*5-1]), .o_out_fmap(xor_out[524*24*24*bW:525*24*24*bW-1]));
convchan2 c_2_525 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[525*5*5:526*5*5-1]), .o_out_fmap(xor_out[525*24*24*bW:526*24*24*bW-1]));
convchan2 c_2_526 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[526*5*5:527*5*5-1]), .o_out_fmap(xor_out[526*24*24*bW:527*24*24*bW-1]));
convchan2 c_2_527 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[527*5*5:528*5*5-1]), .o_out_fmap(xor_out[527*24*24*bW:528*24*24*bW-1]));
convchan2 c_2_528 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[528*5*5:529*5*5-1]), .o_out_fmap(xor_out[528*24*24*bW:529*24*24*bW-1]));
convchan2 c_2_529 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[529*5*5:530*5*5-1]), .o_out_fmap(xor_out[529*24*24*bW:530*24*24*bW-1]));
convchan2 c_2_530 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[530*5*5:531*5*5-1]), .o_out_fmap(xor_out[530*24*24*bW:531*24*24*bW-1]));
convchan2 c_2_531 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[531*5*5:532*5*5-1]), .o_out_fmap(xor_out[531*24*24*bW:532*24*24*bW-1]));
convchan2 c_2_532 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[532*5*5:533*5*5-1]), .o_out_fmap(xor_out[532*24*24*bW:533*24*24*bW-1]));
convchan2 c_2_533 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[533*5*5:534*5*5-1]), .o_out_fmap(xor_out[533*24*24*bW:534*24*24*bW-1]));
convchan2 c_2_534 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[534*5*5:535*5*5-1]), .o_out_fmap(xor_out[534*24*24*bW:535*24*24*bW-1]));
convchan2 c_2_535 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[535*5*5:536*5*5-1]), .o_out_fmap(xor_out[535*24*24*bW:536*24*24*bW-1]));
convchan2 c_2_536 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[536*5*5:537*5*5-1]), .o_out_fmap(xor_out[536*24*24*bW:537*24*24*bW-1]));
convchan2 c_2_537 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[537*5*5:538*5*5-1]), .o_out_fmap(xor_out[537*24*24*bW:538*24*24*bW-1]));
convchan2 c_2_538 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[538*5*5:539*5*5-1]), .o_out_fmap(xor_out[538*24*24*bW:539*24*24*bW-1]));
convchan2 c_2_539 (.i_image(image[8*12*12:9*12*12*+1]), .i_kernel(kernels[539*5*5:540*5*5-1]), .o_out_fmap(xor_out[539*24*24*bW:540*24*24*bW-1]));
convchan2 c_2_540 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[540*5*5:541*5*5-1]), .o_out_fmap(xor_out[540*24*24*bW:541*24*24*bW-1]));
convchan2 c_2_541 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[541*5*5:542*5*5-1]), .o_out_fmap(xor_out[541*24*24*bW:542*24*24*bW-1]));
convchan2 c_2_542 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[542*5*5:543*5*5-1]), .o_out_fmap(xor_out[542*24*24*bW:543*24*24*bW-1]));
convchan2 c_2_543 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[543*5*5:544*5*5-1]), .o_out_fmap(xor_out[543*24*24*bW:544*24*24*bW-1]));
convchan2 c_2_544 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[544*5*5:545*5*5-1]), .o_out_fmap(xor_out[544*24*24*bW:545*24*24*bW-1]));
convchan2 c_2_545 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[545*5*5:546*5*5-1]), .o_out_fmap(xor_out[545*24*24*bW:546*24*24*bW-1]));
convchan2 c_2_546 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[546*5*5:547*5*5-1]), .o_out_fmap(xor_out[546*24*24*bW:547*24*24*bW-1]));
convchan2 c_2_547 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[547*5*5:548*5*5-1]), .o_out_fmap(xor_out[547*24*24*bW:548*24*24*bW-1]));
convchan2 c_2_548 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[548*5*5:549*5*5-1]), .o_out_fmap(xor_out[548*24*24*bW:549*24*24*bW-1]));
convchan2 c_2_549 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[549*5*5:550*5*5-1]), .o_out_fmap(xor_out[549*24*24*bW:550*24*24*bW-1]));
convchan2 c_2_550 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[550*5*5:551*5*5-1]), .o_out_fmap(xor_out[550*24*24*bW:551*24*24*bW-1]));
convchan2 c_2_551 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[551*5*5:552*5*5-1]), .o_out_fmap(xor_out[551*24*24*bW:552*24*24*bW-1]));
convchan2 c_2_552 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[552*5*5:553*5*5-1]), .o_out_fmap(xor_out[552*24*24*bW:553*24*24*bW-1]));
convchan2 c_2_553 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[553*5*5:554*5*5-1]), .o_out_fmap(xor_out[553*24*24*bW:554*24*24*bW-1]));
convchan2 c_2_554 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[554*5*5:555*5*5-1]), .o_out_fmap(xor_out[554*24*24*bW:555*24*24*bW-1]));
convchan2 c_2_555 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[555*5*5:556*5*5-1]), .o_out_fmap(xor_out[555*24*24*bW:556*24*24*bW-1]));
convchan2 c_2_556 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[556*5*5:557*5*5-1]), .o_out_fmap(xor_out[556*24*24*bW:557*24*24*bW-1]));
convchan2 c_2_557 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[557*5*5:558*5*5-1]), .o_out_fmap(xor_out[557*24*24*bW:558*24*24*bW-1]));
convchan2 c_2_558 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[558*5*5:559*5*5-1]), .o_out_fmap(xor_out[558*24*24*bW:559*24*24*bW-1]));
convchan2 c_2_559 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[559*5*5:560*5*5-1]), .o_out_fmap(xor_out[559*24*24*bW:560*24*24*bW-1]));
convchan2 c_2_560 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[560*5*5:561*5*5-1]), .o_out_fmap(xor_out[560*24*24*bW:561*24*24*bW-1]));
convchan2 c_2_561 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[561*5*5:562*5*5-1]), .o_out_fmap(xor_out[561*24*24*bW:562*24*24*bW-1]));
convchan2 c_2_562 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[562*5*5:563*5*5-1]), .o_out_fmap(xor_out[562*24*24*bW:563*24*24*bW-1]));
convchan2 c_2_563 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[563*5*5:564*5*5-1]), .o_out_fmap(xor_out[563*24*24*bW:564*24*24*bW-1]));
convchan2 c_2_564 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[564*5*5:565*5*5-1]), .o_out_fmap(xor_out[564*24*24*bW:565*24*24*bW-1]));
convchan2 c_2_565 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[565*5*5:566*5*5-1]), .o_out_fmap(xor_out[565*24*24*bW:566*24*24*bW-1]));
convchan2 c_2_566 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[566*5*5:567*5*5-1]), .o_out_fmap(xor_out[566*24*24*bW:567*24*24*bW-1]));
convchan2 c_2_567 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[567*5*5:568*5*5-1]), .o_out_fmap(xor_out[567*24*24*bW:568*24*24*bW-1]));
convchan2 c_2_568 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[568*5*5:569*5*5-1]), .o_out_fmap(xor_out[568*24*24*bW:569*24*24*bW-1]));
convchan2 c_2_569 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[569*5*5:570*5*5-1]), .o_out_fmap(xor_out[569*24*24*bW:570*24*24*bW-1]));
convchan2 c_2_570 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[570*5*5:571*5*5-1]), .o_out_fmap(xor_out[570*24*24*bW:571*24*24*bW-1]));
convchan2 c_2_571 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[571*5*5:572*5*5-1]), .o_out_fmap(xor_out[571*24*24*bW:572*24*24*bW-1]));
convchan2 c_2_572 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[572*5*5:573*5*5-1]), .o_out_fmap(xor_out[572*24*24*bW:573*24*24*bW-1]));
convchan2 c_2_573 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[573*5*5:574*5*5-1]), .o_out_fmap(xor_out[573*24*24*bW:574*24*24*bW-1]));
convchan2 c_2_574 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[574*5*5:575*5*5-1]), .o_out_fmap(xor_out[574*24*24*bW:575*24*24*bW-1]));
convchan2 c_2_575 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[575*5*5:576*5*5-1]), .o_out_fmap(xor_out[575*24*24*bW:576*24*24*bW-1]));
convchan2 c_2_576 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[576*5*5:577*5*5-1]), .o_out_fmap(xor_out[576*24*24*bW:577*24*24*bW-1]));
convchan2 c_2_577 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[577*5*5:578*5*5-1]), .o_out_fmap(xor_out[577*24*24*bW:578*24*24*bW-1]));
convchan2 c_2_578 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[578*5*5:579*5*5-1]), .o_out_fmap(xor_out[578*24*24*bW:579*24*24*bW-1]));
convchan2 c_2_579 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[579*5*5:580*5*5-1]), .o_out_fmap(xor_out[579*24*24*bW:580*24*24*bW-1]));
convchan2 c_2_580 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[580*5*5:581*5*5-1]), .o_out_fmap(xor_out[580*24*24*bW:581*24*24*bW-1]));
convchan2 c_2_581 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[581*5*5:582*5*5-1]), .o_out_fmap(xor_out[581*24*24*bW:582*24*24*bW-1]));
convchan2 c_2_582 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[582*5*5:583*5*5-1]), .o_out_fmap(xor_out[582*24*24*bW:583*24*24*bW-1]));
convchan2 c_2_583 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[583*5*5:584*5*5-1]), .o_out_fmap(xor_out[583*24*24*bW:584*24*24*bW-1]));
convchan2 c_2_584 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[584*5*5:585*5*5-1]), .o_out_fmap(xor_out[584*24*24*bW:585*24*24*bW-1]));
convchan2 c_2_585 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[585*5*5:586*5*5-1]), .o_out_fmap(xor_out[585*24*24*bW:586*24*24*bW-1]));
convchan2 c_2_586 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[586*5*5:587*5*5-1]), .o_out_fmap(xor_out[586*24*24*bW:587*24*24*bW-1]));
convchan2 c_2_587 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[587*5*5:588*5*5-1]), .o_out_fmap(xor_out[587*24*24*bW:588*24*24*bW-1]));
convchan2 c_2_588 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[588*5*5:589*5*5-1]), .o_out_fmap(xor_out[588*24*24*bW:589*24*24*bW-1]));
convchan2 c_2_589 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[589*5*5:590*5*5-1]), .o_out_fmap(xor_out[589*24*24*bW:590*24*24*bW-1]));
convchan2 c_2_590 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[590*5*5:591*5*5-1]), .o_out_fmap(xor_out[590*24*24*bW:591*24*24*bW-1]));
convchan2 c_2_591 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[591*5*5:592*5*5-1]), .o_out_fmap(xor_out[591*24*24*bW:592*24*24*bW-1]));
convchan2 c_2_592 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[592*5*5:593*5*5-1]), .o_out_fmap(xor_out[592*24*24*bW:593*24*24*bW-1]));
convchan2 c_2_593 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[593*5*5:594*5*5-1]), .o_out_fmap(xor_out[593*24*24*bW:594*24*24*bW-1]));
convchan2 c_2_594 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[594*5*5:595*5*5-1]), .o_out_fmap(xor_out[594*24*24*bW:595*24*24*bW-1]));
convchan2 c_2_595 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[595*5*5:596*5*5-1]), .o_out_fmap(xor_out[595*24*24*bW:596*24*24*bW-1]));
convchan2 c_2_596 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[596*5*5:597*5*5-1]), .o_out_fmap(xor_out[596*24*24*bW:597*24*24*bW-1]));
convchan2 c_2_597 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[597*5*5:598*5*5-1]), .o_out_fmap(xor_out[597*24*24*bW:598*24*24*bW-1]));
convchan2 c_2_598 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[598*5*5:599*5*5-1]), .o_out_fmap(xor_out[598*24*24*bW:599*24*24*bW-1]));
convchan2 c_2_599 (.i_image(image[9*12*12:10*12*12*+1]), .i_kernel(kernels[599*5*5:600*5*5-1]), .o_out_fmap(xor_out[599*24*24*bW:600*24*24*bW-1]));
convchan2 c_2_600 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[600*5*5:601*5*5-1]), .o_out_fmap(xor_out[600*24*24*bW:601*24*24*bW-1]));
convchan2 c_2_601 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[601*5*5:602*5*5-1]), .o_out_fmap(xor_out[601*24*24*bW:602*24*24*bW-1]));
convchan2 c_2_602 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[602*5*5:603*5*5-1]), .o_out_fmap(xor_out[602*24*24*bW:603*24*24*bW-1]));
convchan2 c_2_603 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[603*5*5:604*5*5-1]), .o_out_fmap(xor_out[603*24*24*bW:604*24*24*bW-1]));
convchan2 c_2_604 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[604*5*5:605*5*5-1]), .o_out_fmap(xor_out[604*24*24*bW:605*24*24*bW-1]));
convchan2 c_2_605 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[605*5*5:606*5*5-1]), .o_out_fmap(xor_out[605*24*24*bW:606*24*24*bW-1]));
convchan2 c_2_606 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[606*5*5:607*5*5-1]), .o_out_fmap(xor_out[606*24*24*bW:607*24*24*bW-1]));
convchan2 c_2_607 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[607*5*5:608*5*5-1]), .o_out_fmap(xor_out[607*24*24*bW:608*24*24*bW-1]));
convchan2 c_2_608 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[608*5*5:609*5*5-1]), .o_out_fmap(xor_out[608*24*24*bW:609*24*24*bW-1]));
convchan2 c_2_609 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[609*5*5:610*5*5-1]), .o_out_fmap(xor_out[609*24*24*bW:610*24*24*bW-1]));
convchan2 c_2_610 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[610*5*5:611*5*5-1]), .o_out_fmap(xor_out[610*24*24*bW:611*24*24*bW-1]));
convchan2 c_2_611 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[611*5*5:612*5*5-1]), .o_out_fmap(xor_out[611*24*24*bW:612*24*24*bW-1]));
convchan2 c_2_612 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[612*5*5:613*5*5-1]), .o_out_fmap(xor_out[612*24*24*bW:613*24*24*bW-1]));
convchan2 c_2_613 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[613*5*5:614*5*5-1]), .o_out_fmap(xor_out[613*24*24*bW:614*24*24*bW-1]));
convchan2 c_2_614 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[614*5*5:615*5*5-1]), .o_out_fmap(xor_out[614*24*24*bW:615*24*24*bW-1]));
convchan2 c_2_615 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[615*5*5:616*5*5-1]), .o_out_fmap(xor_out[615*24*24*bW:616*24*24*bW-1]));
convchan2 c_2_616 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[616*5*5:617*5*5-1]), .o_out_fmap(xor_out[616*24*24*bW:617*24*24*bW-1]));
convchan2 c_2_617 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[617*5*5:618*5*5-1]), .o_out_fmap(xor_out[617*24*24*bW:618*24*24*bW-1]));
convchan2 c_2_618 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[618*5*5:619*5*5-1]), .o_out_fmap(xor_out[618*24*24*bW:619*24*24*bW-1]));
convchan2 c_2_619 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[619*5*5:620*5*5-1]), .o_out_fmap(xor_out[619*24*24*bW:620*24*24*bW-1]));
convchan2 c_2_620 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[620*5*5:621*5*5-1]), .o_out_fmap(xor_out[620*24*24*bW:621*24*24*bW-1]));
convchan2 c_2_621 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[621*5*5:622*5*5-1]), .o_out_fmap(xor_out[621*24*24*bW:622*24*24*bW-1]));
convchan2 c_2_622 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[622*5*5:623*5*5-1]), .o_out_fmap(xor_out[622*24*24*bW:623*24*24*bW-1]));
convchan2 c_2_623 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[623*5*5:624*5*5-1]), .o_out_fmap(xor_out[623*24*24*bW:624*24*24*bW-1]));
convchan2 c_2_624 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[624*5*5:625*5*5-1]), .o_out_fmap(xor_out[624*24*24*bW:625*24*24*bW-1]));
convchan2 c_2_625 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[625*5*5:626*5*5-1]), .o_out_fmap(xor_out[625*24*24*bW:626*24*24*bW-1]));
convchan2 c_2_626 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[626*5*5:627*5*5-1]), .o_out_fmap(xor_out[626*24*24*bW:627*24*24*bW-1]));
convchan2 c_2_627 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[627*5*5:628*5*5-1]), .o_out_fmap(xor_out[627*24*24*bW:628*24*24*bW-1]));
convchan2 c_2_628 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[628*5*5:629*5*5-1]), .o_out_fmap(xor_out[628*24*24*bW:629*24*24*bW-1]));
convchan2 c_2_629 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[629*5*5:630*5*5-1]), .o_out_fmap(xor_out[629*24*24*bW:630*24*24*bW-1]));
convchan2 c_2_630 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[630*5*5:631*5*5-1]), .o_out_fmap(xor_out[630*24*24*bW:631*24*24*bW-1]));
convchan2 c_2_631 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[631*5*5:632*5*5-1]), .o_out_fmap(xor_out[631*24*24*bW:632*24*24*bW-1]));
convchan2 c_2_632 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[632*5*5:633*5*5-1]), .o_out_fmap(xor_out[632*24*24*bW:633*24*24*bW-1]));
convchan2 c_2_633 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[633*5*5:634*5*5-1]), .o_out_fmap(xor_out[633*24*24*bW:634*24*24*bW-1]));
convchan2 c_2_634 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[634*5*5:635*5*5-1]), .o_out_fmap(xor_out[634*24*24*bW:635*24*24*bW-1]));
convchan2 c_2_635 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[635*5*5:636*5*5-1]), .o_out_fmap(xor_out[635*24*24*bW:636*24*24*bW-1]));
convchan2 c_2_636 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[636*5*5:637*5*5-1]), .o_out_fmap(xor_out[636*24*24*bW:637*24*24*bW-1]));
convchan2 c_2_637 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[637*5*5:638*5*5-1]), .o_out_fmap(xor_out[637*24*24*bW:638*24*24*bW-1]));
convchan2 c_2_638 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[638*5*5:639*5*5-1]), .o_out_fmap(xor_out[638*24*24*bW:639*24*24*bW-1]));
convchan2 c_2_639 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[639*5*5:640*5*5-1]), .o_out_fmap(xor_out[639*24*24*bW:640*24*24*bW-1]));
convchan2 c_2_640 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[640*5*5:641*5*5-1]), .o_out_fmap(xor_out[640*24*24*bW:641*24*24*bW-1]));
convchan2 c_2_641 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[641*5*5:642*5*5-1]), .o_out_fmap(xor_out[641*24*24*bW:642*24*24*bW-1]));
convchan2 c_2_642 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[642*5*5:643*5*5-1]), .o_out_fmap(xor_out[642*24*24*bW:643*24*24*bW-1]));
convchan2 c_2_643 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[643*5*5:644*5*5-1]), .o_out_fmap(xor_out[643*24*24*bW:644*24*24*bW-1]));
convchan2 c_2_644 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[644*5*5:645*5*5-1]), .o_out_fmap(xor_out[644*24*24*bW:645*24*24*bW-1]));
convchan2 c_2_645 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[645*5*5:646*5*5-1]), .o_out_fmap(xor_out[645*24*24*bW:646*24*24*bW-1]));
convchan2 c_2_646 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[646*5*5:647*5*5-1]), .o_out_fmap(xor_out[646*24*24*bW:647*24*24*bW-1]));
convchan2 c_2_647 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[647*5*5:648*5*5-1]), .o_out_fmap(xor_out[647*24*24*bW:648*24*24*bW-1]));
convchan2 c_2_648 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[648*5*5:649*5*5-1]), .o_out_fmap(xor_out[648*24*24*bW:649*24*24*bW-1]));
convchan2 c_2_649 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[649*5*5:650*5*5-1]), .o_out_fmap(xor_out[649*24*24*bW:650*24*24*bW-1]));
convchan2 c_2_650 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[650*5*5:651*5*5-1]), .o_out_fmap(xor_out[650*24*24*bW:651*24*24*bW-1]));
convchan2 c_2_651 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[651*5*5:652*5*5-1]), .o_out_fmap(xor_out[651*24*24*bW:652*24*24*bW-1]));
convchan2 c_2_652 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[652*5*5:653*5*5-1]), .o_out_fmap(xor_out[652*24*24*bW:653*24*24*bW-1]));
convchan2 c_2_653 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[653*5*5:654*5*5-1]), .o_out_fmap(xor_out[653*24*24*bW:654*24*24*bW-1]));
convchan2 c_2_654 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[654*5*5:655*5*5-1]), .o_out_fmap(xor_out[654*24*24*bW:655*24*24*bW-1]));
convchan2 c_2_655 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[655*5*5:656*5*5-1]), .o_out_fmap(xor_out[655*24*24*bW:656*24*24*bW-1]));
convchan2 c_2_656 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[656*5*5:657*5*5-1]), .o_out_fmap(xor_out[656*24*24*bW:657*24*24*bW-1]));
convchan2 c_2_657 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[657*5*5:658*5*5-1]), .o_out_fmap(xor_out[657*24*24*bW:658*24*24*bW-1]));
convchan2 c_2_658 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[658*5*5:659*5*5-1]), .o_out_fmap(xor_out[658*24*24*bW:659*24*24*bW-1]));
convchan2 c_2_659 (.i_image(image[10*12*12:11*12*12*+1]), .i_kernel(kernels[659*5*5:660*5*5-1]), .o_out_fmap(xor_out[659*24*24*bW:660*24*24*bW-1]));
convchan2 c_2_660 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[660*5*5:661*5*5-1]), .o_out_fmap(xor_out[660*24*24*bW:661*24*24*bW-1]));
convchan2 c_2_661 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[661*5*5:662*5*5-1]), .o_out_fmap(xor_out[661*24*24*bW:662*24*24*bW-1]));
convchan2 c_2_662 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[662*5*5:663*5*5-1]), .o_out_fmap(xor_out[662*24*24*bW:663*24*24*bW-1]));
convchan2 c_2_663 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[663*5*5:664*5*5-1]), .o_out_fmap(xor_out[663*24*24*bW:664*24*24*bW-1]));
convchan2 c_2_664 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[664*5*5:665*5*5-1]), .o_out_fmap(xor_out[664*24*24*bW:665*24*24*bW-1]));
convchan2 c_2_665 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[665*5*5:666*5*5-1]), .o_out_fmap(xor_out[665*24*24*bW:666*24*24*bW-1]));
convchan2 c_2_666 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[666*5*5:667*5*5-1]), .o_out_fmap(xor_out[666*24*24*bW:667*24*24*bW-1]));
convchan2 c_2_667 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[667*5*5:668*5*5-1]), .o_out_fmap(xor_out[667*24*24*bW:668*24*24*bW-1]));
convchan2 c_2_668 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[668*5*5:669*5*5-1]), .o_out_fmap(xor_out[668*24*24*bW:669*24*24*bW-1]));
convchan2 c_2_669 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[669*5*5:670*5*5-1]), .o_out_fmap(xor_out[669*24*24*bW:670*24*24*bW-1]));
convchan2 c_2_670 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[670*5*5:671*5*5-1]), .o_out_fmap(xor_out[670*24*24*bW:671*24*24*bW-1]));
convchan2 c_2_671 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[671*5*5:672*5*5-1]), .o_out_fmap(xor_out[671*24*24*bW:672*24*24*bW-1]));
convchan2 c_2_672 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[672*5*5:673*5*5-1]), .o_out_fmap(xor_out[672*24*24*bW:673*24*24*bW-1]));
convchan2 c_2_673 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[673*5*5:674*5*5-1]), .o_out_fmap(xor_out[673*24*24*bW:674*24*24*bW-1]));
convchan2 c_2_674 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[674*5*5:675*5*5-1]), .o_out_fmap(xor_out[674*24*24*bW:675*24*24*bW-1]));
convchan2 c_2_675 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[675*5*5:676*5*5-1]), .o_out_fmap(xor_out[675*24*24*bW:676*24*24*bW-1]));
convchan2 c_2_676 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[676*5*5:677*5*5-1]), .o_out_fmap(xor_out[676*24*24*bW:677*24*24*bW-1]));
convchan2 c_2_677 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[677*5*5:678*5*5-1]), .o_out_fmap(xor_out[677*24*24*bW:678*24*24*bW-1]));
convchan2 c_2_678 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[678*5*5:679*5*5-1]), .o_out_fmap(xor_out[678*24*24*bW:679*24*24*bW-1]));
convchan2 c_2_679 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[679*5*5:680*5*5-1]), .o_out_fmap(xor_out[679*24*24*bW:680*24*24*bW-1]));
convchan2 c_2_680 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[680*5*5:681*5*5-1]), .o_out_fmap(xor_out[680*24*24*bW:681*24*24*bW-1]));
convchan2 c_2_681 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[681*5*5:682*5*5-1]), .o_out_fmap(xor_out[681*24*24*bW:682*24*24*bW-1]));
convchan2 c_2_682 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[682*5*5:683*5*5-1]), .o_out_fmap(xor_out[682*24*24*bW:683*24*24*bW-1]));
convchan2 c_2_683 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[683*5*5:684*5*5-1]), .o_out_fmap(xor_out[683*24*24*bW:684*24*24*bW-1]));
convchan2 c_2_684 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[684*5*5:685*5*5-1]), .o_out_fmap(xor_out[684*24*24*bW:685*24*24*bW-1]));
convchan2 c_2_685 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[685*5*5:686*5*5-1]), .o_out_fmap(xor_out[685*24*24*bW:686*24*24*bW-1]));
convchan2 c_2_686 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[686*5*5:687*5*5-1]), .o_out_fmap(xor_out[686*24*24*bW:687*24*24*bW-1]));
convchan2 c_2_687 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[687*5*5:688*5*5-1]), .o_out_fmap(xor_out[687*24*24*bW:688*24*24*bW-1]));
convchan2 c_2_688 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[688*5*5:689*5*5-1]), .o_out_fmap(xor_out[688*24*24*bW:689*24*24*bW-1]));
convchan2 c_2_689 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[689*5*5:690*5*5-1]), .o_out_fmap(xor_out[689*24*24*bW:690*24*24*bW-1]));
convchan2 c_2_690 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[690*5*5:691*5*5-1]), .o_out_fmap(xor_out[690*24*24*bW:691*24*24*bW-1]));
convchan2 c_2_691 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[691*5*5:692*5*5-1]), .o_out_fmap(xor_out[691*24*24*bW:692*24*24*bW-1]));
convchan2 c_2_692 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[692*5*5:693*5*5-1]), .o_out_fmap(xor_out[692*24*24*bW:693*24*24*bW-1]));
convchan2 c_2_693 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[693*5*5:694*5*5-1]), .o_out_fmap(xor_out[693*24*24*bW:694*24*24*bW-1]));
convchan2 c_2_694 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[694*5*5:695*5*5-1]), .o_out_fmap(xor_out[694*24*24*bW:695*24*24*bW-1]));
convchan2 c_2_695 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[695*5*5:696*5*5-1]), .o_out_fmap(xor_out[695*24*24*bW:696*24*24*bW-1]));
convchan2 c_2_696 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[696*5*5:697*5*5-1]), .o_out_fmap(xor_out[696*24*24*bW:697*24*24*bW-1]));
convchan2 c_2_697 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[697*5*5:698*5*5-1]), .o_out_fmap(xor_out[697*24*24*bW:698*24*24*bW-1]));
convchan2 c_2_698 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[698*5*5:699*5*5-1]), .o_out_fmap(xor_out[698*24*24*bW:699*24*24*bW-1]));
convchan2 c_2_699 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[699*5*5:700*5*5-1]), .o_out_fmap(xor_out[699*24*24*bW:700*24*24*bW-1]));
convchan2 c_2_700 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[700*5*5:701*5*5-1]), .o_out_fmap(xor_out[700*24*24*bW:701*24*24*bW-1]));
convchan2 c_2_701 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[701*5*5:702*5*5-1]), .o_out_fmap(xor_out[701*24*24*bW:702*24*24*bW-1]));
convchan2 c_2_702 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[702*5*5:703*5*5-1]), .o_out_fmap(xor_out[702*24*24*bW:703*24*24*bW-1]));
convchan2 c_2_703 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[703*5*5:704*5*5-1]), .o_out_fmap(xor_out[703*24*24*bW:704*24*24*bW-1]));
convchan2 c_2_704 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[704*5*5:705*5*5-1]), .o_out_fmap(xor_out[704*24*24*bW:705*24*24*bW-1]));
convchan2 c_2_705 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[705*5*5:706*5*5-1]), .o_out_fmap(xor_out[705*24*24*bW:706*24*24*bW-1]));
convchan2 c_2_706 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[706*5*5:707*5*5-1]), .o_out_fmap(xor_out[706*24*24*bW:707*24*24*bW-1]));
convchan2 c_2_707 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[707*5*5:708*5*5-1]), .o_out_fmap(xor_out[707*24*24*bW:708*24*24*bW-1]));
convchan2 c_2_708 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[708*5*5:709*5*5-1]), .o_out_fmap(xor_out[708*24*24*bW:709*24*24*bW-1]));
convchan2 c_2_709 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[709*5*5:710*5*5-1]), .o_out_fmap(xor_out[709*24*24*bW:710*24*24*bW-1]));
convchan2 c_2_710 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[710*5*5:711*5*5-1]), .o_out_fmap(xor_out[710*24*24*bW:711*24*24*bW-1]));
convchan2 c_2_711 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[711*5*5:712*5*5-1]), .o_out_fmap(xor_out[711*24*24*bW:712*24*24*bW-1]));
convchan2 c_2_712 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[712*5*5:713*5*5-1]), .o_out_fmap(xor_out[712*24*24*bW:713*24*24*bW-1]));
convchan2 c_2_713 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[713*5*5:714*5*5-1]), .o_out_fmap(xor_out[713*24*24*bW:714*24*24*bW-1]));
convchan2 c_2_714 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[714*5*5:715*5*5-1]), .o_out_fmap(xor_out[714*24*24*bW:715*24*24*bW-1]));
convchan2 c_2_715 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[715*5*5:716*5*5-1]), .o_out_fmap(xor_out[715*24*24*bW:716*24*24*bW-1]));
convchan2 c_2_716 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[716*5*5:717*5*5-1]), .o_out_fmap(xor_out[716*24*24*bW:717*24*24*bW-1]));
convchan2 c_2_717 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[717*5*5:718*5*5-1]), .o_out_fmap(xor_out[717*24*24*bW:718*24*24*bW-1]));
convchan2 c_2_718 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[718*5*5:719*5*5-1]), .o_out_fmap(xor_out[718*24*24*bW:719*24*24*bW-1]));
convchan2 c_2_719 (.i_image(image[11*12*12:12*12*12*+1]), .i_kernel(kernels[719*5*5:720*5*5-1]), .o_out_fmap(xor_out[719*24*24*bW:720*24*24*bW-1]));
convchan2 c_2_720 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[720*5*5:721*5*5-1]), .o_out_fmap(xor_out[720*24*24*bW:721*24*24*bW-1]));
convchan2 c_2_721 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[721*5*5:722*5*5-1]), .o_out_fmap(xor_out[721*24*24*bW:722*24*24*bW-1]));
convchan2 c_2_722 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[722*5*5:723*5*5-1]), .o_out_fmap(xor_out[722*24*24*bW:723*24*24*bW-1]));
convchan2 c_2_723 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[723*5*5:724*5*5-1]), .o_out_fmap(xor_out[723*24*24*bW:724*24*24*bW-1]));
convchan2 c_2_724 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[724*5*5:725*5*5-1]), .o_out_fmap(xor_out[724*24*24*bW:725*24*24*bW-1]));
convchan2 c_2_725 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[725*5*5:726*5*5-1]), .o_out_fmap(xor_out[725*24*24*bW:726*24*24*bW-1]));
convchan2 c_2_726 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[726*5*5:727*5*5-1]), .o_out_fmap(xor_out[726*24*24*bW:727*24*24*bW-1]));
convchan2 c_2_727 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[727*5*5:728*5*5-1]), .o_out_fmap(xor_out[727*24*24*bW:728*24*24*bW-1]));
convchan2 c_2_728 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[728*5*5:729*5*5-1]), .o_out_fmap(xor_out[728*24*24*bW:729*24*24*bW-1]));
convchan2 c_2_729 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[729*5*5:730*5*5-1]), .o_out_fmap(xor_out[729*24*24*bW:730*24*24*bW-1]));
convchan2 c_2_730 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[730*5*5:731*5*5-1]), .o_out_fmap(xor_out[730*24*24*bW:731*24*24*bW-1]));
convchan2 c_2_731 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[731*5*5:732*5*5-1]), .o_out_fmap(xor_out[731*24*24*bW:732*24*24*bW-1]));
convchan2 c_2_732 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[732*5*5:733*5*5-1]), .o_out_fmap(xor_out[732*24*24*bW:733*24*24*bW-1]));
convchan2 c_2_733 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[733*5*5:734*5*5-1]), .o_out_fmap(xor_out[733*24*24*bW:734*24*24*bW-1]));
convchan2 c_2_734 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[734*5*5:735*5*5-1]), .o_out_fmap(xor_out[734*24*24*bW:735*24*24*bW-1]));
convchan2 c_2_735 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[735*5*5:736*5*5-1]), .o_out_fmap(xor_out[735*24*24*bW:736*24*24*bW-1]));
convchan2 c_2_736 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[736*5*5:737*5*5-1]), .o_out_fmap(xor_out[736*24*24*bW:737*24*24*bW-1]));
convchan2 c_2_737 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[737*5*5:738*5*5-1]), .o_out_fmap(xor_out[737*24*24*bW:738*24*24*bW-1]));
convchan2 c_2_738 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[738*5*5:739*5*5-1]), .o_out_fmap(xor_out[738*24*24*bW:739*24*24*bW-1]));
convchan2 c_2_739 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[739*5*5:740*5*5-1]), .o_out_fmap(xor_out[739*24*24*bW:740*24*24*bW-1]));
convchan2 c_2_740 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[740*5*5:741*5*5-1]), .o_out_fmap(xor_out[740*24*24*bW:741*24*24*bW-1]));
convchan2 c_2_741 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[741*5*5:742*5*5-1]), .o_out_fmap(xor_out[741*24*24*bW:742*24*24*bW-1]));
convchan2 c_2_742 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[742*5*5:743*5*5-1]), .o_out_fmap(xor_out[742*24*24*bW:743*24*24*bW-1]));
convchan2 c_2_743 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[743*5*5:744*5*5-1]), .o_out_fmap(xor_out[743*24*24*bW:744*24*24*bW-1]));
convchan2 c_2_744 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[744*5*5:745*5*5-1]), .o_out_fmap(xor_out[744*24*24*bW:745*24*24*bW-1]));
convchan2 c_2_745 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[745*5*5:746*5*5-1]), .o_out_fmap(xor_out[745*24*24*bW:746*24*24*bW-1]));
convchan2 c_2_746 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[746*5*5:747*5*5-1]), .o_out_fmap(xor_out[746*24*24*bW:747*24*24*bW-1]));
convchan2 c_2_747 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[747*5*5:748*5*5-1]), .o_out_fmap(xor_out[747*24*24*bW:748*24*24*bW-1]));
convchan2 c_2_748 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[748*5*5:749*5*5-1]), .o_out_fmap(xor_out[748*24*24*bW:749*24*24*bW-1]));
convchan2 c_2_749 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[749*5*5:750*5*5-1]), .o_out_fmap(xor_out[749*24*24*bW:750*24*24*bW-1]));
convchan2 c_2_750 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[750*5*5:751*5*5-1]), .o_out_fmap(xor_out[750*24*24*bW:751*24*24*bW-1]));
convchan2 c_2_751 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[751*5*5:752*5*5-1]), .o_out_fmap(xor_out[751*24*24*bW:752*24*24*bW-1]));
convchan2 c_2_752 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[752*5*5:753*5*5-1]), .o_out_fmap(xor_out[752*24*24*bW:753*24*24*bW-1]));
convchan2 c_2_753 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[753*5*5:754*5*5-1]), .o_out_fmap(xor_out[753*24*24*bW:754*24*24*bW-1]));
convchan2 c_2_754 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[754*5*5:755*5*5-1]), .o_out_fmap(xor_out[754*24*24*bW:755*24*24*bW-1]));
convchan2 c_2_755 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[755*5*5:756*5*5-1]), .o_out_fmap(xor_out[755*24*24*bW:756*24*24*bW-1]));
convchan2 c_2_756 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[756*5*5:757*5*5-1]), .o_out_fmap(xor_out[756*24*24*bW:757*24*24*bW-1]));
convchan2 c_2_757 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[757*5*5:758*5*5-1]), .o_out_fmap(xor_out[757*24*24*bW:758*24*24*bW-1]));
convchan2 c_2_758 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[758*5*5:759*5*5-1]), .o_out_fmap(xor_out[758*24*24*bW:759*24*24*bW-1]));
convchan2 c_2_759 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[759*5*5:760*5*5-1]), .o_out_fmap(xor_out[759*24*24*bW:760*24*24*bW-1]));
convchan2 c_2_760 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[760*5*5:761*5*5-1]), .o_out_fmap(xor_out[760*24*24*bW:761*24*24*bW-1]));
convchan2 c_2_761 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[761*5*5:762*5*5-1]), .o_out_fmap(xor_out[761*24*24*bW:762*24*24*bW-1]));
convchan2 c_2_762 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[762*5*5:763*5*5-1]), .o_out_fmap(xor_out[762*24*24*bW:763*24*24*bW-1]));
convchan2 c_2_763 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[763*5*5:764*5*5-1]), .o_out_fmap(xor_out[763*24*24*bW:764*24*24*bW-1]));
convchan2 c_2_764 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[764*5*5:765*5*5-1]), .o_out_fmap(xor_out[764*24*24*bW:765*24*24*bW-1]));
convchan2 c_2_765 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[765*5*5:766*5*5-1]), .o_out_fmap(xor_out[765*24*24*bW:766*24*24*bW-1]));
convchan2 c_2_766 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[766*5*5:767*5*5-1]), .o_out_fmap(xor_out[766*24*24*bW:767*24*24*bW-1]));
convchan2 c_2_767 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[767*5*5:768*5*5-1]), .o_out_fmap(xor_out[767*24*24*bW:768*24*24*bW-1]));
convchan2 c_2_768 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[768*5*5:769*5*5-1]), .o_out_fmap(xor_out[768*24*24*bW:769*24*24*bW-1]));
convchan2 c_2_769 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[769*5*5:770*5*5-1]), .o_out_fmap(xor_out[769*24*24*bW:770*24*24*bW-1]));
convchan2 c_2_770 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[770*5*5:771*5*5-1]), .o_out_fmap(xor_out[770*24*24*bW:771*24*24*bW-1]));
convchan2 c_2_771 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[771*5*5:772*5*5-1]), .o_out_fmap(xor_out[771*24*24*bW:772*24*24*bW-1]));
convchan2 c_2_772 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[772*5*5:773*5*5-1]), .o_out_fmap(xor_out[772*24*24*bW:773*24*24*bW-1]));
convchan2 c_2_773 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[773*5*5:774*5*5-1]), .o_out_fmap(xor_out[773*24*24*bW:774*24*24*bW-1]));
convchan2 c_2_774 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[774*5*5:775*5*5-1]), .o_out_fmap(xor_out[774*24*24*bW:775*24*24*bW-1]));
convchan2 c_2_775 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[775*5*5:776*5*5-1]), .o_out_fmap(xor_out[775*24*24*bW:776*24*24*bW-1]));
convchan2 c_2_776 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[776*5*5:777*5*5-1]), .o_out_fmap(xor_out[776*24*24*bW:777*24*24*bW-1]));
convchan2 c_2_777 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[777*5*5:778*5*5-1]), .o_out_fmap(xor_out[777*24*24*bW:778*24*24*bW-1]));
convchan2 c_2_778 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[778*5*5:779*5*5-1]), .o_out_fmap(xor_out[778*24*24*bW:779*24*24*bW-1]));
convchan2 c_2_779 (.i_image(image[12*12*12:13*12*12*+1]), .i_kernel(kernels[779*5*5:780*5*5-1]), .o_out_fmap(xor_out[779*24*24*bW:780*24*24*bW-1]));
convchan2 c_2_780 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[780*5*5:781*5*5-1]), .o_out_fmap(xor_out[780*24*24*bW:781*24*24*bW-1]));
convchan2 c_2_781 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[781*5*5:782*5*5-1]), .o_out_fmap(xor_out[781*24*24*bW:782*24*24*bW-1]));
convchan2 c_2_782 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[782*5*5:783*5*5-1]), .o_out_fmap(xor_out[782*24*24*bW:783*24*24*bW-1]));
convchan2 c_2_783 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[783*5*5:784*5*5-1]), .o_out_fmap(xor_out[783*24*24*bW:784*24*24*bW-1]));
convchan2 c_2_784 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[784*5*5:785*5*5-1]), .o_out_fmap(xor_out[784*24*24*bW:785*24*24*bW-1]));
convchan2 c_2_785 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[785*5*5:786*5*5-1]), .o_out_fmap(xor_out[785*24*24*bW:786*24*24*bW-1]));
convchan2 c_2_786 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[786*5*5:787*5*5-1]), .o_out_fmap(xor_out[786*24*24*bW:787*24*24*bW-1]));
convchan2 c_2_787 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[787*5*5:788*5*5-1]), .o_out_fmap(xor_out[787*24*24*bW:788*24*24*bW-1]));
convchan2 c_2_788 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[788*5*5:789*5*5-1]), .o_out_fmap(xor_out[788*24*24*bW:789*24*24*bW-1]));
convchan2 c_2_789 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[789*5*5:790*5*5-1]), .o_out_fmap(xor_out[789*24*24*bW:790*24*24*bW-1]));
convchan2 c_2_790 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[790*5*5:791*5*5-1]), .o_out_fmap(xor_out[790*24*24*bW:791*24*24*bW-1]));
convchan2 c_2_791 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[791*5*5:792*5*5-1]), .o_out_fmap(xor_out[791*24*24*bW:792*24*24*bW-1]));
convchan2 c_2_792 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[792*5*5:793*5*5-1]), .o_out_fmap(xor_out[792*24*24*bW:793*24*24*bW-1]));
convchan2 c_2_793 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[793*5*5:794*5*5-1]), .o_out_fmap(xor_out[793*24*24*bW:794*24*24*bW-1]));
convchan2 c_2_794 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[794*5*5:795*5*5-1]), .o_out_fmap(xor_out[794*24*24*bW:795*24*24*bW-1]));
convchan2 c_2_795 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[795*5*5:796*5*5-1]), .o_out_fmap(xor_out[795*24*24*bW:796*24*24*bW-1]));
convchan2 c_2_796 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[796*5*5:797*5*5-1]), .o_out_fmap(xor_out[796*24*24*bW:797*24*24*bW-1]));
convchan2 c_2_797 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[797*5*5:798*5*5-1]), .o_out_fmap(xor_out[797*24*24*bW:798*24*24*bW-1]));
convchan2 c_2_798 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[798*5*5:799*5*5-1]), .o_out_fmap(xor_out[798*24*24*bW:799*24*24*bW-1]));
convchan2 c_2_799 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[799*5*5:800*5*5-1]), .o_out_fmap(xor_out[799*24*24*bW:800*24*24*bW-1]));
convchan2 c_2_800 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[800*5*5:801*5*5-1]), .o_out_fmap(xor_out[800*24*24*bW:801*24*24*bW-1]));
convchan2 c_2_801 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[801*5*5:802*5*5-1]), .o_out_fmap(xor_out[801*24*24*bW:802*24*24*bW-1]));
convchan2 c_2_802 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[802*5*5:803*5*5-1]), .o_out_fmap(xor_out[802*24*24*bW:803*24*24*bW-1]));
convchan2 c_2_803 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[803*5*5:804*5*5-1]), .o_out_fmap(xor_out[803*24*24*bW:804*24*24*bW-1]));
convchan2 c_2_804 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[804*5*5:805*5*5-1]), .o_out_fmap(xor_out[804*24*24*bW:805*24*24*bW-1]));
convchan2 c_2_805 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[805*5*5:806*5*5-1]), .o_out_fmap(xor_out[805*24*24*bW:806*24*24*bW-1]));
convchan2 c_2_806 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[806*5*5:807*5*5-1]), .o_out_fmap(xor_out[806*24*24*bW:807*24*24*bW-1]));
convchan2 c_2_807 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[807*5*5:808*5*5-1]), .o_out_fmap(xor_out[807*24*24*bW:808*24*24*bW-1]));
convchan2 c_2_808 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[808*5*5:809*5*5-1]), .o_out_fmap(xor_out[808*24*24*bW:809*24*24*bW-1]));
convchan2 c_2_809 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[809*5*5:810*5*5-1]), .o_out_fmap(xor_out[809*24*24*bW:810*24*24*bW-1]));
convchan2 c_2_810 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[810*5*5:811*5*5-1]), .o_out_fmap(xor_out[810*24*24*bW:811*24*24*bW-1]));
convchan2 c_2_811 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[811*5*5:812*5*5-1]), .o_out_fmap(xor_out[811*24*24*bW:812*24*24*bW-1]));
convchan2 c_2_812 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[812*5*5:813*5*5-1]), .o_out_fmap(xor_out[812*24*24*bW:813*24*24*bW-1]));
convchan2 c_2_813 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[813*5*5:814*5*5-1]), .o_out_fmap(xor_out[813*24*24*bW:814*24*24*bW-1]));
convchan2 c_2_814 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[814*5*5:815*5*5-1]), .o_out_fmap(xor_out[814*24*24*bW:815*24*24*bW-1]));
convchan2 c_2_815 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[815*5*5:816*5*5-1]), .o_out_fmap(xor_out[815*24*24*bW:816*24*24*bW-1]));
convchan2 c_2_816 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[816*5*5:817*5*5-1]), .o_out_fmap(xor_out[816*24*24*bW:817*24*24*bW-1]));
convchan2 c_2_817 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[817*5*5:818*5*5-1]), .o_out_fmap(xor_out[817*24*24*bW:818*24*24*bW-1]));
convchan2 c_2_818 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[818*5*5:819*5*5-1]), .o_out_fmap(xor_out[818*24*24*bW:819*24*24*bW-1]));
convchan2 c_2_819 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[819*5*5:820*5*5-1]), .o_out_fmap(xor_out[819*24*24*bW:820*24*24*bW-1]));
convchan2 c_2_820 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[820*5*5:821*5*5-1]), .o_out_fmap(xor_out[820*24*24*bW:821*24*24*bW-1]));
convchan2 c_2_821 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[821*5*5:822*5*5-1]), .o_out_fmap(xor_out[821*24*24*bW:822*24*24*bW-1]));
convchan2 c_2_822 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[822*5*5:823*5*5-1]), .o_out_fmap(xor_out[822*24*24*bW:823*24*24*bW-1]));
convchan2 c_2_823 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[823*5*5:824*5*5-1]), .o_out_fmap(xor_out[823*24*24*bW:824*24*24*bW-1]));
convchan2 c_2_824 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[824*5*5:825*5*5-1]), .o_out_fmap(xor_out[824*24*24*bW:825*24*24*bW-1]));
convchan2 c_2_825 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[825*5*5:826*5*5-1]), .o_out_fmap(xor_out[825*24*24*bW:826*24*24*bW-1]));
convchan2 c_2_826 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[826*5*5:827*5*5-1]), .o_out_fmap(xor_out[826*24*24*bW:827*24*24*bW-1]));
convchan2 c_2_827 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[827*5*5:828*5*5-1]), .o_out_fmap(xor_out[827*24*24*bW:828*24*24*bW-1]));
convchan2 c_2_828 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[828*5*5:829*5*5-1]), .o_out_fmap(xor_out[828*24*24*bW:829*24*24*bW-1]));
convchan2 c_2_829 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[829*5*5:830*5*5-1]), .o_out_fmap(xor_out[829*24*24*bW:830*24*24*bW-1]));
convchan2 c_2_830 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[830*5*5:831*5*5-1]), .o_out_fmap(xor_out[830*24*24*bW:831*24*24*bW-1]));
convchan2 c_2_831 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[831*5*5:832*5*5-1]), .o_out_fmap(xor_out[831*24*24*bW:832*24*24*bW-1]));
convchan2 c_2_832 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[832*5*5:833*5*5-1]), .o_out_fmap(xor_out[832*24*24*bW:833*24*24*bW-1]));
convchan2 c_2_833 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[833*5*5:834*5*5-1]), .o_out_fmap(xor_out[833*24*24*bW:834*24*24*bW-1]));
convchan2 c_2_834 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[834*5*5:835*5*5-1]), .o_out_fmap(xor_out[834*24*24*bW:835*24*24*bW-1]));
convchan2 c_2_835 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[835*5*5:836*5*5-1]), .o_out_fmap(xor_out[835*24*24*bW:836*24*24*bW-1]));
convchan2 c_2_836 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[836*5*5:837*5*5-1]), .o_out_fmap(xor_out[836*24*24*bW:837*24*24*bW-1]));
convchan2 c_2_837 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[837*5*5:838*5*5-1]), .o_out_fmap(xor_out[837*24*24*bW:838*24*24*bW-1]));
convchan2 c_2_838 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[838*5*5:839*5*5-1]), .o_out_fmap(xor_out[838*24*24*bW:839*24*24*bW-1]));
convchan2 c_2_839 (.i_image(image[13*12*12:14*12*12*+1]), .i_kernel(kernels[839*5*5:840*5*5-1]), .o_out_fmap(xor_out[839*24*24*bW:840*24*24*bW-1]));
convchan2 c_2_840 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[840*5*5:841*5*5-1]), .o_out_fmap(xor_out[840*24*24*bW:841*24*24*bW-1]));
convchan2 c_2_841 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[841*5*5:842*5*5-1]), .o_out_fmap(xor_out[841*24*24*bW:842*24*24*bW-1]));
convchan2 c_2_842 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[842*5*5:843*5*5-1]), .o_out_fmap(xor_out[842*24*24*bW:843*24*24*bW-1]));
convchan2 c_2_843 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[843*5*5:844*5*5-1]), .o_out_fmap(xor_out[843*24*24*bW:844*24*24*bW-1]));
convchan2 c_2_844 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[844*5*5:845*5*5-1]), .o_out_fmap(xor_out[844*24*24*bW:845*24*24*bW-1]));
convchan2 c_2_845 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[845*5*5:846*5*5-1]), .o_out_fmap(xor_out[845*24*24*bW:846*24*24*bW-1]));
convchan2 c_2_846 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[846*5*5:847*5*5-1]), .o_out_fmap(xor_out[846*24*24*bW:847*24*24*bW-1]));
convchan2 c_2_847 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[847*5*5:848*5*5-1]), .o_out_fmap(xor_out[847*24*24*bW:848*24*24*bW-1]));
convchan2 c_2_848 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[848*5*5:849*5*5-1]), .o_out_fmap(xor_out[848*24*24*bW:849*24*24*bW-1]));
convchan2 c_2_849 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[849*5*5:850*5*5-1]), .o_out_fmap(xor_out[849*24*24*bW:850*24*24*bW-1]));
convchan2 c_2_850 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[850*5*5:851*5*5-1]), .o_out_fmap(xor_out[850*24*24*bW:851*24*24*bW-1]));
convchan2 c_2_851 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[851*5*5:852*5*5-1]), .o_out_fmap(xor_out[851*24*24*bW:852*24*24*bW-1]));
convchan2 c_2_852 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[852*5*5:853*5*5-1]), .o_out_fmap(xor_out[852*24*24*bW:853*24*24*bW-1]));
convchan2 c_2_853 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[853*5*5:854*5*5-1]), .o_out_fmap(xor_out[853*24*24*bW:854*24*24*bW-1]));
convchan2 c_2_854 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[854*5*5:855*5*5-1]), .o_out_fmap(xor_out[854*24*24*bW:855*24*24*bW-1]));
convchan2 c_2_855 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[855*5*5:856*5*5-1]), .o_out_fmap(xor_out[855*24*24*bW:856*24*24*bW-1]));
convchan2 c_2_856 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[856*5*5:857*5*5-1]), .o_out_fmap(xor_out[856*24*24*bW:857*24*24*bW-1]));
convchan2 c_2_857 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[857*5*5:858*5*5-1]), .o_out_fmap(xor_out[857*24*24*bW:858*24*24*bW-1]));
convchan2 c_2_858 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[858*5*5:859*5*5-1]), .o_out_fmap(xor_out[858*24*24*bW:859*24*24*bW-1]));
convchan2 c_2_859 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[859*5*5:860*5*5-1]), .o_out_fmap(xor_out[859*24*24*bW:860*24*24*bW-1]));
convchan2 c_2_860 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[860*5*5:861*5*5-1]), .o_out_fmap(xor_out[860*24*24*bW:861*24*24*bW-1]));
convchan2 c_2_861 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[861*5*5:862*5*5-1]), .o_out_fmap(xor_out[861*24*24*bW:862*24*24*bW-1]));
convchan2 c_2_862 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[862*5*5:863*5*5-1]), .o_out_fmap(xor_out[862*24*24*bW:863*24*24*bW-1]));
convchan2 c_2_863 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[863*5*5:864*5*5-1]), .o_out_fmap(xor_out[863*24*24*bW:864*24*24*bW-1]));
convchan2 c_2_864 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[864*5*5:865*5*5-1]), .o_out_fmap(xor_out[864*24*24*bW:865*24*24*bW-1]));
convchan2 c_2_865 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[865*5*5:866*5*5-1]), .o_out_fmap(xor_out[865*24*24*bW:866*24*24*bW-1]));
convchan2 c_2_866 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[866*5*5:867*5*5-1]), .o_out_fmap(xor_out[866*24*24*bW:867*24*24*bW-1]));
convchan2 c_2_867 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[867*5*5:868*5*5-1]), .o_out_fmap(xor_out[867*24*24*bW:868*24*24*bW-1]));
convchan2 c_2_868 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[868*5*5:869*5*5-1]), .o_out_fmap(xor_out[868*24*24*bW:869*24*24*bW-1]));
convchan2 c_2_869 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[869*5*5:870*5*5-1]), .o_out_fmap(xor_out[869*24*24*bW:870*24*24*bW-1]));
convchan2 c_2_870 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[870*5*5:871*5*5-1]), .o_out_fmap(xor_out[870*24*24*bW:871*24*24*bW-1]));
convchan2 c_2_871 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[871*5*5:872*5*5-1]), .o_out_fmap(xor_out[871*24*24*bW:872*24*24*bW-1]));
convchan2 c_2_872 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[872*5*5:873*5*5-1]), .o_out_fmap(xor_out[872*24*24*bW:873*24*24*bW-1]));
convchan2 c_2_873 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[873*5*5:874*5*5-1]), .o_out_fmap(xor_out[873*24*24*bW:874*24*24*bW-1]));
convchan2 c_2_874 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[874*5*5:875*5*5-1]), .o_out_fmap(xor_out[874*24*24*bW:875*24*24*bW-1]));
convchan2 c_2_875 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[875*5*5:876*5*5-1]), .o_out_fmap(xor_out[875*24*24*bW:876*24*24*bW-1]));
convchan2 c_2_876 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[876*5*5:877*5*5-1]), .o_out_fmap(xor_out[876*24*24*bW:877*24*24*bW-1]));
convchan2 c_2_877 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[877*5*5:878*5*5-1]), .o_out_fmap(xor_out[877*24*24*bW:878*24*24*bW-1]));
convchan2 c_2_878 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[878*5*5:879*5*5-1]), .o_out_fmap(xor_out[878*24*24*bW:879*24*24*bW-1]));
convchan2 c_2_879 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[879*5*5:880*5*5-1]), .o_out_fmap(xor_out[879*24*24*bW:880*24*24*bW-1]));
convchan2 c_2_880 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[880*5*5:881*5*5-1]), .o_out_fmap(xor_out[880*24*24*bW:881*24*24*bW-1]));
convchan2 c_2_881 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[881*5*5:882*5*5-1]), .o_out_fmap(xor_out[881*24*24*bW:882*24*24*bW-1]));
convchan2 c_2_882 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[882*5*5:883*5*5-1]), .o_out_fmap(xor_out[882*24*24*bW:883*24*24*bW-1]));
convchan2 c_2_883 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[883*5*5:884*5*5-1]), .o_out_fmap(xor_out[883*24*24*bW:884*24*24*bW-1]));
convchan2 c_2_884 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[884*5*5:885*5*5-1]), .o_out_fmap(xor_out[884*24*24*bW:885*24*24*bW-1]));
convchan2 c_2_885 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[885*5*5:886*5*5-1]), .o_out_fmap(xor_out[885*24*24*bW:886*24*24*bW-1]));
convchan2 c_2_886 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[886*5*5:887*5*5-1]), .o_out_fmap(xor_out[886*24*24*bW:887*24*24*bW-1]));
convchan2 c_2_887 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[887*5*5:888*5*5-1]), .o_out_fmap(xor_out[887*24*24*bW:888*24*24*bW-1]));
convchan2 c_2_888 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[888*5*5:889*5*5-1]), .o_out_fmap(xor_out[888*24*24*bW:889*24*24*bW-1]));
convchan2 c_2_889 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[889*5*5:890*5*5-1]), .o_out_fmap(xor_out[889*24*24*bW:890*24*24*bW-1]));
convchan2 c_2_890 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[890*5*5:891*5*5-1]), .o_out_fmap(xor_out[890*24*24*bW:891*24*24*bW-1]));
convchan2 c_2_891 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[891*5*5:892*5*5-1]), .o_out_fmap(xor_out[891*24*24*bW:892*24*24*bW-1]));
convchan2 c_2_892 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[892*5*5:893*5*5-1]), .o_out_fmap(xor_out[892*24*24*bW:893*24*24*bW-1]));
convchan2 c_2_893 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[893*5*5:894*5*5-1]), .o_out_fmap(xor_out[893*24*24*bW:894*24*24*bW-1]));
convchan2 c_2_894 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[894*5*5:895*5*5-1]), .o_out_fmap(xor_out[894*24*24*bW:895*24*24*bW-1]));
convchan2 c_2_895 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[895*5*5:896*5*5-1]), .o_out_fmap(xor_out[895*24*24*bW:896*24*24*bW-1]));
convchan2 c_2_896 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[896*5*5:897*5*5-1]), .o_out_fmap(xor_out[896*24*24*bW:897*24*24*bW-1]));
convchan2 c_2_897 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[897*5*5:898*5*5-1]), .o_out_fmap(xor_out[897*24*24*bW:898*24*24*bW-1]));
convchan2 c_2_898 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[898*5*5:899*5*5-1]), .o_out_fmap(xor_out[898*24*24*bW:899*24*24*bW-1]));
convchan2 c_2_899 (.i_image(image[14*12*12:15*12*12*+1]), .i_kernel(kernels[899*5*5:900*5*5-1]), .o_out_fmap(xor_out[899*24*24*bW:900*24*24*bW-1]));
convchan2 c_2_900 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[900*5*5:901*5*5-1]), .o_out_fmap(xor_out[900*24*24*bW:901*24*24*bW-1]));
convchan2 c_2_901 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[901*5*5:902*5*5-1]), .o_out_fmap(xor_out[901*24*24*bW:902*24*24*bW-1]));
convchan2 c_2_902 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[902*5*5:903*5*5-1]), .o_out_fmap(xor_out[902*24*24*bW:903*24*24*bW-1]));
convchan2 c_2_903 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[903*5*5:904*5*5-1]), .o_out_fmap(xor_out[903*24*24*bW:904*24*24*bW-1]));
convchan2 c_2_904 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[904*5*5:905*5*5-1]), .o_out_fmap(xor_out[904*24*24*bW:905*24*24*bW-1]));
convchan2 c_2_905 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[905*5*5:906*5*5-1]), .o_out_fmap(xor_out[905*24*24*bW:906*24*24*bW-1]));
convchan2 c_2_906 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[906*5*5:907*5*5-1]), .o_out_fmap(xor_out[906*24*24*bW:907*24*24*bW-1]));
convchan2 c_2_907 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[907*5*5:908*5*5-1]), .o_out_fmap(xor_out[907*24*24*bW:908*24*24*bW-1]));
convchan2 c_2_908 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[908*5*5:909*5*5-1]), .o_out_fmap(xor_out[908*24*24*bW:909*24*24*bW-1]));
convchan2 c_2_909 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[909*5*5:910*5*5-1]), .o_out_fmap(xor_out[909*24*24*bW:910*24*24*bW-1]));
convchan2 c_2_910 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[910*5*5:911*5*5-1]), .o_out_fmap(xor_out[910*24*24*bW:911*24*24*bW-1]));
convchan2 c_2_911 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[911*5*5:912*5*5-1]), .o_out_fmap(xor_out[911*24*24*bW:912*24*24*bW-1]));
convchan2 c_2_912 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[912*5*5:913*5*5-1]), .o_out_fmap(xor_out[912*24*24*bW:913*24*24*bW-1]));
convchan2 c_2_913 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[913*5*5:914*5*5-1]), .o_out_fmap(xor_out[913*24*24*bW:914*24*24*bW-1]));
convchan2 c_2_914 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[914*5*5:915*5*5-1]), .o_out_fmap(xor_out[914*24*24*bW:915*24*24*bW-1]));
convchan2 c_2_915 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[915*5*5:916*5*5-1]), .o_out_fmap(xor_out[915*24*24*bW:916*24*24*bW-1]));
convchan2 c_2_916 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[916*5*5:917*5*5-1]), .o_out_fmap(xor_out[916*24*24*bW:917*24*24*bW-1]));
convchan2 c_2_917 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[917*5*5:918*5*5-1]), .o_out_fmap(xor_out[917*24*24*bW:918*24*24*bW-1]));
convchan2 c_2_918 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[918*5*5:919*5*5-1]), .o_out_fmap(xor_out[918*24*24*bW:919*24*24*bW-1]));
convchan2 c_2_919 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[919*5*5:920*5*5-1]), .o_out_fmap(xor_out[919*24*24*bW:920*24*24*bW-1]));
convchan2 c_2_920 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[920*5*5:921*5*5-1]), .o_out_fmap(xor_out[920*24*24*bW:921*24*24*bW-1]));
convchan2 c_2_921 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[921*5*5:922*5*5-1]), .o_out_fmap(xor_out[921*24*24*bW:922*24*24*bW-1]));
convchan2 c_2_922 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[922*5*5:923*5*5-1]), .o_out_fmap(xor_out[922*24*24*bW:923*24*24*bW-1]));
convchan2 c_2_923 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[923*5*5:924*5*5-1]), .o_out_fmap(xor_out[923*24*24*bW:924*24*24*bW-1]));
convchan2 c_2_924 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[924*5*5:925*5*5-1]), .o_out_fmap(xor_out[924*24*24*bW:925*24*24*bW-1]));
convchan2 c_2_925 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[925*5*5:926*5*5-1]), .o_out_fmap(xor_out[925*24*24*bW:926*24*24*bW-1]));
convchan2 c_2_926 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[926*5*5:927*5*5-1]), .o_out_fmap(xor_out[926*24*24*bW:927*24*24*bW-1]));
convchan2 c_2_927 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[927*5*5:928*5*5-1]), .o_out_fmap(xor_out[927*24*24*bW:928*24*24*bW-1]));
convchan2 c_2_928 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[928*5*5:929*5*5-1]), .o_out_fmap(xor_out[928*24*24*bW:929*24*24*bW-1]));
convchan2 c_2_929 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[929*5*5:930*5*5-1]), .o_out_fmap(xor_out[929*24*24*bW:930*24*24*bW-1]));
convchan2 c_2_930 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[930*5*5:931*5*5-1]), .o_out_fmap(xor_out[930*24*24*bW:931*24*24*bW-1]));
convchan2 c_2_931 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[931*5*5:932*5*5-1]), .o_out_fmap(xor_out[931*24*24*bW:932*24*24*bW-1]));
convchan2 c_2_932 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[932*5*5:933*5*5-1]), .o_out_fmap(xor_out[932*24*24*bW:933*24*24*bW-1]));
convchan2 c_2_933 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[933*5*5:934*5*5-1]), .o_out_fmap(xor_out[933*24*24*bW:934*24*24*bW-1]));
convchan2 c_2_934 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[934*5*5:935*5*5-1]), .o_out_fmap(xor_out[934*24*24*bW:935*24*24*bW-1]));
convchan2 c_2_935 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[935*5*5:936*5*5-1]), .o_out_fmap(xor_out[935*24*24*bW:936*24*24*bW-1]));
convchan2 c_2_936 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[936*5*5:937*5*5-1]), .o_out_fmap(xor_out[936*24*24*bW:937*24*24*bW-1]));
convchan2 c_2_937 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[937*5*5:938*5*5-1]), .o_out_fmap(xor_out[937*24*24*bW:938*24*24*bW-1]));
convchan2 c_2_938 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[938*5*5:939*5*5-1]), .o_out_fmap(xor_out[938*24*24*bW:939*24*24*bW-1]));
convchan2 c_2_939 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[939*5*5:940*5*5-1]), .o_out_fmap(xor_out[939*24*24*bW:940*24*24*bW-1]));
convchan2 c_2_940 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[940*5*5:941*5*5-1]), .o_out_fmap(xor_out[940*24*24*bW:941*24*24*bW-1]));
convchan2 c_2_941 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[941*5*5:942*5*5-1]), .o_out_fmap(xor_out[941*24*24*bW:942*24*24*bW-1]));
convchan2 c_2_942 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[942*5*5:943*5*5-1]), .o_out_fmap(xor_out[942*24*24*bW:943*24*24*bW-1]));
convchan2 c_2_943 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[943*5*5:944*5*5-1]), .o_out_fmap(xor_out[943*24*24*bW:944*24*24*bW-1]));
convchan2 c_2_944 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[944*5*5:945*5*5-1]), .o_out_fmap(xor_out[944*24*24*bW:945*24*24*bW-1]));
convchan2 c_2_945 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[945*5*5:946*5*5-1]), .o_out_fmap(xor_out[945*24*24*bW:946*24*24*bW-1]));
convchan2 c_2_946 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[946*5*5:947*5*5-1]), .o_out_fmap(xor_out[946*24*24*bW:947*24*24*bW-1]));
convchan2 c_2_947 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[947*5*5:948*5*5-1]), .o_out_fmap(xor_out[947*24*24*bW:948*24*24*bW-1]));
convchan2 c_2_948 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[948*5*5:949*5*5-1]), .o_out_fmap(xor_out[948*24*24*bW:949*24*24*bW-1]));
convchan2 c_2_949 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[949*5*5:950*5*5-1]), .o_out_fmap(xor_out[949*24*24*bW:950*24*24*bW-1]));
convchan2 c_2_950 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[950*5*5:951*5*5-1]), .o_out_fmap(xor_out[950*24*24*bW:951*24*24*bW-1]));
convchan2 c_2_951 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[951*5*5:952*5*5-1]), .o_out_fmap(xor_out[951*24*24*bW:952*24*24*bW-1]));
convchan2 c_2_952 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[952*5*5:953*5*5-1]), .o_out_fmap(xor_out[952*24*24*bW:953*24*24*bW-1]));
convchan2 c_2_953 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[953*5*5:954*5*5-1]), .o_out_fmap(xor_out[953*24*24*bW:954*24*24*bW-1]));
convchan2 c_2_954 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[954*5*5:955*5*5-1]), .o_out_fmap(xor_out[954*24*24*bW:955*24*24*bW-1]));
convchan2 c_2_955 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[955*5*5:956*5*5-1]), .o_out_fmap(xor_out[955*24*24*bW:956*24*24*bW-1]));
convchan2 c_2_956 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[956*5*5:957*5*5-1]), .o_out_fmap(xor_out[956*24*24*bW:957*24*24*bW-1]));
convchan2 c_2_957 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[957*5*5:958*5*5-1]), .o_out_fmap(xor_out[957*24*24*bW:958*24*24*bW-1]));
convchan2 c_2_958 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[958*5*5:959*5*5-1]), .o_out_fmap(xor_out[958*24*24*bW:959*24*24*bW-1]));
convchan2 c_2_959 (.i_image(image[15*12*12:16*12*12*+1]), .i_kernel(kernels[959*5*5:960*5*5-1]), .o_out_fmap(xor_out[959*24*24*bW:960*24*24*bW-1]));
convchan2 c_2_960 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[960*5*5:961*5*5-1]), .o_out_fmap(xor_out[960*24*24*bW:961*24*24*bW-1]));
convchan2 c_2_961 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[961*5*5:962*5*5-1]), .o_out_fmap(xor_out[961*24*24*bW:962*24*24*bW-1]));
convchan2 c_2_962 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[962*5*5:963*5*5-1]), .o_out_fmap(xor_out[962*24*24*bW:963*24*24*bW-1]));
convchan2 c_2_963 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[963*5*5:964*5*5-1]), .o_out_fmap(xor_out[963*24*24*bW:964*24*24*bW-1]));
convchan2 c_2_964 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[964*5*5:965*5*5-1]), .o_out_fmap(xor_out[964*24*24*bW:965*24*24*bW-1]));
convchan2 c_2_965 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[965*5*5:966*5*5-1]), .o_out_fmap(xor_out[965*24*24*bW:966*24*24*bW-1]));
convchan2 c_2_966 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[966*5*5:967*5*5-1]), .o_out_fmap(xor_out[966*24*24*bW:967*24*24*bW-1]));
convchan2 c_2_967 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[967*5*5:968*5*5-1]), .o_out_fmap(xor_out[967*24*24*bW:968*24*24*bW-1]));
convchan2 c_2_968 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[968*5*5:969*5*5-1]), .o_out_fmap(xor_out[968*24*24*bW:969*24*24*bW-1]));
convchan2 c_2_969 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[969*5*5:970*5*5-1]), .o_out_fmap(xor_out[969*24*24*bW:970*24*24*bW-1]));
convchan2 c_2_970 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[970*5*5:971*5*5-1]), .o_out_fmap(xor_out[970*24*24*bW:971*24*24*bW-1]));
convchan2 c_2_971 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[971*5*5:972*5*5-1]), .o_out_fmap(xor_out[971*24*24*bW:972*24*24*bW-1]));
convchan2 c_2_972 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[972*5*5:973*5*5-1]), .o_out_fmap(xor_out[972*24*24*bW:973*24*24*bW-1]));
convchan2 c_2_973 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[973*5*5:974*5*5-1]), .o_out_fmap(xor_out[973*24*24*bW:974*24*24*bW-1]));
convchan2 c_2_974 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[974*5*5:975*5*5-1]), .o_out_fmap(xor_out[974*24*24*bW:975*24*24*bW-1]));
convchan2 c_2_975 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[975*5*5:976*5*5-1]), .o_out_fmap(xor_out[975*24*24*bW:976*24*24*bW-1]));
convchan2 c_2_976 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[976*5*5:977*5*5-1]), .o_out_fmap(xor_out[976*24*24*bW:977*24*24*bW-1]));
convchan2 c_2_977 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[977*5*5:978*5*5-1]), .o_out_fmap(xor_out[977*24*24*bW:978*24*24*bW-1]));
convchan2 c_2_978 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[978*5*5:979*5*5-1]), .o_out_fmap(xor_out[978*24*24*bW:979*24*24*bW-1]));
convchan2 c_2_979 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[979*5*5:980*5*5-1]), .o_out_fmap(xor_out[979*24*24*bW:980*24*24*bW-1]));
convchan2 c_2_980 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[980*5*5:981*5*5-1]), .o_out_fmap(xor_out[980*24*24*bW:981*24*24*bW-1]));
convchan2 c_2_981 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[981*5*5:982*5*5-1]), .o_out_fmap(xor_out[981*24*24*bW:982*24*24*bW-1]));
convchan2 c_2_982 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[982*5*5:983*5*5-1]), .o_out_fmap(xor_out[982*24*24*bW:983*24*24*bW-1]));
convchan2 c_2_983 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[983*5*5:984*5*5-1]), .o_out_fmap(xor_out[983*24*24*bW:984*24*24*bW-1]));
convchan2 c_2_984 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[984*5*5:985*5*5-1]), .o_out_fmap(xor_out[984*24*24*bW:985*24*24*bW-1]));
convchan2 c_2_985 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[985*5*5:986*5*5-1]), .o_out_fmap(xor_out[985*24*24*bW:986*24*24*bW-1]));
convchan2 c_2_986 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[986*5*5:987*5*5-1]), .o_out_fmap(xor_out[986*24*24*bW:987*24*24*bW-1]));
convchan2 c_2_987 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[987*5*5:988*5*5-1]), .o_out_fmap(xor_out[987*24*24*bW:988*24*24*bW-1]));
convchan2 c_2_988 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[988*5*5:989*5*5-1]), .o_out_fmap(xor_out[988*24*24*bW:989*24*24*bW-1]));
convchan2 c_2_989 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[989*5*5:990*5*5-1]), .o_out_fmap(xor_out[989*24*24*bW:990*24*24*bW-1]));
convchan2 c_2_990 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[990*5*5:991*5*5-1]), .o_out_fmap(xor_out[990*24*24*bW:991*24*24*bW-1]));
convchan2 c_2_991 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[991*5*5:992*5*5-1]), .o_out_fmap(xor_out[991*24*24*bW:992*24*24*bW-1]));
convchan2 c_2_992 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[992*5*5:993*5*5-1]), .o_out_fmap(xor_out[992*24*24*bW:993*24*24*bW-1]));
convchan2 c_2_993 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[993*5*5:994*5*5-1]), .o_out_fmap(xor_out[993*24*24*bW:994*24*24*bW-1]));
convchan2 c_2_994 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[994*5*5:995*5*5-1]), .o_out_fmap(xor_out[994*24*24*bW:995*24*24*bW-1]));
convchan2 c_2_995 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[995*5*5:996*5*5-1]), .o_out_fmap(xor_out[995*24*24*bW:996*24*24*bW-1]));
convchan2 c_2_996 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[996*5*5:997*5*5-1]), .o_out_fmap(xor_out[996*24*24*bW:997*24*24*bW-1]));
convchan2 c_2_997 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[997*5*5:998*5*5-1]), .o_out_fmap(xor_out[997*24*24*bW:998*24*24*bW-1]));
convchan2 c_2_998 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[998*5*5:999*5*5-1]), .o_out_fmap(xor_out[998*24*24*bW:999*24*24*bW-1]));
convchan2 c_2_999 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[999*5*5:1000*5*5-1]), .o_out_fmap(xor_out[999*24*24*bW:1000*24*24*bW-1]));
convchan2 c_2_1000 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[1000*5*5:1001*5*5-1]), .o_out_fmap(xor_out[1000*24*24*bW:1001*24*24*bW-1]));
convchan2 c_2_1001 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[1001*5*5:1002*5*5-1]), .o_out_fmap(xor_out[1001*24*24*bW:1002*24*24*bW-1]));
convchan2 c_2_1002 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[1002*5*5:1003*5*5-1]), .o_out_fmap(xor_out[1002*24*24*bW:1003*24*24*bW-1]));
convchan2 c_2_1003 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[1003*5*5:1004*5*5-1]), .o_out_fmap(xor_out[1003*24*24*bW:1004*24*24*bW-1]));
convchan2 c_2_1004 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[1004*5*5:1005*5*5-1]), .o_out_fmap(xor_out[1004*24*24*bW:1005*24*24*bW-1]));
convchan2 c_2_1005 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[1005*5*5:1006*5*5-1]), .o_out_fmap(xor_out[1005*24*24*bW:1006*24*24*bW-1]));
convchan2 c_2_1006 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[1006*5*5:1007*5*5-1]), .o_out_fmap(xor_out[1006*24*24*bW:1007*24*24*bW-1]));
convchan2 c_2_1007 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[1007*5*5:1008*5*5-1]), .o_out_fmap(xor_out[1007*24*24*bW:1008*24*24*bW-1]));
convchan2 c_2_1008 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[1008*5*5:1009*5*5-1]), .o_out_fmap(xor_out[1008*24*24*bW:1009*24*24*bW-1]));
convchan2 c_2_1009 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[1009*5*5:1010*5*5-1]), .o_out_fmap(xor_out[1009*24*24*bW:1010*24*24*bW-1]));
convchan2 c_2_1010 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[1010*5*5:1011*5*5-1]), .o_out_fmap(xor_out[1010*24*24*bW:1011*24*24*bW-1]));
convchan2 c_2_1011 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[1011*5*5:1012*5*5-1]), .o_out_fmap(xor_out[1011*24*24*bW:1012*24*24*bW-1]));
convchan2 c_2_1012 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[1012*5*5:1013*5*5-1]), .o_out_fmap(xor_out[1012*24*24*bW:1013*24*24*bW-1]));
convchan2 c_2_1013 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[1013*5*5:1014*5*5-1]), .o_out_fmap(xor_out[1013*24*24*bW:1014*24*24*bW-1]));
convchan2 c_2_1014 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[1014*5*5:1015*5*5-1]), .o_out_fmap(xor_out[1014*24*24*bW:1015*24*24*bW-1]));
convchan2 c_2_1015 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[1015*5*5:1016*5*5-1]), .o_out_fmap(xor_out[1015*24*24*bW:1016*24*24*bW-1]));
convchan2 c_2_1016 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[1016*5*5:1017*5*5-1]), .o_out_fmap(xor_out[1016*24*24*bW:1017*24*24*bW-1]));
convchan2 c_2_1017 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[1017*5*5:1018*5*5-1]), .o_out_fmap(xor_out[1017*24*24*bW:1018*24*24*bW-1]));
convchan2 c_2_1018 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[1018*5*5:1019*5*5-1]), .o_out_fmap(xor_out[1018*24*24*bW:1019*24*24*bW-1]));
convchan2 c_2_1019 (.i_image(image[16*12*12:17*12*12*+1]), .i_kernel(kernels[1019*5*5:1020*5*5-1]), .o_out_fmap(xor_out[1019*24*24*bW:1020*24*24*bW-1]));
convchan2 c_2_1020 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1020*5*5:1021*5*5-1]), .o_out_fmap(xor_out[1020*24*24*bW:1021*24*24*bW-1]));
convchan2 c_2_1021 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1021*5*5:1022*5*5-1]), .o_out_fmap(xor_out[1021*24*24*bW:1022*24*24*bW-1]));
convchan2 c_2_1022 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1022*5*5:1023*5*5-1]), .o_out_fmap(xor_out[1022*24*24*bW:1023*24*24*bW-1]));
convchan2 c_2_1023 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1023*5*5:1024*5*5-1]), .o_out_fmap(xor_out[1023*24*24*bW:1024*24*24*bW-1]));
convchan2 c_2_1024 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1024*5*5:1025*5*5-1]), .o_out_fmap(xor_out[1024*24*24*bW:1025*24*24*bW-1]));
convchan2 c_2_1025 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1025*5*5:1026*5*5-1]), .o_out_fmap(xor_out[1025*24*24*bW:1026*24*24*bW-1]));
convchan2 c_2_1026 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1026*5*5:1027*5*5-1]), .o_out_fmap(xor_out[1026*24*24*bW:1027*24*24*bW-1]));
convchan2 c_2_1027 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1027*5*5:1028*5*5-1]), .o_out_fmap(xor_out[1027*24*24*bW:1028*24*24*bW-1]));
convchan2 c_2_1028 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1028*5*5:1029*5*5-1]), .o_out_fmap(xor_out[1028*24*24*bW:1029*24*24*bW-1]));
convchan2 c_2_1029 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1029*5*5:1030*5*5-1]), .o_out_fmap(xor_out[1029*24*24*bW:1030*24*24*bW-1]));
convchan2 c_2_1030 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1030*5*5:1031*5*5-1]), .o_out_fmap(xor_out[1030*24*24*bW:1031*24*24*bW-1]));
convchan2 c_2_1031 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1031*5*5:1032*5*5-1]), .o_out_fmap(xor_out[1031*24*24*bW:1032*24*24*bW-1]));
convchan2 c_2_1032 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1032*5*5:1033*5*5-1]), .o_out_fmap(xor_out[1032*24*24*bW:1033*24*24*bW-1]));
convchan2 c_2_1033 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1033*5*5:1034*5*5-1]), .o_out_fmap(xor_out[1033*24*24*bW:1034*24*24*bW-1]));
convchan2 c_2_1034 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1034*5*5:1035*5*5-1]), .o_out_fmap(xor_out[1034*24*24*bW:1035*24*24*bW-1]));
convchan2 c_2_1035 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1035*5*5:1036*5*5-1]), .o_out_fmap(xor_out[1035*24*24*bW:1036*24*24*bW-1]));
convchan2 c_2_1036 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1036*5*5:1037*5*5-1]), .o_out_fmap(xor_out[1036*24*24*bW:1037*24*24*bW-1]));
convchan2 c_2_1037 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1037*5*5:1038*5*5-1]), .o_out_fmap(xor_out[1037*24*24*bW:1038*24*24*bW-1]));
convchan2 c_2_1038 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1038*5*5:1039*5*5-1]), .o_out_fmap(xor_out[1038*24*24*bW:1039*24*24*bW-1]));
convchan2 c_2_1039 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1039*5*5:1040*5*5-1]), .o_out_fmap(xor_out[1039*24*24*bW:1040*24*24*bW-1]));
convchan2 c_2_1040 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1040*5*5:1041*5*5-1]), .o_out_fmap(xor_out[1040*24*24*bW:1041*24*24*bW-1]));
convchan2 c_2_1041 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1041*5*5:1042*5*5-1]), .o_out_fmap(xor_out[1041*24*24*bW:1042*24*24*bW-1]));
convchan2 c_2_1042 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1042*5*5:1043*5*5-1]), .o_out_fmap(xor_out[1042*24*24*bW:1043*24*24*bW-1]));
convchan2 c_2_1043 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1043*5*5:1044*5*5-1]), .o_out_fmap(xor_out[1043*24*24*bW:1044*24*24*bW-1]));
convchan2 c_2_1044 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1044*5*5:1045*5*5-1]), .o_out_fmap(xor_out[1044*24*24*bW:1045*24*24*bW-1]));
convchan2 c_2_1045 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1045*5*5:1046*5*5-1]), .o_out_fmap(xor_out[1045*24*24*bW:1046*24*24*bW-1]));
convchan2 c_2_1046 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1046*5*5:1047*5*5-1]), .o_out_fmap(xor_out[1046*24*24*bW:1047*24*24*bW-1]));
convchan2 c_2_1047 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1047*5*5:1048*5*5-1]), .o_out_fmap(xor_out[1047*24*24*bW:1048*24*24*bW-1]));
convchan2 c_2_1048 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1048*5*5:1049*5*5-1]), .o_out_fmap(xor_out[1048*24*24*bW:1049*24*24*bW-1]));
convchan2 c_2_1049 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1049*5*5:1050*5*5-1]), .o_out_fmap(xor_out[1049*24*24*bW:1050*24*24*bW-1]));
convchan2 c_2_1050 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1050*5*5:1051*5*5-1]), .o_out_fmap(xor_out[1050*24*24*bW:1051*24*24*bW-1]));
convchan2 c_2_1051 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1051*5*5:1052*5*5-1]), .o_out_fmap(xor_out[1051*24*24*bW:1052*24*24*bW-1]));
convchan2 c_2_1052 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1052*5*5:1053*5*5-1]), .o_out_fmap(xor_out[1052*24*24*bW:1053*24*24*bW-1]));
convchan2 c_2_1053 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1053*5*5:1054*5*5-1]), .o_out_fmap(xor_out[1053*24*24*bW:1054*24*24*bW-1]));
convchan2 c_2_1054 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1054*5*5:1055*5*5-1]), .o_out_fmap(xor_out[1054*24*24*bW:1055*24*24*bW-1]));
convchan2 c_2_1055 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1055*5*5:1056*5*5-1]), .o_out_fmap(xor_out[1055*24*24*bW:1056*24*24*bW-1]));
convchan2 c_2_1056 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1056*5*5:1057*5*5-1]), .o_out_fmap(xor_out[1056*24*24*bW:1057*24*24*bW-1]));
convchan2 c_2_1057 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1057*5*5:1058*5*5-1]), .o_out_fmap(xor_out[1057*24*24*bW:1058*24*24*bW-1]));
convchan2 c_2_1058 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1058*5*5:1059*5*5-1]), .o_out_fmap(xor_out[1058*24*24*bW:1059*24*24*bW-1]));
convchan2 c_2_1059 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1059*5*5:1060*5*5-1]), .o_out_fmap(xor_out[1059*24*24*bW:1060*24*24*bW-1]));
convchan2 c_2_1060 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1060*5*5:1061*5*5-1]), .o_out_fmap(xor_out[1060*24*24*bW:1061*24*24*bW-1]));
convchan2 c_2_1061 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1061*5*5:1062*5*5-1]), .o_out_fmap(xor_out[1061*24*24*bW:1062*24*24*bW-1]));
convchan2 c_2_1062 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1062*5*5:1063*5*5-1]), .o_out_fmap(xor_out[1062*24*24*bW:1063*24*24*bW-1]));
convchan2 c_2_1063 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1063*5*5:1064*5*5-1]), .o_out_fmap(xor_out[1063*24*24*bW:1064*24*24*bW-1]));
convchan2 c_2_1064 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1064*5*5:1065*5*5-1]), .o_out_fmap(xor_out[1064*24*24*bW:1065*24*24*bW-1]));
convchan2 c_2_1065 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1065*5*5:1066*5*5-1]), .o_out_fmap(xor_out[1065*24*24*bW:1066*24*24*bW-1]));
convchan2 c_2_1066 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1066*5*5:1067*5*5-1]), .o_out_fmap(xor_out[1066*24*24*bW:1067*24*24*bW-1]));
convchan2 c_2_1067 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1067*5*5:1068*5*5-1]), .o_out_fmap(xor_out[1067*24*24*bW:1068*24*24*bW-1]));
convchan2 c_2_1068 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1068*5*5:1069*5*5-1]), .o_out_fmap(xor_out[1068*24*24*bW:1069*24*24*bW-1]));
convchan2 c_2_1069 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1069*5*5:1070*5*5-1]), .o_out_fmap(xor_out[1069*24*24*bW:1070*24*24*bW-1]));
convchan2 c_2_1070 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1070*5*5:1071*5*5-1]), .o_out_fmap(xor_out[1070*24*24*bW:1071*24*24*bW-1]));
convchan2 c_2_1071 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1071*5*5:1072*5*5-1]), .o_out_fmap(xor_out[1071*24*24*bW:1072*24*24*bW-1]));
convchan2 c_2_1072 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1072*5*5:1073*5*5-1]), .o_out_fmap(xor_out[1072*24*24*bW:1073*24*24*bW-1]));
convchan2 c_2_1073 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1073*5*5:1074*5*5-1]), .o_out_fmap(xor_out[1073*24*24*bW:1074*24*24*bW-1]));
convchan2 c_2_1074 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1074*5*5:1075*5*5-1]), .o_out_fmap(xor_out[1074*24*24*bW:1075*24*24*bW-1]));
convchan2 c_2_1075 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1075*5*5:1076*5*5-1]), .o_out_fmap(xor_out[1075*24*24*bW:1076*24*24*bW-1]));
convchan2 c_2_1076 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1076*5*5:1077*5*5-1]), .o_out_fmap(xor_out[1076*24*24*bW:1077*24*24*bW-1]));
convchan2 c_2_1077 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1077*5*5:1078*5*5-1]), .o_out_fmap(xor_out[1077*24*24*bW:1078*24*24*bW-1]));
convchan2 c_2_1078 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1078*5*5:1079*5*5-1]), .o_out_fmap(xor_out[1078*24*24*bW:1079*24*24*bW-1]));
convchan2 c_2_1079 (.i_image(image[17*12*12:18*12*12*+1]), .i_kernel(kernels[1079*5*5:1080*5*5-1]), .o_out_fmap(xor_out[1079*24*24*bW:1080*24*24*bW-1]));

accbin2 ab_2_0 (.i_accbin_in(xor_out[0*18*24*24*bW:1*18*24*24*bW-1]), .kernel_offset(kernel_offset[0*bW:1*bW-1]), .o_accbin_out(conv_one_out[0*8*8:1*8*8-1]));
accbin2 ab_2_1 (.i_accbin_in(xor_out[1*18*24*24*bW:2*18*24*24*bW-1]), .kernel_offset(kernel_offset[1*bW:2*bW-1]), .o_accbin_out(conv_one_out[1*8*8:2*8*8-1]));
accbin2 ab_2_2 (.i_accbin_in(xor_out[2*18*24*24*bW:3*18*24*24*bW-1]), .kernel_offset(kernel_offset[2*bW:3*bW-1]), .o_accbin_out(conv_one_out[2*8*8:3*8*8-1]));
accbin2 ab_2_3 (.i_accbin_in(xor_out[3*18*24*24*bW:4*18*24*24*bW-1]), .kernel_offset(kernel_offset[3*bW:4*bW-1]), .o_accbin_out(conv_one_out[3*8*8:4*8*8-1]));
accbin2 ab_2_4 (.i_accbin_in(xor_out[4*18*24*24*bW:5*18*24*24*bW-1]), .kernel_offset(kernel_offset[4*bW:5*bW-1]), .o_accbin_out(conv_one_out[4*8*8:5*8*8-1]));
accbin2 ab_2_5 (.i_accbin_in(xor_out[5*18*24*24*bW:6*18*24*24*bW-1]), .kernel_offset(kernel_offset[5*bW:6*bW-1]), .o_accbin_out(conv_one_out[5*8*8:6*8*8-1]));
accbin2 ab_2_6 (.i_accbin_in(xor_out[6*18*24*24*bW:7*18*24*24*bW-1]), .kernel_offset(kernel_offset[6*bW:7*bW-1]), .o_accbin_out(conv_one_out[6*8*8:7*8*8-1]));
accbin2 ab_2_7 (.i_accbin_in(xor_out[7*18*24*24*bW:8*18*24*24*bW-1]), .kernel_offset(kernel_offset[7*bW:8*bW-1]), .o_accbin_out(conv_one_out[7*8*8:8*8*8-1]));
accbin2 ab_2_8 (.i_accbin_in(xor_out[8*18*24*24*bW:9*18*24*24*bW-1]), .kernel_offset(kernel_offset[8*bW:9*bW-1]), .o_accbin_out(conv_one_out[8*8*8:9*8*8-1]));
accbin2 ab_2_9 (.i_accbin_in(xor_out[9*18*24*24*bW:10*18*24*24*bW-1]), .kernel_offset(kernel_offset[9*bW:10*bW-1]), .o_accbin_out(conv_one_out[9*8*8:10*8*8-1]));
accbin2 ab_2_10 (.i_accbin_in(xor_out[10*18*24*24*bW:11*18*24*24*bW-1]), .kernel_offset(kernel_offset[10*bW:11*bW-1]), .o_accbin_out(conv_one_out[10*8*8:11*8*8-1]));
accbin2 ab_2_11 (.i_accbin_in(xor_out[11*18*24*24*bW:12*18*24*24*bW-1]), .kernel_offset(kernel_offset[11*bW:12*bW-1]), .o_accbin_out(conv_one_out[11*8*8:12*8*8-1]));
accbin2 ab_2_12 (.i_accbin_in(xor_out[12*18*24*24*bW:13*18*24*24*bW-1]), .kernel_offset(kernel_offset[12*bW:13*bW-1]), .o_accbin_out(conv_one_out[12*8*8:13*8*8-1]));
accbin2 ab_2_13 (.i_accbin_in(xor_out[13*18*24*24*bW:14*18*24*24*bW-1]), .kernel_offset(kernel_offset[13*bW:14*bW-1]), .o_accbin_out(conv_one_out[13*8*8:14*8*8-1]));
accbin2 ab_2_14 (.i_accbin_in(xor_out[14*18*24*24*bW:15*18*24*24*bW-1]), .kernel_offset(kernel_offset[14*bW:15*bW-1]), .o_accbin_out(conv_one_out[14*8*8:15*8*8-1]));
accbin2 ab_2_15 (.i_accbin_in(xor_out[15*18*24*24*bW:16*18*24*24*bW-1]), .kernel_offset(kernel_offset[15*bW:16*bW-1]), .o_accbin_out(conv_one_out[15*8*8:16*8*8-1]));
accbin2 ab_2_16 (.i_accbin_in(xor_out[16*18*24*24*bW:17*18*24*24*bW-1]), .kernel_offset(kernel_offset[16*bW:17*bW-1]), .o_accbin_out(conv_one_out[16*8*8:17*8*8-1]));
accbin2 ab_2_17 (.i_accbin_in(xor_out[17*18*24*24*bW:18*18*24*24*bW-1]), .kernel_offset(kernel_offset[17*bW:18*bW-1]), .o_accbin_out(conv_one_out[17*8*8:18*8*8-1]));
accbin2 ab_2_18 (.i_accbin_in(xor_out[18*18*24*24*bW:19*18*24*24*bW-1]), .kernel_offset(kernel_offset[18*bW:19*bW-1]), .o_accbin_out(conv_one_out[18*8*8:19*8*8-1]));
accbin2 ab_2_19 (.i_accbin_in(xor_out[19*18*24*24*bW:20*18*24*24*bW-1]), .kernel_offset(kernel_offset[19*bW:20*bW-1]), .o_accbin_out(conv_one_out[19*8*8:20*8*8-1]));
accbin2 ab_2_20 (.i_accbin_in(xor_out[20*18*24*24*bW:21*18*24*24*bW-1]), .kernel_offset(kernel_offset[20*bW:21*bW-1]), .o_accbin_out(conv_one_out[20*8*8:21*8*8-1]));
accbin2 ab_2_21 (.i_accbin_in(xor_out[21*18*24*24*bW:22*18*24*24*bW-1]), .kernel_offset(kernel_offset[21*bW:22*bW-1]), .o_accbin_out(conv_one_out[21*8*8:22*8*8-1]));
accbin2 ab_2_22 (.i_accbin_in(xor_out[22*18*24*24*bW:23*18*24*24*bW-1]), .kernel_offset(kernel_offset[22*bW:23*bW-1]), .o_accbin_out(conv_one_out[22*8*8:23*8*8-1]));
accbin2 ab_2_23 (.i_accbin_in(xor_out[23*18*24*24*bW:24*18*24*24*bW-1]), .kernel_offset(kernel_offset[23*bW:24*bW-1]), .o_accbin_out(conv_one_out[23*8*8:24*8*8-1]));
accbin2 ab_2_24 (.i_accbin_in(xor_out[24*18*24*24*bW:25*18*24*24*bW-1]), .kernel_offset(kernel_offset[24*bW:25*bW-1]), .o_accbin_out(conv_one_out[24*8*8:25*8*8-1]));
accbin2 ab_2_25 (.i_accbin_in(xor_out[25*18*24*24*bW:26*18*24*24*bW-1]), .kernel_offset(kernel_offset[25*bW:26*bW-1]), .o_accbin_out(conv_one_out[25*8*8:26*8*8-1]));
accbin2 ab_2_26 (.i_accbin_in(xor_out[26*18*24*24*bW:27*18*24*24*bW-1]), .kernel_offset(kernel_offset[26*bW:27*bW-1]), .o_accbin_out(conv_one_out[26*8*8:27*8*8-1]));
accbin2 ab_2_27 (.i_accbin_in(xor_out[27*18*24*24*bW:28*18*24*24*bW-1]), .kernel_offset(kernel_offset[27*bW:28*bW-1]), .o_accbin_out(conv_one_out[27*8*8:28*8*8-1]));
accbin2 ab_2_28 (.i_accbin_in(xor_out[28*18*24*24*bW:29*18*24*24*bW-1]), .kernel_offset(kernel_offset[28*bW:29*bW-1]), .o_accbin_out(conv_one_out[28*8*8:29*8*8-1]));
accbin2 ab_2_29 (.i_accbin_in(xor_out[29*18*24*24*bW:30*18*24*24*bW-1]), .kernel_offset(kernel_offset[29*bW:30*bW-1]), .o_accbin_out(conv_one_out[29*8*8:30*8*8-1]));
accbin2 ab_2_30 (.i_accbin_in(xor_out[30*18*24*24*bW:31*18*24*24*bW-1]), .kernel_offset(kernel_offset[30*bW:31*bW-1]), .o_accbin_out(conv_one_out[30*8*8:31*8*8-1]));
accbin2 ab_2_31 (.i_accbin_in(xor_out[31*18*24*24*bW:32*18*24*24*bW-1]), .kernel_offset(kernel_offset[31*bW:32*bW-1]), .o_accbin_out(conv_one_out[31*8*8:32*8*8-1]));
accbin2 ab_2_32 (.i_accbin_in(xor_out[32*18*24*24*bW:33*18*24*24*bW-1]), .kernel_offset(kernel_offset[32*bW:33*bW-1]), .o_accbin_out(conv_one_out[32*8*8:33*8*8-1]));
accbin2 ab_2_33 (.i_accbin_in(xor_out[33*18*24*24*bW:34*18*24*24*bW-1]), .kernel_offset(kernel_offset[33*bW:34*bW-1]), .o_accbin_out(conv_one_out[33*8*8:34*8*8-1]));
accbin2 ab_2_34 (.i_accbin_in(xor_out[34*18*24*24*bW:35*18*24*24*bW-1]), .kernel_offset(kernel_offset[34*bW:35*bW-1]), .o_accbin_out(conv_one_out[34*8*8:35*8*8-1]));
accbin2 ab_2_35 (.i_accbin_in(xor_out[35*18*24*24*bW:36*18*24*24*bW-1]), .kernel_offset(kernel_offset[35*bW:36*bW-1]), .o_accbin_out(conv_one_out[35*8*8:36*8*8-1]));
accbin2 ab_2_36 (.i_accbin_in(xor_out[36*18*24*24*bW:37*18*24*24*bW-1]), .kernel_offset(kernel_offset[36*bW:37*bW-1]), .o_accbin_out(conv_one_out[36*8*8:37*8*8-1]));
accbin2 ab_2_37 (.i_accbin_in(xor_out[37*18*24*24*bW:38*18*24*24*bW-1]), .kernel_offset(kernel_offset[37*bW:38*bW-1]), .o_accbin_out(conv_one_out[37*8*8:38*8*8-1]));
accbin2 ab_2_38 (.i_accbin_in(xor_out[38*18*24*24*bW:39*18*24*24*bW-1]), .kernel_offset(kernel_offset[38*bW:39*bW-1]), .o_accbin_out(conv_one_out[38*8*8:39*8*8-1]));
accbin2 ab_2_39 (.i_accbin_in(xor_out[39*18*24*24*bW:40*18*24*24*bW-1]), .kernel_offset(kernel_offset[39*bW:40*bW-1]), .o_accbin_out(conv_one_out[39*8*8:40*8*8-1]));
accbin2 ab_2_40 (.i_accbin_in(xor_out[40*18*24*24*bW:41*18*24*24*bW-1]), .kernel_offset(kernel_offset[40*bW:41*bW-1]), .o_accbin_out(conv_one_out[40*8*8:41*8*8-1]));
accbin2 ab_2_41 (.i_accbin_in(xor_out[41*18*24*24*bW:42*18*24*24*bW-1]), .kernel_offset(kernel_offset[41*bW:42*bW-1]), .o_accbin_out(conv_one_out[41*8*8:42*8*8-1]));
accbin2 ab_2_42 (.i_accbin_in(xor_out[42*18*24*24*bW:43*18*24*24*bW-1]), .kernel_offset(kernel_offset[42*bW:43*bW-1]), .o_accbin_out(conv_one_out[42*8*8:43*8*8-1]));
accbin2 ab_2_43 (.i_accbin_in(xor_out[43*18*24*24*bW:44*18*24*24*bW-1]), .kernel_offset(kernel_offset[43*bW:44*bW-1]), .o_accbin_out(conv_one_out[43*8*8:44*8*8-1]));
accbin2 ab_2_44 (.i_accbin_in(xor_out[44*18*24*24*bW:45*18*24*24*bW-1]), .kernel_offset(kernel_offset[44*bW:45*bW-1]), .o_accbin_out(conv_one_out[44*8*8:45*8*8-1]));
accbin2 ab_2_45 (.i_accbin_in(xor_out[45*18*24*24*bW:46*18*24*24*bW-1]), .kernel_offset(kernel_offset[45*bW:46*bW-1]), .o_accbin_out(conv_one_out[45*8*8:46*8*8-1]));
accbin2 ab_2_46 (.i_accbin_in(xor_out[46*18*24*24*bW:47*18*24*24*bW-1]), .kernel_offset(kernel_offset[46*bW:47*bW-1]), .o_accbin_out(conv_one_out[46*8*8:47*8*8-1]));
accbin2 ab_2_47 (.i_accbin_in(xor_out[47*18*24*24*bW:48*18*24*24*bW-1]), .kernel_offset(kernel_offset[47*bW:48*bW-1]), .o_accbin_out(conv_one_out[47*8*8:48*8*8-1]));
accbin2 ab_2_48 (.i_accbin_in(xor_out[48*18*24*24*bW:49*18*24*24*bW-1]), .kernel_offset(kernel_offset[48*bW:49*bW-1]), .o_accbin_out(conv_one_out[48*8*8:49*8*8-1]));
accbin2 ab_2_49 (.i_accbin_in(xor_out[49*18*24*24*bW:50*18*24*24*bW-1]), .kernel_offset(kernel_offset[49*bW:50*bW-1]), .o_accbin_out(conv_one_out[49*8*8:50*8*8-1]));
accbin2 ab_2_50 (.i_accbin_in(xor_out[50*18*24*24*bW:51*18*24*24*bW-1]), .kernel_offset(kernel_offset[50*bW:51*bW-1]), .o_accbin_out(conv_one_out[50*8*8:51*8*8-1]));
accbin2 ab_2_51 (.i_accbin_in(xor_out[51*18*24*24*bW:52*18*24*24*bW-1]), .kernel_offset(kernel_offset[51*bW:52*bW-1]), .o_accbin_out(conv_one_out[51*8*8:52*8*8-1]));
accbin2 ab_2_52 (.i_accbin_in(xor_out[52*18*24*24*bW:53*18*24*24*bW-1]), .kernel_offset(kernel_offset[52*bW:53*bW-1]), .o_accbin_out(conv_one_out[52*8*8:53*8*8-1]));
accbin2 ab_2_53 (.i_accbin_in(xor_out[53*18*24*24*bW:54*18*24*24*bW-1]), .kernel_offset(kernel_offset[53*bW:54*bW-1]), .o_accbin_out(conv_one_out[53*8*8:54*8*8-1]));
accbin2 ab_2_54 (.i_accbin_in(xor_out[54*18*24*24*bW:55*18*24*24*bW-1]), .kernel_offset(kernel_offset[54*bW:55*bW-1]), .o_accbin_out(conv_one_out[54*8*8:55*8*8-1]));
accbin2 ab_2_55 (.i_accbin_in(xor_out[55*18*24*24*bW:56*18*24*24*bW-1]), .kernel_offset(kernel_offset[55*bW:56*bW-1]), .o_accbin_out(conv_one_out[55*8*8:56*8*8-1]));
accbin2 ab_2_56 (.i_accbin_in(xor_out[56*18*24*24*bW:57*18*24*24*bW-1]), .kernel_offset(kernel_offset[56*bW:57*bW-1]), .o_accbin_out(conv_one_out[56*8*8:57*8*8-1]));
accbin2 ab_2_57 (.i_accbin_in(xor_out[57*18*24*24*bW:58*18*24*24*bW-1]), .kernel_offset(kernel_offset[57*bW:58*bW-1]), .o_accbin_out(conv_one_out[57*8*8:58*8*8-1]));
accbin2 ab_2_58 (.i_accbin_in(xor_out[58*18*24*24*bW:59*18*24*24*bW-1]), .kernel_offset(kernel_offset[58*bW:59*bW-1]), .o_accbin_out(conv_one_out[58*8*8:59*8*8-1]));
accbin2 ab_2_59 (.i_accbin_in(xor_out[59*18*24*24*bW:60*18*24*24*bW-1]), .kernel_offset(kernel_offset[59*bW:60*bW-1]), .o_accbin_out(conv_one_out[59*8*8:60*8*8-1]));

endmodule