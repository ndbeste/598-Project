module conv2
    #( parameter bW = 8 )
    (
    input  logic            image          [0:  17][0:11][0:11],
    input  logic            kernels        [0:1079][0: 4][0: 4],
    input  logic  [bW-1:0]  kernel_offset  [0:  59],
    output logic            conv_two_out   [0:  59][0: 7][0: 7]
    );

logic       xor_out [0:1079][0:23][0:23];

convchan2 c_2_0 (.image, .kernel(kernels[0]), .conv_out(xor_out[0]));
convchan2 c_2_1 (.image, .kernel(kernels[1]), .conv_out(xor_out[1]));
convchan2 c_2_2 (.image, .kernel(kernels[2]), .conv_out(xor_out[2]));
convchan2 c_2_3 (.image, .kernel(kernels[3]), .conv_out(xor_out[3]));
convchan2 c_2_4 (.image, .kernel(kernels[4]), .conv_out(xor_out[4]));
convchan2 c_2_5 (.image, .kernel(kernels[5]), .conv_out(xor_out[5]));
convchan2 c_2_6 (.image, .kernel(kernels[6]), .conv_out(xor_out[6]));
convchan2 c_2_7 (.image, .kernel(kernels[7]), .conv_out(xor_out[7]));
convchan2 c_2_8 (.image, .kernel(kernels[8]), .conv_out(xor_out[8]));
convchan2 c_2_9 (.image, .kernel(kernels[9]), .conv_out(xor_out[9]));
convchan2 c_2_10 (.image, .kernel(kernels[10]), .conv_out(xor_out[10]));
convchan2 c_2_11 (.image, .kernel(kernels[11]), .conv_out(xor_out[11]));
convchan2 c_2_12 (.image, .kernel(kernels[12]), .conv_out(xor_out[12]));
convchan2 c_2_13 (.image, .kernel(kernels[13]), .conv_out(xor_out[13]));
convchan2 c_2_14 (.image, .kernel(kernels[14]), .conv_out(xor_out[14]));
convchan2 c_2_15 (.image, .kernel(kernels[15]), .conv_out(xor_out[15]));
convchan2 c_2_16 (.image, .kernel(kernels[16]), .conv_out(xor_out[16]));
convchan2 c_2_17 (.image, .kernel(kernels[17]), .conv_out(xor_out[17]));
convchan2 c_2_18 (.image, .kernel(kernels[18]), .conv_out(xor_out[18]));
convchan2 c_2_19 (.image, .kernel(kernels[19]), .conv_out(xor_out[19]));
convchan2 c_2_20 (.image, .kernel(kernels[20]), .conv_out(xor_out[20]));
convchan2 c_2_21 (.image, .kernel(kernels[21]), .conv_out(xor_out[21]));
convchan2 c_2_22 (.image, .kernel(kernels[22]), .conv_out(xor_out[22]));
convchan2 c_2_23 (.image, .kernel(kernels[23]), .conv_out(xor_out[23]));
convchan2 c_2_24 (.image, .kernel(kernels[24]), .conv_out(xor_out[24]));
convchan2 c_2_25 (.image, .kernel(kernels[25]), .conv_out(xor_out[25]));
convchan2 c_2_26 (.image, .kernel(kernels[26]), .conv_out(xor_out[26]));
convchan2 c_2_27 (.image, .kernel(kernels[27]), .conv_out(xor_out[27]));
convchan2 c_2_28 (.image, .kernel(kernels[28]), .conv_out(xor_out[28]));
convchan2 c_2_29 (.image, .kernel(kernels[29]), .conv_out(xor_out[29]));
convchan2 c_2_30 (.image, .kernel(kernels[30]), .conv_out(xor_out[30]));
convchan2 c_2_31 (.image, .kernel(kernels[31]), .conv_out(xor_out[31]));
convchan2 c_2_32 (.image, .kernel(kernels[32]), .conv_out(xor_out[32]));
convchan2 c_2_33 (.image, .kernel(kernels[33]), .conv_out(xor_out[33]));
convchan2 c_2_34 (.image, .kernel(kernels[34]), .conv_out(xor_out[34]));
convchan2 c_2_35 (.image, .kernel(kernels[35]), .conv_out(xor_out[35]));
convchan2 c_2_36 (.image, .kernel(kernels[36]), .conv_out(xor_out[36]));
convchan2 c_2_37 (.image, .kernel(kernels[37]), .conv_out(xor_out[37]));
convchan2 c_2_38 (.image, .kernel(kernels[38]), .conv_out(xor_out[38]));
convchan2 c_2_39 (.image, .kernel(kernels[39]), .conv_out(xor_out[39]));
convchan2 c_2_40 (.image, .kernel(kernels[40]), .conv_out(xor_out[40]));
convchan2 c_2_41 (.image, .kernel(kernels[41]), .conv_out(xor_out[41]));
convchan2 c_2_42 (.image, .kernel(kernels[42]), .conv_out(xor_out[42]));
convchan2 c_2_43 (.image, .kernel(kernels[43]), .conv_out(xor_out[43]));
convchan2 c_2_44 (.image, .kernel(kernels[44]), .conv_out(xor_out[44]));
convchan2 c_2_45 (.image, .kernel(kernels[45]), .conv_out(xor_out[45]));
convchan2 c_2_46 (.image, .kernel(kernels[46]), .conv_out(xor_out[46]));
convchan2 c_2_47 (.image, .kernel(kernels[47]), .conv_out(xor_out[47]));
convchan2 c_2_48 (.image, .kernel(kernels[48]), .conv_out(xor_out[48]));
convchan2 c_2_49 (.image, .kernel(kernels[49]), .conv_out(xor_out[49]));
convchan2 c_2_50 (.image, .kernel(kernels[50]), .conv_out(xor_out[50]));
convchan2 c_2_51 (.image, .kernel(kernels[51]), .conv_out(xor_out[51]));
convchan2 c_2_52 (.image, .kernel(kernels[52]), .conv_out(xor_out[52]));
convchan2 c_2_53 (.image, .kernel(kernels[53]), .conv_out(xor_out[53]));
convchan2 c_2_54 (.image, .kernel(kernels[54]), .conv_out(xor_out[54]));
convchan2 c_2_55 (.image, .kernel(kernels[55]), .conv_out(xor_out[55]));
convchan2 c_2_56 (.image, .kernel(kernels[56]), .conv_out(xor_out[56]));
convchan2 c_2_57 (.image, .kernel(kernels[57]), .conv_out(xor_out[57]));
convchan2 c_2_58 (.image, .kernel(kernels[58]), .conv_out(xor_out[58]));
convchan2 c_2_59 (.image, .kernel(kernels[59]), .conv_out(xor_out[59]));
convchan2 c_2_60 (.image, .kernel(kernels[60]), .conv_out(xor_out[60]));
convchan2 c_2_61 (.image, .kernel(kernels[61]), .conv_out(xor_out[61]));
convchan2 c_2_62 (.image, .kernel(kernels[62]), .conv_out(xor_out[62]));
convchan2 c_2_63 (.image, .kernel(kernels[63]), .conv_out(xor_out[63]));
convchan2 c_2_64 (.image, .kernel(kernels[64]), .conv_out(xor_out[64]));
convchan2 c_2_65 (.image, .kernel(kernels[65]), .conv_out(xor_out[65]));
convchan2 c_2_66 (.image, .kernel(kernels[66]), .conv_out(xor_out[66]));
convchan2 c_2_67 (.image, .kernel(kernels[67]), .conv_out(xor_out[67]));
convchan2 c_2_68 (.image, .kernel(kernels[68]), .conv_out(xor_out[68]));
convchan2 c_2_69 (.image, .kernel(kernels[69]), .conv_out(xor_out[69]));
convchan2 c_2_70 (.image, .kernel(kernels[70]), .conv_out(xor_out[70]));
convchan2 c_2_71 (.image, .kernel(kernels[71]), .conv_out(xor_out[71]));
convchan2 c_2_72 (.image, .kernel(kernels[72]), .conv_out(xor_out[72]));
convchan2 c_2_73 (.image, .kernel(kernels[73]), .conv_out(xor_out[73]));
convchan2 c_2_74 (.image, .kernel(kernels[74]), .conv_out(xor_out[74]));
convchan2 c_2_75 (.image, .kernel(kernels[75]), .conv_out(xor_out[75]));
convchan2 c_2_76 (.image, .kernel(kernels[76]), .conv_out(xor_out[76]));
convchan2 c_2_77 (.image, .kernel(kernels[77]), .conv_out(xor_out[77]));
convchan2 c_2_78 (.image, .kernel(kernels[78]), .conv_out(xor_out[78]));
convchan2 c_2_79 (.image, .kernel(kernels[79]), .conv_out(xor_out[79]));
convchan2 c_2_80 (.image, .kernel(kernels[80]), .conv_out(xor_out[80]));
convchan2 c_2_81 (.image, .kernel(kernels[81]), .conv_out(xor_out[81]));
convchan2 c_2_82 (.image, .kernel(kernels[82]), .conv_out(xor_out[82]));
convchan2 c_2_83 (.image, .kernel(kernels[83]), .conv_out(xor_out[83]));
convchan2 c_2_84 (.image, .kernel(kernels[84]), .conv_out(xor_out[84]));
convchan2 c_2_85 (.image, .kernel(kernels[85]), .conv_out(xor_out[85]));
convchan2 c_2_86 (.image, .kernel(kernels[86]), .conv_out(xor_out[86]));
convchan2 c_2_87 (.image, .kernel(kernels[87]), .conv_out(xor_out[87]));
convchan2 c_2_88 (.image, .kernel(kernels[88]), .conv_out(xor_out[88]));
convchan2 c_2_89 (.image, .kernel(kernels[89]), .conv_out(xor_out[89]));
convchan2 c_2_90 (.image, .kernel(kernels[90]), .conv_out(xor_out[90]));
convchan2 c_2_91 (.image, .kernel(kernels[91]), .conv_out(xor_out[91]));
convchan2 c_2_92 (.image, .kernel(kernels[92]), .conv_out(xor_out[92]));
convchan2 c_2_93 (.image, .kernel(kernels[93]), .conv_out(xor_out[93]));
convchan2 c_2_94 (.image, .kernel(kernels[94]), .conv_out(xor_out[94]));
convchan2 c_2_95 (.image, .kernel(kernels[95]), .conv_out(xor_out[95]));
convchan2 c_2_96 (.image, .kernel(kernels[96]), .conv_out(xor_out[96]));
convchan2 c_2_97 (.image, .kernel(kernels[97]), .conv_out(xor_out[97]));
convchan2 c_2_98 (.image, .kernel(kernels[98]), .conv_out(xor_out[98]));
convchan2 c_2_99 (.image, .kernel(kernels[99]), .conv_out(xor_out[99]));
convchan2 c_2_100 (.image, .kernel(kernels[100]), .conv_out(xor_out[100]));
convchan2 c_2_101 (.image, .kernel(kernels[101]), .conv_out(xor_out[101]));
convchan2 c_2_102 (.image, .kernel(kernels[102]), .conv_out(xor_out[102]));
convchan2 c_2_103 (.image, .kernel(kernels[103]), .conv_out(xor_out[103]));
convchan2 c_2_104 (.image, .kernel(kernels[104]), .conv_out(xor_out[104]));
convchan2 c_2_105 (.image, .kernel(kernels[105]), .conv_out(xor_out[105]));
convchan2 c_2_106 (.image, .kernel(kernels[106]), .conv_out(xor_out[106]));
convchan2 c_2_107 (.image, .kernel(kernels[107]), .conv_out(xor_out[107]));
convchan2 c_2_108 (.image, .kernel(kernels[108]), .conv_out(xor_out[108]));
convchan2 c_2_109 (.image, .kernel(kernels[109]), .conv_out(xor_out[109]));
convchan2 c_2_110 (.image, .kernel(kernels[110]), .conv_out(xor_out[110]));
convchan2 c_2_111 (.image, .kernel(kernels[111]), .conv_out(xor_out[111]));
convchan2 c_2_112 (.image, .kernel(kernels[112]), .conv_out(xor_out[112]));
convchan2 c_2_113 (.image, .kernel(kernels[113]), .conv_out(xor_out[113]));
convchan2 c_2_114 (.image, .kernel(kernels[114]), .conv_out(xor_out[114]));
convchan2 c_2_115 (.image, .kernel(kernels[115]), .conv_out(xor_out[115]));
convchan2 c_2_116 (.image, .kernel(kernels[116]), .conv_out(xor_out[116]));
convchan2 c_2_117 (.image, .kernel(kernels[117]), .conv_out(xor_out[117]));
convchan2 c_2_118 (.image, .kernel(kernels[118]), .conv_out(xor_out[118]));
convchan2 c_2_119 (.image, .kernel(kernels[119]), .conv_out(xor_out[119]));
convchan2 c_2_120 (.image, .kernel(kernels[120]), .conv_out(xor_out[120]));
convchan2 c_2_121 (.image, .kernel(kernels[121]), .conv_out(xor_out[121]));
convchan2 c_2_122 (.image, .kernel(kernels[122]), .conv_out(xor_out[122]));
convchan2 c_2_123 (.image, .kernel(kernels[123]), .conv_out(xor_out[123]));
convchan2 c_2_124 (.image, .kernel(kernels[124]), .conv_out(xor_out[124]));
convchan2 c_2_125 (.image, .kernel(kernels[125]), .conv_out(xor_out[125]));
convchan2 c_2_126 (.image, .kernel(kernels[126]), .conv_out(xor_out[126]));
convchan2 c_2_127 (.image, .kernel(kernels[127]), .conv_out(xor_out[127]));
convchan2 c_2_128 (.image, .kernel(kernels[128]), .conv_out(xor_out[128]));
convchan2 c_2_129 (.image, .kernel(kernels[129]), .conv_out(xor_out[129]));
convchan2 c_2_130 (.image, .kernel(kernels[130]), .conv_out(xor_out[130]));
convchan2 c_2_131 (.image, .kernel(kernels[131]), .conv_out(xor_out[131]));
convchan2 c_2_132 (.image, .kernel(kernels[132]), .conv_out(xor_out[132]));
convchan2 c_2_133 (.image, .kernel(kernels[133]), .conv_out(xor_out[133]));
convchan2 c_2_134 (.image, .kernel(kernels[134]), .conv_out(xor_out[134]));
convchan2 c_2_135 (.image, .kernel(kernels[135]), .conv_out(xor_out[135]));
convchan2 c_2_136 (.image, .kernel(kernels[136]), .conv_out(xor_out[136]));
convchan2 c_2_137 (.image, .kernel(kernels[137]), .conv_out(xor_out[137]));
convchan2 c_2_138 (.image, .kernel(kernels[138]), .conv_out(xor_out[138]));
convchan2 c_2_139 (.image, .kernel(kernels[139]), .conv_out(xor_out[139]));
convchan2 c_2_140 (.image, .kernel(kernels[140]), .conv_out(xor_out[140]));
convchan2 c_2_141 (.image, .kernel(kernels[141]), .conv_out(xor_out[141]));
convchan2 c_2_142 (.image, .kernel(kernels[142]), .conv_out(xor_out[142]));
convchan2 c_2_143 (.image, .kernel(kernels[143]), .conv_out(xor_out[143]));
convchan2 c_2_144 (.image, .kernel(kernels[144]), .conv_out(xor_out[144]));
convchan2 c_2_145 (.image, .kernel(kernels[145]), .conv_out(xor_out[145]));
convchan2 c_2_146 (.image, .kernel(kernels[146]), .conv_out(xor_out[146]));
convchan2 c_2_147 (.image, .kernel(kernels[147]), .conv_out(xor_out[147]));
convchan2 c_2_148 (.image, .kernel(kernels[148]), .conv_out(xor_out[148]));
convchan2 c_2_149 (.image, .kernel(kernels[149]), .conv_out(xor_out[149]));
convchan2 c_2_150 (.image, .kernel(kernels[150]), .conv_out(xor_out[150]));
convchan2 c_2_151 (.image, .kernel(kernels[151]), .conv_out(xor_out[151]));
convchan2 c_2_152 (.image, .kernel(kernels[152]), .conv_out(xor_out[152]));
convchan2 c_2_153 (.image, .kernel(kernels[153]), .conv_out(xor_out[153]));
convchan2 c_2_154 (.image, .kernel(kernels[154]), .conv_out(xor_out[154]));
convchan2 c_2_155 (.image, .kernel(kernels[155]), .conv_out(xor_out[155]));
convchan2 c_2_156 (.image, .kernel(kernels[156]), .conv_out(xor_out[156]));
convchan2 c_2_157 (.image, .kernel(kernels[157]), .conv_out(xor_out[157]));
convchan2 c_2_158 (.image, .kernel(kernels[158]), .conv_out(xor_out[158]));
convchan2 c_2_159 (.image, .kernel(kernels[159]), .conv_out(xor_out[159]));
convchan2 c_2_160 (.image, .kernel(kernels[160]), .conv_out(xor_out[160]));
convchan2 c_2_161 (.image, .kernel(kernels[161]), .conv_out(xor_out[161]));
convchan2 c_2_162 (.image, .kernel(kernels[162]), .conv_out(xor_out[162]));
convchan2 c_2_163 (.image, .kernel(kernels[163]), .conv_out(xor_out[163]));
convchan2 c_2_164 (.image, .kernel(kernels[164]), .conv_out(xor_out[164]));
convchan2 c_2_165 (.image, .kernel(kernels[165]), .conv_out(xor_out[165]));
convchan2 c_2_166 (.image, .kernel(kernels[166]), .conv_out(xor_out[166]));
convchan2 c_2_167 (.image, .kernel(kernels[167]), .conv_out(xor_out[167]));
convchan2 c_2_168 (.image, .kernel(kernels[168]), .conv_out(xor_out[168]));
convchan2 c_2_169 (.image, .kernel(kernels[169]), .conv_out(xor_out[169]));
convchan2 c_2_170 (.image, .kernel(kernels[170]), .conv_out(xor_out[170]));
convchan2 c_2_171 (.image, .kernel(kernels[171]), .conv_out(xor_out[171]));
convchan2 c_2_172 (.image, .kernel(kernels[172]), .conv_out(xor_out[172]));
convchan2 c_2_173 (.image, .kernel(kernels[173]), .conv_out(xor_out[173]));
convchan2 c_2_174 (.image, .kernel(kernels[174]), .conv_out(xor_out[174]));
convchan2 c_2_175 (.image, .kernel(kernels[175]), .conv_out(xor_out[175]));
convchan2 c_2_176 (.image, .kernel(kernels[176]), .conv_out(xor_out[176]));
convchan2 c_2_177 (.image, .kernel(kernels[177]), .conv_out(xor_out[177]));
convchan2 c_2_178 (.image, .kernel(kernels[178]), .conv_out(xor_out[178]));
convchan2 c_2_179 (.image, .kernel(kernels[179]), .conv_out(xor_out[179]));
convchan2 c_2_180 (.image, .kernel(kernels[180]), .conv_out(xor_out[180]));
convchan2 c_2_181 (.image, .kernel(kernels[181]), .conv_out(xor_out[181]));
convchan2 c_2_182 (.image, .kernel(kernels[182]), .conv_out(xor_out[182]));
convchan2 c_2_183 (.image, .kernel(kernels[183]), .conv_out(xor_out[183]));
convchan2 c_2_184 (.image, .kernel(kernels[184]), .conv_out(xor_out[184]));
convchan2 c_2_185 (.image, .kernel(kernels[185]), .conv_out(xor_out[185]));
convchan2 c_2_186 (.image, .kernel(kernels[186]), .conv_out(xor_out[186]));
convchan2 c_2_187 (.image, .kernel(kernels[187]), .conv_out(xor_out[187]));
convchan2 c_2_188 (.image, .kernel(kernels[188]), .conv_out(xor_out[188]));
convchan2 c_2_189 (.image, .kernel(kernels[189]), .conv_out(xor_out[189]));
convchan2 c_2_190 (.image, .kernel(kernels[190]), .conv_out(xor_out[190]));
convchan2 c_2_191 (.image, .kernel(kernels[191]), .conv_out(xor_out[191]));
convchan2 c_2_192 (.image, .kernel(kernels[192]), .conv_out(xor_out[192]));
convchan2 c_2_193 (.image, .kernel(kernels[193]), .conv_out(xor_out[193]));
convchan2 c_2_194 (.image, .kernel(kernels[194]), .conv_out(xor_out[194]));
convchan2 c_2_195 (.image, .kernel(kernels[195]), .conv_out(xor_out[195]));
convchan2 c_2_196 (.image, .kernel(kernels[196]), .conv_out(xor_out[196]));
convchan2 c_2_197 (.image, .kernel(kernels[197]), .conv_out(xor_out[197]));
convchan2 c_2_198 (.image, .kernel(kernels[198]), .conv_out(xor_out[198]));
convchan2 c_2_199 (.image, .kernel(kernels[199]), .conv_out(xor_out[199]));
convchan2 c_2_200 (.image, .kernel(kernels[200]), .conv_out(xor_out[200]));
convchan2 c_2_201 (.image, .kernel(kernels[201]), .conv_out(xor_out[201]));
convchan2 c_2_202 (.image, .kernel(kernels[202]), .conv_out(xor_out[202]));
convchan2 c_2_203 (.image, .kernel(kernels[203]), .conv_out(xor_out[203]));
convchan2 c_2_204 (.image, .kernel(kernels[204]), .conv_out(xor_out[204]));
convchan2 c_2_205 (.image, .kernel(kernels[205]), .conv_out(xor_out[205]));
convchan2 c_2_206 (.image, .kernel(kernels[206]), .conv_out(xor_out[206]));
convchan2 c_2_207 (.image, .kernel(kernels[207]), .conv_out(xor_out[207]));
convchan2 c_2_208 (.image, .kernel(kernels[208]), .conv_out(xor_out[208]));
convchan2 c_2_209 (.image, .kernel(kernels[209]), .conv_out(xor_out[209]));
convchan2 c_2_210 (.image, .kernel(kernels[210]), .conv_out(xor_out[210]));
convchan2 c_2_211 (.image, .kernel(kernels[211]), .conv_out(xor_out[211]));
convchan2 c_2_212 (.image, .kernel(kernels[212]), .conv_out(xor_out[212]));
convchan2 c_2_213 (.image, .kernel(kernels[213]), .conv_out(xor_out[213]));
convchan2 c_2_214 (.image, .kernel(kernels[214]), .conv_out(xor_out[214]));
convchan2 c_2_215 (.image, .kernel(kernels[215]), .conv_out(xor_out[215]));
convchan2 c_2_216 (.image, .kernel(kernels[216]), .conv_out(xor_out[216]));
convchan2 c_2_217 (.image, .kernel(kernels[217]), .conv_out(xor_out[217]));
convchan2 c_2_218 (.image, .kernel(kernels[218]), .conv_out(xor_out[218]));
convchan2 c_2_219 (.image, .kernel(kernels[219]), .conv_out(xor_out[219]));
convchan2 c_2_220 (.image, .kernel(kernels[220]), .conv_out(xor_out[220]));
convchan2 c_2_221 (.image, .kernel(kernels[221]), .conv_out(xor_out[221]));
convchan2 c_2_222 (.image, .kernel(kernels[222]), .conv_out(xor_out[222]));
convchan2 c_2_223 (.image, .kernel(kernels[223]), .conv_out(xor_out[223]));
convchan2 c_2_224 (.image, .kernel(kernels[224]), .conv_out(xor_out[224]));
convchan2 c_2_225 (.image, .kernel(kernels[225]), .conv_out(xor_out[225]));
convchan2 c_2_226 (.image, .kernel(kernels[226]), .conv_out(xor_out[226]));
convchan2 c_2_227 (.image, .kernel(kernels[227]), .conv_out(xor_out[227]));
convchan2 c_2_228 (.image, .kernel(kernels[228]), .conv_out(xor_out[228]));
convchan2 c_2_229 (.image, .kernel(kernels[229]), .conv_out(xor_out[229]));
convchan2 c_2_230 (.image, .kernel(kernels[230]), .conv_out(xor_out[230]));
convchan2 c_2_231 (.image, .kernel(kernels[231]), .conv_out(xor_out[231]));
convchan2 c_2_232 (.image, .kernel(kernels[232]), .conv_out(xor_out[232]));
convchan2 c_2_233 (.image, .kernel(kernels[233]), .conv_out(xor_out[233]));
convchan2 c_2_234 (.image, .kernel(kernels[234]), .conv_out(xor_out[234]));
convchan2 c_2_235 (.image, .kernel(kernels[235]), .conv_out(xor_out[235]));
convchan2 c_2_236 (.image, .kernel(kernels[236]), .conv_out(xor_out[236]));
convchan2 c_2_237 (.image, .kernel(kernels[237]), .conv_out(xor_out[237]));
convchan2 c_2_238 (.image, .kernel(kernels[238]), .conv_out(xor_out[238]));
convchan2 c_2_239 (.image, .kernel(kernels[239]), .conv_out(xor_out[239]));
convchan2 c_2_240 (.image, .kernel(kernels[240]), .conv_out(xor_out[240]));
convchan2 c_2_241 (.image, .kernel(kernels[241]), .conv_out(xor_out[241]));
convchan2 c_2_242 (.image, .kernel(kernels[242]), .conv_out(xor_out[242]));
convchan2 c_2_243 (.image, .kernel(kernels[243]), .conv_out(xor_out[243]));
convchan2 c_2_244 (.image, .kernel(kernels[244]), .conv_out(xor_out[244]));
convchan2 c_2_245 (.image, .kernel(kernels[245]), .conv_out(xor_out[245]));
convchan2 c_2_246 (.image, .kernel(kernels[246]), .conv_out(xor_out[246]));
convchan2 c_2_247 (.image, .kernel(kernels[247]), .conv_out(xor_out[247]));
convchan2 c_2_248 (.image, .kernel(kernels[248]), .conv_out(xor_out[248]));
convchan2 c_2_249 (.image, .kernel(kernels[249]), .conv_out(xor_out[249]));
convchan2 c_2_250 (.image, .kernel(kernels[250]), .conv_out(xor_out[250]));
convchan2 c_2_251 (.image, .kernel(kernels[251]), .conv_out(xor_out[251]));
convchan2 c_2_252 (.image, .kernel(kernels[252]), .conv_out(xor_out[252]));
convchan2 c_2_253 (.image, .kernel(kernels[253]), .conv_out(xor_out[253]));
convchan2 c_2_254 (.image, .kernel(kernels[254]), .conv_out(xor_out[254]));
convchan2 c_2_255 (.image, .kernel(kernels[255]), .conv_out(xor_out[255]));
convchan2 c_2_256 (.image, .kernel(kernels[256]), .conv_out(xor_out[256]));
convchan2 c_2_257 (.image, .kernel(kernels[257]), .conv_out(xor_out[257]));
convchan2 c_2_258 (.image, .kernel(kernels[258]), .conv_out(xor_out[258]));
convchan2 c_2_259 (.image, .kernel(kernels[259]), .conv_out(xor_out[259]));
convchan2 c_2_260 (.image, .kernel(kernels[260]), .conv_out(xor_out[260]));
convchan2 c_2_261 (.image, .kernel(kernels[261]), .conv_out(xor_out[261]));
convchan2 c_2_262 (.image, .kernel(kernels[262]), .conv_out(xor_out[262]));
convchan2 c_2_263 (.image, .kernel(kernels[263]), .conv_out(xor_out[263]));
convchan2 c_2_264 (.image, .kernel(kernels[264]), .conv_out(xor_out[264]));
convchan2 c_2_265 (.image, .kernel(kernels[265]), .conv_out(xor_out[265]));
convchan2 c_2_266 (.image, .kernel(kernels[266]), .conv_out(xor_out[266]));
convchan2 c_2_267 (.image, .kernel(kernels[267]), .conv_out(xor_out[267]));
convchan2 c_2_268 (.image, .kernel(kernels[268]), .conv_out(xor_out[268]));
convchan2 c_2_269 (.image, .kernel(kernels[269]), .conv_out(xor_out[269]));
convchan2 c_2_270 (.image, .kernel(kernels[270]), .conv_out(xor_out[270]));
convchan2 c_2_271 (.image, .kernel(kernels[271]), .conv_out(xor_out[271]));
convchan2 c_2_272 (.image, .kernel(kernels[272]), .conv_out(xor_out[272]));
convchan2 c_2_273 (.image, .kernel(kernels[273]), .conv_out(xor_out[273]));
convchan2 c_2_274 (.image, .kernel(kernels[274]), .conv_out(xor_out[274]));
convchan2 c_2_275 (.image, .kernel(kernels[275]), .conv_out(xor_out[275]));
convchan2 c_2_276 (.image, .kernel(kernels[276]), .conv_out(xor_out[276]));
convchan2 c_2_277 (.image, .kernel(kernels[277]), .conv_out(xor_out[277]));
convchan2 c_2_278 (.image, .kernel(kernels[278]), .conv_out(xor_out[278]));
convchan2 c_2_279 (.image, .kernel(kernels[279]), .conv_out(xor_out[279]));
convchan2 c_2_280 (.image, .kernel(kernels[280]), .conv_out(xor_out[280]));
convchan2 c_2_281 (.image, .kernel(kernels[281]), .conv_out(xor_out[281]));
convchan2 c_2_282 (.image, .kernel(kernels[282]), .conv_out(xor_out[282]));
convchan2 c_2_283 (.image, .kernel(kernels[283]), .conv_out(xor_out[283]));
convchan2 c_2_284 (.image, .kernel(kernels[284]), .conv_out(xor_out[284]));
convchan2 c_2_285 (.image, .kernel(kernels[285]), .conv_out(xor_out[285]));
convchan2 c_2_286 (.image, .kernel(kernels[286]), .conv_out(xor_out[286]));
convchan2 c_2_287 (.image, .kernel(kernels[287]), .conv_out(xor_out[287]));
convchan2 c_2_288 (.image, .kernel(kernels[288]), .conv_out(xor_out[288]));
convchan2 c_2_289 (.image, .kernel(kernels[289]), .conv_out(xor_out[289]));
convchan2 c_2_290 (.image, .kernel(kernels[290]), .conv_out(xor_out[290]));
convchan2 c_2_291 (.image, .kernel(kernels[291]), .conv_out(xor_out[291]));
convchan2 c_2_292 (.image, .kernel(kernels[292]), .conv_out(xor_out[292]));
convchan2 c_2_293 (.image, .kernel(kernels[293]), .conv_out(xor_out[293]));
convchan2 c_2_294 (.image, .kernel(kernels[294]), .conv_out(xor_out[294]));
convchan2 c_2_295 (.image, .kernel(kernels[295]), .conv_out(xor_out[295]));
convchan2 c_2_296 (.image, .kernel(kernels[296]), .conv_out(xor_out[296]));
convchan2 c_2_297 (.image, .kernel(kernels[297]), .conv_out(xor_out[297]));
convchan2 c_2_298 (.image, .kernel(kernels[298]), .conv_out(xor_out[298]));
convchan2 c_2_299 (.image, .kernel(kernels[299]), .conv_out(xor_out[299]));
convchan2 c_2_300 (.image, .kernel(kernels[300]), .conv_out(xor_out[300]));
convchan2 c_2_301 (.image, .kernel(kernels[301]), .conv_out(xor_out[301]));
convchan2 c_2_302 (.image, .kernel(kernels[302]), .conv_out(xor_out[302]));
convchan2 c_2_303 (.image, .kernel(kernels[303]), .conv_out(xor_out[303]));
convchan2 c_2_304 (.image, .kernel(kernels[304]), .conv_out(xor_out[304]));
convchan2 c_2_305 (.image, .kernel(kernels[305]), .conv_out(xor_out[305]));
convchan2 c_2_306 (.image, .kernel(kernels[306]), .conv_out(xor_out[306]));
convchan2 c_2_307 (.image, .kernel(kernels[307]), .conv_out(xor_out[307]));
convchan2 c_2_308 (.image, .kernel(kernels[308]), .conv_out(xor_out[308]));
convchan2 c_2_309 (.image, .kernel(kernels[309]), .conv_out(xor_out[309]));
convchan2 c_2_310 (.image, .kernel(kernels[310]), .conv_out(xor_out[310]));
convchan2 c_2_311 (.image, .kernel(kernels[311]), .conv_out(xor_out[311]));
convchan2 c_2_312 (.image, .kernel(kernels[312]), .conv_out(xor_out[312]));
convchan2 c_2_313 (.image, .kernel(kernels[313]), .conv_out(xor_out[313]));
convchan2 c_2_314 (.image, .kernel(kernels[314]), .conv_out(xor_out[314]));
convchan2 c_2_315 (.image, .kernel(kernels[315]), .conv_out(xor_out[315]));
convchan2 c_2_316 (.image, .kernel(kernels[316]), .conv_out(xor_out[316]));
convchan2 c_2_317 (.image, .kernel(kernels[317]), .conv_out(xor_out[317]));
convchan2 c_2_318 (.image, .kernel(kernels[318]), .conv_out(xor_out[318]));
convchan2 c_2_319 (.image, .kernel(kernels[319]), .conv_out(xor_out[319]));
convchan2 c_2_320 (.image, .kernel(kernels[320]), .conv_out(xor_out[320]));
convchan2 c_2_321 (.image, .kernel(kernels[321]), .conv_out(xor_out[321]));
convchan2 c_2_322 (.image, .kernel(kernels[322]), .conv_out(xor_out[322]));
convchan2 c_2_323 (.image, .kernel(kernels[323]), .conv_out(xor_out[323]));
convchan2 c_2_324 (.image, .kernel(kernels[324]), .conv_out(xor_out[324]));
convchan2 c_2_325 (.image, .kernel(kernels[325]), .conv_out(xor_out[325]));
convchan2 c_2_326 (.image, .kernel(kernels[326]), .conv_out(xor_out[326]));
convchan2 c_2_327 (.image, .kernel(kernels[327]), .conv_out(xor_out[327]));
convchan2 c_2_328 (.image, .kernel(kernels[328]), .conv_out(xor_out[328]));
convchan2 c_2_329 (.image, .kernel(kernels[329]), .conv_out(xor_out[329]));
convchan2 c_2_330 (.image, .kernel(kernels[330]), .conv_out(xor_out[330]));
convchan2 c_2_331 (.image, .kernel(kernels[331]), .conv_out(xor_out[331]));
convchan2 c_2_332 (.image, .kernel(kernels[332]), .conv_out(xor_out[332]));
convchan2 c_2_333 (.image, .kernel(kernels[333]), .conv_out(xor_out[333]));
convchan2 c_2_334 (.image, .kernel(kernels[334]), .conv_out(xor_out[334]));
convchan2 c_2_335 (.image, .kernel(kernels[335]), .conv_out(xor_out[335]));
convchan2 c_2_336 (.image, .kernel(kernels[336]), .conv_out(xor_out[336]));
convchan2 c_2_337 (.image, .kernel(kernels[337]), .conv_out(xor_out[337]));
convchan2 c_2_338 (.image, .kernel(kernels[338]), .conv_out(xor_out[338]));
convchan2 c_2_339 (.image, .kernel(kernels[339]), .conv_out(xor_out[339]));
convchan2 c_2_340 (.image, .kernel(kernels[340]), .conv_out(xor_out[340]));
convchan2 c_2_341 (.image, .kernel(kernels[341]), .conv_out(xor_out[341]));
convchan2 c_2_342 (.image, .kernel(kernels[342]), .conv_out(xor_out[342]));
convchan2 c_2_343 (.image, .kernel(kernels[343]), .conv_out(xor_out[343]));
convchan2 c_2_344 (.image, .kernel(kernels[344]), .conv_out(xor_out[344]));
convchan2 c_2_345 (.image, .kernel(kernels[345]), .conv_out(xor_out[345]));
convchan2 c_2_346 (.image, .kernel(kernels[346]), .conv_out(xor_out[346]));
convchan2 c_2_347 (.image, .kernel(kernels[347]), .conv_out(xor_out[347]));
convchan2 c_2_348 (.image, .kernel(kernels[348]), .conv_out(xor_out[348]));
convchan2 c_2_349 (.image, .kernel(kernels[349]), .conv_out(xor_out[349]));
convchan2 c_2_350 (.image, .kernel(kernels[350]), .conv_out(xor_out[350]));
convchan2 c_2_351 (.image, .kernel(kernels[351]), .conv_out(xor_out[351]));
convchan2 c_2_352 (.image, .kernel(kernels[352]), .conv_out(xor_out[352]));
convchan2 c_2_353 (.image, .kernel(kernels[353]), .conv_out(xor_out[353]));
convchan2 c_2_354 (.image, .kernel(kernels[354]), .conv_out(xor_out[354]));
convchan2 c_2_355 (.image, .kernel(kernels[355]), .conv_out(xor_out[355]));
convchan2 c_2_356 (.image, .kernel(kernels[356]), .conv_out(xor_out[356]));
convchan2 c_2_357 (.image, .kernel(kernels[357]), .conv_out(xor_out[357]));
convchan2 c_2_358 (.image, .kernel(kernels[358]), .conv_out(xor_out[358]));
convchan2 c_2_359 (.image, .kernel(kernels[359]), .conv_out(xor_out[359]));
convchan2 c_2_360 (.image, .kernel(kernels[360]), .conv_out(xor_out[360]));
convchan2 c_2_361 (.image, .kernel(kernels[361]), .conv_out(xor_out[361]));
convchan2 c_2_362 (.image, .kernel(kernels[362]), .conv_out(xor_out[362]));
convchan2 c_2_363 (.image, .kernel(kernels[363]), .conv_out(xor_out[363]));
convchan2 c_2_364 (.image, .kernel(kernels[364]), .conv_out(xor_out[364]));
convchan2 c_2_365 (.image, .kernel(kernels[365]), .conv_out(xor_out[365]));
convchan2 c_2_366 (.image, .kernel(kernels[366]), .conv_out(xor_out[366]));
convchan2 c_2_367 (.image, .kernel(kernels[367]), .conv_out(xor_out[367]));
convchan2 c_2_368 (.image, .kernel(kernels[368]), .conv_out(xor_out[368]));
convchan2 c_2_369 (.image, .kernel(kernels[369]), .conv_out(xor_out[369]));
convchan2 c_2_370 (.image, .kernel(kernels[370]), .conv_out(xor_out[370]));
convchan2 c_2_371 (.image, .kernel(kernels[371]), .conv_out(xor_out[371]));
convchan2 c_2_372 (.image, .kernel(kernels[372]), .conv_out(xor_out[372]));
convchan2 c_2_373 (.image, .kernel(kernels[373]), .conv_out(xor_out[373]));
convchan2 c_2_374 (.image, .kernel(kernels[374]), .conv_out(xor_out[374]));
convchan2 c_2_375 (.image, .kernel(kernels[375]), .conv_out(xor_out[375]));
convchan2 c_2_376 (.image, .kernel(kernels[376]), .conv_out(xor_out[376]));
convchan2 c_2_377 (.image, .kernel(kernels[377]), .conv_out(xor_out[377]));
convchan2 c_2_378 (.image, .kernel(kernels[378]), .conv_out(xor_out[378]));
convchan2 c_2_379 (.image, .kernel(kernels[379]), .conv_out(xor_out[379]));
convchan2 c_2_380 (.image, .kernel(kernels[380]), .conv_out(xor_out[380]));
convchan2 c_2_381 (.image, .kernel(kernels[381]), .conv_out(xor_out[381]));
convchan2 c_2_382 (.image, .kernel(kernels[382]), .conv_out(xor_out[382]));
convchan2 c_2_383 (.image, .kernel(kernels[383]), .conv_out(xor_out[383]));
convchan2 c_2_384 (.image, .kernel(kernels[384]), .conv_out(xor_out[384]));
convchan2 c_2_385 (.image, .kernel(kernels[385]), .conv_out(xor_out[385]));
convchan2 c_2_386 (.image, .kernel(kernels[386]), .conv_out(xor_out[386]));
convchan2 c_2_387 (.image, .kernel(kernels[387]), .conv_out(xor_out[387]));
convchan2 c_2_388 (.image, .kernel(kernels[388]), .conv_out(xor_out[388]));
convchan2 c_2_389 (.image, .kernel(kernels[389]), .conv_out(xor_out[389]));
convchan2 c_2_390 (.image, .kernel(kernels[390]), .conv_out(xor_out[390]));
convchan2 c_2_391 (.image, .kernel(kernels[391]), .conv_out(xor_out[391]));
convchan2 c_2_392 (.image, .kernel(kernels[392]), .conv_out(xor_out[392]));
convchan2 c_2_393 (.image, .kernel(kernels[393]), .conv_out(xor_out[393]));
convchan2 c_2_394 (.image, .kernel(kernels[394]), .conv_out(xor_out[394]));
convchan2 c_2_395 (.image, .kernel(kernels[395]), .conv_out(xor_out[395]));
convchan2 c_2_396 (.image, .kernel(kernels[396]), .conv_out(xor_out[396]));
convchan2 c_2_397 (.image, .kernel(kernels[397]), .conv_out(xor_out[397]));
convchan2 c_2_398 (.image, .kernel(kernels[398]), .conv_out(xor_out[398]));
convchan2 c_2_399 (.image, .kernel(kernels[399]), .conv_out(xor_out[399]));
convchan2 c_2_400 (.image, .kernel(kernels[400]), .conv_out(xor_out[400]));
convchan2 c_2_401 (.image, .kernel(kernels[401]), .conv_out(xor_out[401]));
convchan2 c_2_402 (.image, .kernel(kernels[402]), .conv_out(xor_out[402]));
convchan2 c_2_403 (.image, .kernel(kernels[403]), .conv_out(xor_out[403]));
convchan2 c_2_404 (.image, .kernel(kernels[404]), .conv_out(xor_out[404]));
convchan2 c_2_405 (.image, .kernel(kernels[405]), .conv_out(xor_out[405]));
convchan2 c_2_406 (.image, .kernel(kernels[406]), .conv_out(xor_out[406]));
convchan2 c_2_407 (.image, .kernel(kernels[407]), .conv_out(xor_out[407]));
convchan2 c_2_408 (.image, .kernel(kernels[408]), .conv_out(xor_out[408]));
convchan2 c_2_409 (.image, .kernel(kernels[409]), .conv_out(xor_out[409]));
convchan2 c_2_410 (.image, .kernel(kernels[410]), .conv_out(xor_out[410]));
convchan2 c_2_411 (.image, .kernel(kernels[411]), .conv_out(xor_out[411]));
convchan2 c_2_412 (.image, .kernel(kernels[412]), .conv_out(xor_out[412]));
convchan2 c_2_413 (.image, .kernel(kernels[413]), .conv_out(xor_out[413]));
convchan2 c_2_414 (.image, .kernel(kernels[414]), .conv_out(xor_out[414]));
convchan2 c_2_415 (.image, .kernel(kernels[415]), .conv_out(xor_out[415]));
convchan2 c_2_416 (.image, .kernel(kernels[416]), .conv_out(xor_out[416]));
convchan2 c_2_417 (.image, .kernel(kernels[417]), .conv_out(xor_out[417]));
convchan2 c_2_418 (.image, .kernel(kernels[418]), .conv_out(xor_out[418]));
convchan2 c_2_419 (.image, .kernel(kernels[419]), .conv_out(xor_out[419]));
convchan2 c_2_420 (.image, .kernel(kernels[420]), .conv_out(xor_out[420]));
convchan2 c_2_421 (.image, .kernel(kernels[421]), .conv_out(xor_out[421]));
convchan2 c_2_422 (.image, .kernel(kernels[422]), .conv_out(xor_out[422]));
convchan2 c_2_423 (.image, .kernel(kernels[423]), .conv_out(xor_out[423]));
convchan2 c_2_424 (.image, .kernel(kernels[424]), .conv_out(xor_out[424]));
convchan2 c_2_425 (.image, .kernel(kernels[425]), .conv_out(xor_out[425]));
convchan2 c_2_426 (.image, .kernel(kernels[426]), .conv_out(xor_out[426]));
convchan2 c_2_427 (.image, .kernel(kernels[427]), .conv_out(xor_out[427]));
convchan2 c_2_428 (.image, .kernel(kernels[428]), .conv_out(xor_out[428]));
convchan2 c_2_429 (.image, .kernel(kernels[429]), .conv_out(xor_out[429]));
convchan2 c_2_430 (.image, .kernel(kernels[430]), .conv_out(xor_out[430]));
convchan2 c_2_431 (.image, .kernel(kernels[431]), .conv_out(xor_out[431]));
convchan2 c_2_432 (.image, .kernel(kernels[432]), .conv_out(xor_out[432]));
convchan2 c_2_433 (.image, .kernel(kernels[433]), .conv_out(xor_out[433]));
convchan2 c_2_434 (.image, .kernel(kernels[434]), .conv_out(xor_out[434]));
convchan2 c_2_435 (.image, .kernel(kernels[435]), .conv_out(xor_out[435]));
convchan2 c_2_436 (.image, .kernel(kernels[436]), .conv_out(xor_out[436]));
convchan2 c_2_437 (.image, .kernel(kernels[437]), .conv_out(xor_out[437]));
convchan2 c_2_438 (.image, .kernel(kernels[438]), .conv_out(xor_out[438]));
convchan2 c_2_439 (.image, .kernel(kernels[439]), .conv_out(xor_out[439]));
convchan2 c_2_440 (.image, .kernel(kernels[440]), .conv_out(xor_out[440]));
convchan2 c_2_441 (.image, .kernel(kernels[441]), .conv_out(xor_out[441]));
convchan2 c_2_442 (.image, .kernel(kernels[442]), .conv_out(xor_out[442]));
convchan2 c_2_443 (.image, .kernel(kernels[443]), .conv_out(xor_out[443]));
convchan2 c_2_444 (.image, .kernel(kernels[444]), .conv_out(xor_out[444]));
convchan2 c_2_445 (.image, .kernel(kernels[445]), .conv_out(xor_out[445]));
convchan2 c_2_446 (.image, .kernel(kernels[446]), .conv_out(xor_out[446]));
convchan2 c_2_447 (.image, .kernel(kernels[447]), .conv_out(xor_out[447]));
convchan2 c_2_448 (.image, .kernel(kernels[448]), .conv_out(xor_out[448]));
convchan2 c_2_449 (.image, .kernel(kernels[449]), .conv_out(xor_out[449]));
convchan2 c_2_450 (.image, .kernel(kernels[450]), .conv_out(xor_out[450]));
convchan2 c_2_451 (.image, .kernel(kernels[451]), .conv_out(xor_out[451]));
convchan2 c_2_452 (.image, .kernel(kernels[452]), .conv_out(xor_out[452]));
convchan2 c_2_453 (.image, .kernel(kernels[453]), .conv_out(xor_out[453]));
convchan2 c_2_454 (.image, .kernel(kernels[454]), .conv_out(xor_out[454]));
convchan2 c_2_455 (.image, .kernel(kernels[455]), .conv_out(xor_out[455]));
convchan2 c_2_456 (.image, .kernel(kernels[456]), .conv_out(xor_out[456]));
convchan2 c_2_457 (.image, .kernel(kernels[457]), .conv_out(xor_out[457]));
convchan2 c_2_458 (.image, .kernel(kernels[458]), .conv_out(xor_out[458]));
convchan2 c_2_459 (.image, .kernel(kernels[459]), .conv_out(xor_out[459]));
convchan2 c_2_460 (.image, .kernel(kernels[460]), .conv_out(xor_out[460]));
convchan2 c_2_461 (.image, .kernel(kernels[461]), .conv_out(xor_out[461]));
convchan2 c_2_462 (.image, .kernel(kernels[462]), .conv_out(xor_out[462]));
convchan2 c_2_463 (.image, .kernel(kernels[463]), .conv_out(xor_out[463]));
convchan2 c_2_464 (.image, .kernel(kernels[464]), .conv_out(xor_out[464]));
convchan2 c_2_465 (.image, .kernel(kernels[465]), .conv_out(xor_out[465]));
convchan2 c_2_466 (.image, .kernel(kernels[466]), .conv_out(xor_out[466]));
convchan2 c_2_467 (.image, .kernel(kernels[467]), .conv_out(xor_out[467]));
convchan2 c_2_468 (.image, .kernel(kernels[468]), .conv_out(xor_out[468]));
convchan2 c_2_469 (.image, .kernel(kernels[469]), .conv_out(xor_out[469]));
convchan2 c_2_470 (.image, .kernel(kernels[470]), .conv_out(xor_out[470]));
convchan2 c_2_471 (.image, .kernel(kernels[471]), .conv_out(xor_out[471]));
convchan2 c_2_472 (.image, .kernel(kernels[472]), .conv_out(xor_out[472]));
convchan2 c_2_473 (.image, .kernel(kernels[473]), .conv_out(xor_out[473]));
convchan2 c_2_474 (.image, .kernel(kernels[474]), .conv_out(xor_out[474]));
convchan2 c_2_475 (.image, .kernel(kernels[475]), .conv_out(xor_out[475]));
convchan2 c_2_476 (.image, .kernel(kernels[476]), .conv_out(xor_out[476]));
convchan2 c_2_477 (.image, .kernel(kernels[477]), .conv_out(xor_out[477]));
convchan2 c_2_478 (.image, .kernel(kernels[478]), .conv_out(xor_out[478]));
convchan2 c_2_479 (.image, .kernel(kernels[479]), .conv_out(xor_out[479]));
convchan2 c_2_480 (.image, .kernel(kernels[480]), .conv_out(xor_out[480]));
convchan2 c_2_481 (.image, .kernel(kernels[481]), .conv_out(xor_out[481]));
convchan2 c_2_482 (.image, .kernel(kernels[482]), .conv_out(xor_out[482]));
convchan2 c_2_483 (.image, .kernel(kernels[483]), .conv_out(xor_out[483]));
convchan2 c_2_484 (.image, .kernel(kernels[484]), .conv_out(xor_out[484]));
convchan2 c_2_485 (.image, .kernel(kernels[485]), .conv_out(xor_out[485]));
convchan2 c_2_486 (.image, .kernel(kernels[486]), .conv_out(xor_out[486]));
convchan2 c_2_487 (.image, .kernel(kernels[487]), .conv_out(xor_out[487]));
convchan2 c_2_488 (.image, .kernel(kernels[488]), .conv_out(xor_out[488]));
convchan2 c_2_489 (.image, .kernel(kernels[489]), .conv_out(xor_out[489]));
convchan2 c_2_490 (.image, .kernel(kernels[490]), .conv_out(xor_out[490]));
convchan2 c_2_491 (.image, .kernel(kernels[491]), .conv_out(xor_out[491]));
convchan2 c_2_492 (.image, .kernel(kernels[492]), .conv_out(xor_out[492]));
convchan2 c_2_493 (.image, .kernel(kernels[493]), .conv_out(xor_out[493]));
convchan2 c_2_494 (.image, .kernel(kernels[494]), .conv_out(xor_out[494]));
convchan2 c_2_495 (.image, .kernel(kernels[495]), .conv_out(xor_out[495]));
convchan2 c_2_496 (.image, .kernel(kernels[496]), .conv_out(xor_out[496]));
convchan2 c_2_497 (.image, .kernel(kernels[497]), .conv_out(xor_out[497]));
convchan2 c_2_498 (.image, .kernel(kernels[498]), .conv_out(xor_out[498]));
convchan2 c_2_499 (.image, .kernel(kernels[499]), .conv_out(xor_out[499]));
convchan2 c_2_500 (.image, .kernel(kernels[500]), .conv_out(xor_out[500]));
convchan2 c_2_501 (.image, .kernel(kernels[501]), .conv_out(xor_out[501]));
convchan2 c_2_502 (.image, .kernel(kernels[502]), .conv_out(xor_out[502]));
convchan2 c_2_503 (.image, .kernel(kernels[503]), .conv_out(xor_out[503]));
convchan2 c_2_504 (.image, .kernel(kernels[504]), .conv_out(xor_out[504]));
convchan2 c_2_505 (.image, .kernel(kernels[505]), .conv_out(xor_out[505]));
convchan2 c_2_506 (.image, .kernel(kernels[506]), .conv_out(xor_out[506]));
convchan2 c_2_507 (.image, .kernel(kernels[507]), .conv_out(xor_out[507]));
convchan2 c_2_508 (.image, .kernel(kernels[508]), .conv_out(xor_out[508]));
convchan2 c_2_509 (.image, .kernel(kernels[509]), .conv_out(xor_out[509]));
convchan2 c_2_510 (.image, .kernel(kernels[510]), .conv_out(xor_out[510]));
convchan2 c_2_511 (.image, .kernel(kernels[511]), .conv_out(xor_out[511]));
convchan2 c_2_512 (.image, .kernel(kernels[512]), .conv_out(xor_out[512]));
convchan2 c_2_513 (.image, .kernel(kernels[513]), .conv_out(xor_out[513]));
convchan2 c_2_514 (.image, .kernel(kernels[514]), .conv_out(xor_out[514]));
convchan2 c_2_515 (.image, .kernel(kernels[515]), .conv_out(xor_out[515]));
convchan2 c_2_516 (.image, .kernel(kernels[516]), .conv_out(xor_out[516]));
convchan2 c_2_517 (.image, .kernel(kernels[517]), .conv_out(xor_out[517]));
convchan2 c_2_518 (.image, .kernel(kernels[518]), .conv_out(xor_out[518]));
convchan2 c_2_519 (.image, .kernel(kernels[519]), .conv_out(xor_out[519]));
convchan2 c_2_520 (.image, .kernel(kernels[520]), .conv_out(xor_out[520]));
convchan2 c_2_521 (.image, .kernel(kernels[521]), .conv_out(xor_out[521]));
convchan2 c_2_522 (.image, .kernel(kernels[522]), .conv_out(xor_out[522]));
convchan2 c_2_523 (.image, .kernel(kernels[523]), .conv_out(xor_out[523]));
convchan2 c_2_524 (.image, .kernel(kernels[524]), .conv_out(xor_out[524]));
convchan2 c_2_525 (.image, .kernel(kernels[525]), .conv_out(xor_out[525]));
convchan2 c_2_526 (.image, .kernel(kernels[526]), .conv_out(xor_out[526]));
convchan2 c_2_527 (.image, .kernel(kernels[527]), .conv_out(xor_out[527]));
convchan2 c_2_528 (.image, .kernel(kernels[528]), .conv_out(xor_out[528]));
convchan2 c_2_529 (.image, .kernel(kernels[529]), .conv_out(xor_out[529]));
convchan2 c_2_530 (.image, .kernel(kernels[530]), .conv_out(xor_out[530]));
convchan2 c_2_531 (.image, .kernel(kernels[531]), .conv_out(xor_out[531]));
convchan2 c_2_532 (.image, .kernel(kernels[532]), .conv_out(xor_out[532]));
convchan2 c_2_533 (.image, .kernel(kernels[533]), .conv_out(xor_out[533]));
convchan2 c_2_534 (.image, .kernel(kernels[534]), .conv_out(xor_out[534]));
convchan2 c_2_535 (.image, .kernel(kernels[535]), .conv_out(xor_out[535]));
convchan2 c_2_536 (.image, .kernel(kernels[536]), .conv_out(xor_out[536]));
convchan2 c_2_537 (.image, .kernel(kernels[537]), .conv_out(xor_out[537]));
convchan2 c_2_538 (.image, .kernel(kernels[538]), .conv_out(xor_out[538]));
convchan2 c_2_539 (.image, .kernel(kernels[539]), .conv_out(xor_out[539]));
convchan2 c_2_540 (.image, .kernel(kernels[540]), .conv_out(xor_out[540]));
convchan2 c_2_541 (.image, .kernel(kernels[541]), .conv_out(xor_out[541]));
convchan2 c_2_542 (.image, .kernel(kernels[542]), .conv_out(xor_out[542]));
convchan2 c_2_543 (.image, .kernel(kernels[543]), .conv_out(xor_out[543]));
convchan2 c_2_544 (.image, .kernel(kernels[544]), .conv_out(xor_out[544]));
convchan2 c_2_545 (.image, .kernel(kernels[545]), .conv_out(xor_out[545]));
convchan2 c_2_546 (.image, .kernel(kernels[546]), .conv_out(xor_out[546]));
convchan2 c_2_547 (.image, .kernel(kernels[547]), .conv_out(xor_out[547]));
convchan2 c_2_548 (.image, .kernel(kernels[548]), .conv_out(xor_out[548]));
convchan2 c_2_549 (.image, .kernel(kernels[549]), .conv_out(xor_out[549]));
convchan2 c_2_550 (.image, .kernel(kernels[550]), .conv_out(xor_out[550]));
convchan2 c_2_551 (.image, .kernel(kernels[551]), .conv_out(xor_out[551]));
convchan2 c_2_552 (.image, .kernel(kernels[552]), .conv_out(xor_out[552]));
convchan2 c_2_553 (.image, .kernel(kernels[553]), .conv_out(xor_out[553]));
convchan2 c_2_554 (.image, .kernel(kernels[554]), .conv_out(xor_out[554]));
convchan2 c_2_555 (.image, .kernel(kernels[555]), .conv_out(xor_out[555]));
convchan2 c_2_556 (.image, .kernel(kernels[556]), .conv_out(xor_out[556]));
convchan2 c_2_557 (.image, .kernel(kernels[557]), .conv_out(xor_out[557]));
convchan2 c_2_558 (.image, .kernel(kernels[558]), .conv_out(xor_out[558]));
convchan2 c_2_559 (.image, .kernel(kernels[559]), .conv_out(xor_out[559]));
convchan2 c_2_560 (.image, .kernel(kernels[560]), .conv_out(xor_out[560]));
convchan2 c_2_561 (.image, .kernel(kernels[561]), .conv_out(xor_out[561]));
convchan2 c_2_562 (.image, .kernel(kernels[562]), .conv_out(xor_out[562]));
convchan2 c_2_563 (.image, .kernel(kernels[563]), .conv_out(xor_out[563]));
convchan2 c_2_564 (.image, .kernel(kernels[564]), .conv_out(xor_out[564]));
convchan2 c_2_565 (.image, .kernel(kernels[565]), .conv_out(xor_out[565]));
convchan2 c_2_566 (.image, .kernel(kernels[566]), .conv_out(xor_out[566]));
convchan2 c_2_567 (.image, .kernel(kernels[567]), .conv_out(xor_out[567]));
convchan2 c_2_568 (.image, .kernel(kernels[568]), .conv_out(xor_out[568]));
convchan2 c_2_569 (.image, .kernel(kernels[569]), .conv_out(xor_out[569]));
convchan2 c_2_570 (.image, .kernel(kernels[570]), .conv_out(xor_out[570]));
convchan2 c_2_571 (.image, .kernel(kernels[571]), .conv_out(xor_out[571]));
convchan2 c_2_572 (.image, .kernel(kernels[572]), .conv_out(xor_out[572]));
convchan2 c_2_573 (.image, .kernel(kernels[573]), .conv_out(xor_out[573]));
convchan2 c_2_574 (.image, .kernel(kernels[574]), .conv_out(xor_out[574]));
convchan2 c_2_575 (.image, .kernel(kernels[575]), .conv_out(xor_out[575]));
convchan2 c_2_576 (.image, .kernel(kernels[576]), .conv_out(xor_out[576]));
convchan2 c_2_577 (.image, .kernel(kernels[577]), .conv_out(xor_out[577]));
convchan2 c_2_578 (.image, .kernel(kernels[578]), .conv_out(xor_out[578]));
convchan2 c_2_579 (.image, .kernel(kernels[579]), .conv_out(xor_out[579]));
convchan2 c_2_580 (.image, .kernel(kernels[580]), .conv_out(xor_out[580]));
convchan2 c_2_581 (.image, .kernel(kernels[581]), .conv_out(xor_out[581]));
convchan2 c_2_582 (.image, .kernel(kernels[582]), .conv_out(xor_out[582]));
convchan2 c_2_583 (.image, .kernel(kernels[583]), .conv_out(xor_out[583]));
convchan2 c_2_584 (.image, .kernel(kernels[584]), .conv_out(xor_out[584]));
convchan2 c_2_585 (.image, .kernel(kernels[585]), .conv_out(xor_out[585]));
convchan2 c_2_586 (.image, .kernel(kernels[586]), .conv_out(xor_out[586]));
convchan2 c_2_587 (.image, .kernel(kernels[587]), .conv_out(xor_out[587]));
convchan2 c_2_588 (.image, .kernel(kernels[588]), .conv_out(xor_out[588]));
convchan2 c_2_589 (.image, .kernel(kernels[589]), .conv_out(xor_out[589]));
convchan2 c_2_590 (.image, .kernel(kernels[590]), .conv_out(xor_out[590]));
convchan2 c_2_591 (.image, .kernel(kernels[591]), .conv_out(xor_out[591]));
convchan2 c_2_592 (.image, .kernel(kernels[592]), .conv_out(xor_out[592]));
convchan2 c_2_593 (.image, .kernel(kernels[593]), .conv_out(xor_out[593]));
convchan2 c_2_594 (.image, .kernel(kernels[594]), .conv_out(xor_out[594]));
convchan2 c_2_595 (.image, .kernel(kernels[595]), .conv_out(xor_out[595]));
convchan2 c_2_596 (.image, .kernel(kernels[596]), .conv_out(xor_out[596]));
convchan2 c_2_597 (.image, .kernel(kernels[597]), .conv_out(xor_out[597]));
convchan2 c_2_598 (.image, .kernel(kernels[598]), .conv_out(xor_out[598]));
convchan2 c_2_599 (.image, .kernel(kernels[599]), .conv_out(xor_out[599]));
convchan2 c_2_600 (.image, .kernel(kernels[600]), .conv_out(xor_out[600]));
convchan2 c_2_601 (.image, .kernel(kernels[601]), .conv_out(xor_out[601]));
convchan2 c_2_602 (.image, .kernel(kernels[602]), .conv_out(xor_out[602]));
convchan2 c_2_603 (.image, .kernel(kernels[603]), .conv_out(xor_out[603]));
convchan2 c_2_604 (.image, .kernel(kernels[604]), .conv_out(xor_out[604]));
convchan2 c_2_605 (.image, .kernel(kernels[605]), .conv_out(xor_out[605]));
convchan2 c_2_606 (.image, .kernel(kernels[606]), .conv_out(xor_out[606]));
convchan2 c_2_607 (.image, .kernel(kernels[607]), .conv_out(xor_out[607]));
convchan2 c_2_608 (.image, .kernel(kernels[608]), .conv_out(xor_out[608]));
convchan2 c_2_609 (.image, .kernel(kernels[609]), .conv_out(xor_out[609]));
convchan2 c_2_610 (.image, .kernel(kernels[610]), .conv_out(xor_out[610]));
convchan2 c_2_611 (.image, .kernel(kernels[611]), .conv_out(xor_out[611]));
convchan2 c_2_612 (.image, .kernel(kernels[612]), .conv_out(xor_out[612]));
convchan2 c_2_613 (.image, .kernel(kernels[613]), .conv_out(xor_out[613]));
convchan2 c_2_614 (.image, .kernel(kernels[614]), .conv_out(xor_out[614]));
convchan2 c_2_615 (.image, .kernel(kernels[615]), .conv_out(xor_out[615]));
convchan2 c_2_616 (.image, .kernel(kernels[616]), .conv_out(xor_out[616]));
convchan2 c_2_617 (.image, .kernel(kernels[617]), .conv_out(xor_out[617]));
convchan2 c_2_618 (.image, .kernel(kernels[618]), .conv_out(xor_out[618]));
convchan2 c_2_619 (.image, .kernel(kernels[619]), .conv_out(xor_out[619]));
convchan2 c_2_620 (.image, .kernel(kernels[620]), .conv_out(xor_out[620]));
convchan2 c_2_621 (.image, .kernel(kernels[621]), .conv_out(xor_out[621]));
convchan2 c_2_622 (.image, .kernel(kernels[622]), .conv_out(xor_out[622]));
convchan2 c_2_623 (.image, .kernel(kernels[623]), .conv_out(xor_out[623]));
convchan2 c_2_624 (.image, .kernel(kernels[624]), .conv_out(xor_out[624]));
convchan2 c_2_625 (.image, .kernel(kernels[625]), .conv_out(xor_out[625]));
convchan2 c_2_626 (.image, .kernel(kernels[626]), .conv_out(xor_out[626]));
convchan2 c_2_627 (.image, .kernel(kernels[627]), .conv_out(xor_out[627]));
convchan2 c_2_628 (.image, .kernel(kernels[628]), .conv_out(xor_out[628]));
convchan2 c_2_629 (.image, .kernel(kernels[629]), .conv_out(xor_out[629]));
convchan2 c_2_630 (.image, .kernel(kernels[630]), .conv_out(xor_out[630]));
convchan2 c_2_631 (.image, .kernel(kernels[631]), .conv_out(xor_out[631]));
convchan2 c_2_632 (.image, .kernel(kernels[632]), .conv_out(xor_out[632]));
convchan2 c_2_633 (.image, .kernel(kernels[633]), .conv_out(xor_out[633]));
convchan2 c_2_634 (.image, .kernel(kernels[634]), .conv_out(xor_out[634]));
convchan2 c_2_635 (.image, .kernel(kernels[635]), .conv_out(xor_out[635]));
convchan2 c_2_636 (.image, .kernel(kernels[636]), .conv_out(xor_out[636]));
convchan2 c_2_637 (.image, .kernel(kernels[637]), .conv_out(xor_out[637]));
convchan2 c_2_638 (.image, .kernel(kernels[638]), .conv_out(xor_out[638]));
convchan2 c_2_639 (.image, .kernel(kernels[639]), .conv_out(xor_out[639]));
convchan2 c_2_640 (.image, .kernel(kernels[640]), .conv_out(xor_out[640]));
convchan2 c_2_641 (.image, .kernel(kernels[641]), .conv_out(xor_out[641]));
convchan2 c_2_642 (.image, .kernel(kernels[642]), .conv_out(xor_out[642]));
convchan2 c_2_643 (.image, .kernel(kernels[643]), .conv_out(xor_out[643]));
convchan2 c_2_644 (.image, .kernel(kernels[644]), .conv_out(xor_out[644]));
convchan2 c_2_645 (.image, .kernel(kernels[645]), .conv_out(xor_out[645]));
convchan2 c_2_646 (.image, .kernel(kernels[646]), .conv_out(xor_out[646]));
convchan2 c_2_647 (.image, .kernel(kernels[647]), .conv_out(xor_out[647]));
convchan2 c_2_648 (.image, .kernel(kernels[648]), .conv_out(xor_out[648]));
convchan2 c_2_649 (.image, .kernel(kernels[649]), .conv_out(xor_out[649]));
convchan2 c_2_650 (.image, .kernel(kernels[650]), .conv_out(xor_out[650]));
convchan2 c_2_651 (.image, .kernel(kernels[651]), .conv_out(xor_out[651]));
convchan2 c_2_652 (.image, .kernel(kernels[652]), .conv_out(xor_out[652]));
convchan2 c_2_653 (.image, .kernel(kernels[653]), .conv_out(xor_out[653]));
convchan2 c_2_654 (.image, .kernel(kernels[654]), .conv_out(xor_out[654]));
convchan2 c_2_655 (.image, .kernel(kernels[655]), .conv_out(xor_out[655]));
convchan2 c_2_656 (.image, .kernel(kernels[656]), .conv_out(xor_out[656]));
convchan2 c_2_657 (.image, .kernel(kernels[657]), .conv_out(xor_out[657]));
convchan2 c_2_658 (.image, .kernel(kernels[658]), .conv_out(xor_out[658]));
convchan2 c_2_659 (.image, .kernel(kernels[659]), .conv_out(xor_out[659]));
convchan2 c_2_660 (.image, .kernel(kernels[660]), .conv_out(xor_out[660]));
convchan2 c_2_661 (.image, .kernel(kernels[661]), .conv_out(xor_out[661]));
convchan2 c_2_662 (.image, .kernel(kernels[662]), .conv_out(xor_out[662]));
convchan2 c_2_663 (.image, .kernel(kernels[663]), .conv_out(xor_out[663]));
convchan2 c_2_664 (.image, .kernel(kernels[664]), .conv_out(xor_out[664]));
convchan2 c_2_665 (.image, .kernel(kernels[665]), .conv_out(xor_out[665]));
convchan2 c_2_666 (.image, .kernel(kernels[666]), .conv_out(xor_out[666]));
convchan2 c_2_667 (.image, .kernel(kernels[667]), .conv_out(xor_out[667]));
convchan2 c_2_668 (.image, .kernel(kernels[668]), .conv_out(xor_out[668]));
convchan2 c_2_669 (.image, .kernel(kernels[669]), .conv_out(xor_out[669]));
convchan2 c_2_670 (.image, .kernel(kernels[670]), .conv_out(xor_out[670]));
convchan2 c_2_671 (.image, .kernel(kernels[671]), .conv_out(xor_out[671]));
convchan2 c_2_672 (.image, .kernel(kernels[672]), .conv_out(xor_out[672]));
convchan2 c_2_673 (.image, .kernel(kernels[673]), .conv_out(xor_out[673]));
convchan2 c_2_674 (.image, .kernel(kernels[674]), .conv_out(xor_out[674]));
convchan2 c_2_675 (.image, .kernel(kernels[675]), .conv_out(xor_out[675]));
convchan2 c_2_676 (.image, .kernel(kernels[676]), .conv_out(xor_out[676]));
convchan2 c_2_677 (.image, .kernel(kernels[677]), .conv_out(xor_out[677]));
convchan2 c_2_678 (.image, .kernel(kernels[678]), .conv_out(xor_out[678]));
convchan2 c_2_679 (.image, .kernel(kernels[679]), .conv_out(xor_out[679]));
convchan2 c_2_680 (.image, .kernel(kernels[680]), .conv_out(xor_out[680]));
convchan2 c_2_681 (.image, .kernel(kernels[681]), .conv_out(xor_out[681]));
convchan2 c_2_682 (.image, .kernel(kernels[682]), .conv_out(xor_out[682]));
convchan2 c_2_683 (.image, .kernel(kernels[683]), .conv_out(xor_out[683]));
convchan2 c_2_684 (.image, .kernel(kernels[684]), .conv_out(xor_out[684]));
convchan2 c_2_685 (.image, .kernel(kernels[685]), .conv_out(xor_out[685]));
convchan2 c_2_686 (.image, .kernel(kernels[686]), .conv_out(xor_out[686]));
convchan2 c_2_687 (.image, .kernel(kernels[687]), .conv_out(xor_out[687]));
convchan2 c_2_688 (.image, .kernel(kernels[688]), .conv_out(xor_out[688]));
convchan2 c_2_689 (.image, .kernel(kernels[689]), .conv_out(xor_out[689]));
convchan2 c_2_690 (.image, .kernel(kernels[690]), .conv_out(xor_out[690]));
convchan2 c_2_691 (.image, .kernel(kernels[691]), .conv_out(xor_out[691]));
convchan2 c_2_692 (.image, .kernel(kernels[692]), .conv_out(xor_out[692]));
convchan2 c_2_693 (.image, .kernel(kernels[693]), .conv_out(xor_out[693]));
convchan2 c_2_694 (.image, .kernel(kernels[694]), .conv_out(xor_out[694]));
convchan2 c_2_695 (.image, .kernel(kernels[695]), .conv_out(xor_out[695]));
convchan2 c_2_696 (.image, .kernel(kernels[696]), .conv_out(xor_out[696]));
convchan2 c_2_697 (.image, .kernel(kernels[697]), .conv_out(xor_out[697]));
convchan2 c_2_698 (.image, .kernel(kernels[698]), .conv_out(xor_out[698]));
convchan2 c_2_699 (.image, .kernel(kernels[699]), .conv_out(xor_out[699]));
convchan2 c_2_700 (.image, .kernel(kernels[700]), .conv_out(xor_out[700]));
convchan2 c_2_701 (.image, .kernel(kernels[701]), .conv_out(xor_out[701]));
convchan2 c_2_702 (.image, .kernel(kernels[702]), .conv_out(xor_out[702]));
convchan2 c_2_703 (.image, .kernel(kernels[703]), .conv_out(xor_out[703]));
convchan2 c_2_704 (.image, .kernel(kernels[704]), .conv_out(xor_out[704]));
convchan2 c_2_705 (.image, .kernel(kernels[705]), .conv_out(xor_out[705]));
convchan2 c_2_706 (.image, .kernel(kernels[706]), .conv_out(xor_out[706]));
convchan2 c_2_707 (.image, .kernel(kernels[707]), .conv_out(xor_out[707]));
convchan2 c_2_708 (.image, .kernel(kernels[708]), .conv_out(xor_out[708]));
convchan2 c_2_709 (.image, .kernel(kernels[709]), .conv_out(xor_out[709]));
convchan2 c_2_710 (.image, .kernel(kernels[710]), .conv_out(xor_out[710]));
convchan2 c_2_711 (.image, .kernel(kernels[711]), .conv_out(xor_out[711]));
convchan2 c_2_712 (.image, .kernel(kernels[712]), .conv_out(xor_out[712]));
convchan2 c_2_713 (.image, .kernel(kernels[713]), .conv_out(xor_out[713]));
convchan2 c_2_714 (.image, .kernel(kernels[714]), .conv_out(xor_out[714]));
convchan2 c_2_715 (.image, .kernel(kernels[715]), .conv_out(xor_out[715]));
convchan2 c_2_716 (.image, .kernel(kernels[716]), .conv_out(xor_out[716]));
convchan2 c_2_717 (.image, .kernel(kernels[717]), .conv_out(xor_out[717]));
convchan2 c_2_718 (.image, .kernel(kernels[718]), .conv_out(xor_out[718]));
convchan2 c_2_719 (.image, .kernel(kernels[719]), .conv_out(xor_out[719]));
convchan2 c_2_720 (.image, .kernel(kernels[720]), .conv_out(xor_out[720]));
convchan2 c_2_721 (.image, .kernel(kernels[721]), .conv_out(xor_out[721]));
convchan2 c_2_722 (.image, .kernel(kernels[722]), .conv_out(xor_out[722]));
convchan2 c_2_723 (.image, .kernel(kernels[723]), .conv_out(xor_out[723]));
convchan2 c_2_724 (.image, .kernel(kernels[724]), .conv_out(xor_out[724]));
convchan2 c_2_725 (.image, .kernel(kernels[725]), .conv_out(xor_out[725]));
convchan2 c_2_726 (.image, .kernel(kernels[726]), .conv_out(xor_out[726]));
convchan2 c_2_727 (.image, .kernel(kernels[727]), .conv_out(xor_out[727]));
convchan2 c_2_728 (.image, .kernel(kernels[728]), .conv_out(xor_out[728]));
convchan2 c_2_729 (.image, .kernel(kernels[729]), .conv_out(xor_out[729]));
convchan2 c_2_730 (.image, .kernel(kernels[730]), .conv_out(xor_out[730]));
convchan2 c_2_731 (.image, .kernel(kernels[731]), .conv_out(xor_out[731]));
convchan2 c_2_732 (.image, .kernel(kernels[732]), .conv_out(xor_out[732]));
convchan2 c_2_733 (.image, .kernel(kernels[733]), .conv_out(xor_out[733]));
convchan2 c_2_734 (.image, .kernel(kernels[734]), .conv_out(xor_out[734]));
convchan2 c_2_735 (.image, .kernel(kernels[735]), .conv_out(xor_out[735]));
convchan2 c_2_736 (.image, .kernel(kernels[736]), .conv_out(xor_out[736]));
convchan2 c_2_737 (.image, .kernel(kernels[737]), .conv_out(xor_out[737]));
convchan2 c_2_738 (.image, .kernel(kernels[738]), .conv_out(xor_out[738]));
convchan2 c_2_739 (.image, .kernel(kernels[739]), .conv_out(xor_out[739]));
convchan2 c_2_740 (.image, .kernel(kernels[740]), .conv_out(xor_out[740]));
convchan2 c_2_741 (.image, .kernel(kernels[741]), .conv_out(xor_out[741]));
convchan2 c_2_742 (.image, .kernel(kernels[742]), .conv_out(xor_out[742]));
convchan2 c_2_743 (.image, .kernel(kernels[743]), .conv_out(xor_out[743]));
convchan2 c_2_744 (.image, .kernel(kernels[744]), .conv_out(xor_out[744]));
convchan2 c_2_745 (.image, .kernel(kernels[745]), .conv_out(xor_out[745]));
convchan2 c_2_746 (.image, .kernel(kernels[746]), .conv_out(xor_out[746]));
convchan2 c_2_747 (.image, .kernel(kernels[747]), .conv_out(xor_out[747]));
convchan2 c_2_748 (.image, .kernel(kernels[748]), .conv_out(xor_out[748]));
convchan2 c_2_749 (.image, .kernel(kernels[749]), .conv_out(xor_out[749]));
convchan2 c_2_750 (.image, .kernel(kernels[750]), .conv_out(xor_out[750]));
convchan2 c_2_751 (.image, .kernel(kernels[751]), .conv_out(xor_out[751]));
convchan2 c_2_752 (.image, .kernel(kernels[752]), .conv_out(xor_out[752]));
convchan2 c_2_753 (.image, .kernel(kernels[753]), .conv_out(xor_out[753]));
convchan2 c_2_754 (.image, .kernel(kernels[754]), .conv_out(xor_out[754]));
convchan2 c_2_755 (.image, .kernel(kernels[755]), .conv_out(xor_out[755]));
convchan2 c_2_756 (.image, .kernel(kernels[756]), .conv_out(xor_out[756]));
convchan2 c_2_757 (.image, .kernel(kernels[757]), .conv_out(xor_out[757]));
convchan2 c_2_758 (.image, .kernel(kernels[758]), .conv_out(xor_out[758]));
convchan2 c_2_759 (.image, .kernel(kernels[759]), .conv_out(xor_out[759]));
convchan2 c_2_760 (.image, .kernel(kernels[760]), .conv_out(xor_out[760]));
convchan2 c_2_761 (.image, .kernel(kernels[761]), .conv_out(xor_out[761]));
convchan2 c_2_762 (.image, .kernel(kernels[762]), .conv_out(xor_out[762]));
convchan2 c_2_763 (.image, .kernel(kernels[763]), .conv_out(xor_out[763]));
convchan2 c_2_764 (.image, .kernel(kernels[764]), .conv_out(xor_out[764]));
convchan2 c_2_765 (.image, .kernel(kernels[765]), .conv_out(xor_out[765]));
convchan2 c_2_766 (.image, .kernel(kernels[766]), .conv_out(xor_out[766]));
convchan2 c_2_767 (.image, .kernel(kernels[767]), .conv_out(xor_out[767]));
convchan2 c_2_768 (.image, .kernel(kernels[768]), .conv_out(xor_out[768]));
convchan2 c_2_769 (.image, .kernel(kernels[769]), .conv_out(xor_out[769]));
convchan2 c_2_770 (.image, .kernel(kernels[770]), .conv_out(xor_out[770]));
convchan2 c_2_771 (.image, .kernel(kernels[771]), .conv_out(xor_out[771]));
convchan2 c_2_772 (.image, .kernel(kernels[772]), .conv_out(xor_out[772]));
convchan2 c_2_773 (.image, .kernel(kernels[773]), .conv_out(xor_out[773]));
convchan2 c_2_774 (.image, .kernel(kernels[774]), .conv_out(xor_out[774]));
convchan2 c_2_775 (.image, .kernel(kernels[775]), .conv_out(xor_out[775]));
convchan2 c_2_776 (.image, .kernel(kernels[776]), .conv_out(xor_out[776]));
convchan2 c_2_777 (.image, .kernel(kernels[777]), .conv_out(xor_out[777]));
convchan2 c_2_778 (.image, .kernel(kernels[778]), .conv_out(xor_out[778]));
convchan2 c_2_779 (.image, .kernel(kernels[779]), .conv_out(xor_out[779]));
convchan2 c_2_780 (.image, .kernel(kernels[780]), .conv_out(xor_out[780]));
convchan2 c_2_781 (.image, .kernel(kernels[781]), .conv_out(xor_out[781]));
convchan2 c_2_782 (.image, .kernel(kernels[782]), .conv_out(xor_out[782]));
convchan2 c_2_783 (.image, .kernel(kernels[783]), .conv_out(xor_out[783]));
convchan2 c_2_784 (.image, .kernel(kernels[784]), .conv_out(xor_out[784]));
convchan2 c_2_785 (.image, .kernel(kernels[785]), .conv_out(xor_out[785]));
convchan2 c_2_786 (.image, .kernel(kernels[786]), .conv_out(xor_out[786]));
convchan2 c_2_787 (.image, .kernel(kernels[787]), .conv_out(xor_out[787]));
convchan2 c_2_788 (.image, .kernel(kernels[788]), .conv_out(xor_out[788]));
convchan2 c_2_789 (.image, .kernel(kernels[789]), .conv_out(xor_out[789]));
convchan2 c_2_790 (.image, .kernel(kernels[790]), .conv_out(xor_out[790]));
convchan2 c_2_791 (.image, .kernel(kernels[791]), .conv_out(xor_out[791]));
convchan2 c_2_792 (.image, .kernel(kernels[792]), .conv_out(xor_out[792]));
convchan2 c_2_793 (.image, .kernel(kernels[793]), .conv_out(xor_out[793]));
convchan2 c_2_794 (.image, .kernel(kernels[794]), .conv_out(xor_out[794]));
convchan2 c_2_795 (.image, .kernel(kernels[795]), .conv_out(xor_out[795]));
convchan2 c_2_796 (.image, .kernel(kernels[796]), .conv_out(xor_out[796]));
convchan2 c_2_797 (.image, .kernel(kernels[797]), .conv_out(xor_out[797]));
convchan2 c_2_798 (.image, .kernel(kernels[798]), .conv_out(xor_out[798]));
convchan2 c_2_799 (.image, .kernel(kernels[799]), .conv_out(xor_out[799]));
convchan2 c_2_800 (.image, .kernel(kernels[800]), .conv_out(xor_out[800]));
convchan2 c_2_801 (.image, .kernel(kernels[801]), .conv_out(xor_out[801]));
convchan2 c_2_802 (.image, .kernel(kernels[802]), .conv_out(xor_out[802]));
convchan2 c_2_803 (.image, .kernel(kernels[803]), .conv_out(xor_out[803]));
convchan2 c_2_804 (.image, .kernel(kernels[804]), .conv_out(xor_out[804]));
convchan2 c_2_805 (.image, .kernel(kernels[805]), .conv_out(xor_out[805]));
convchan2 c_2_806 (.image, .kernel(kernels[806]), .conv_out(xor_out[806]));
convchan2 c_2_807 (.image, .kernel(kernels[807]), .conv_out(xor_out[807]));
convchan2 c_2_808 (.image, .kernel(kernels[808]), .conv_out(xor_out[808]));
convchan2 c_2_809 (.image, .kernel(kernels[809]), .conv_out(xor_out[809]));
convchan2 c_2_810 (.image, .kernel(kernels[810]), .conv_out(xor_out[810]));
convchan2 c_2_811 (.image, .kernel(kernels[811]), .conv_out(xor_out[811]));
convchan2 c_2_812 (.image, .kernel(kernels[812]), .conv_out(xor_out[812]));
convchan2 c_2_813 (.image, .kernel(kernels[813]), .conv_out(xor_out[813]));
convchan2 c_2_814 (.image, .kernel(kernels[814]), .conv_out(xor_out[814]));
convchan2 c_2_815 (.image, .kernel(kernels[815]), .conv_out(xor_out[815]));
convchan2 c_2_816 (.image, .kernel(kernels[816]), .conv_out(xor_out[816]));
convchan2 c_2_817 (.image, .kernel(kernels[817]), .conv_out(xor_out[817]));
convchan2 c_2_818 (.image, .kernel(kernels[818]), .conv_out(xor_out[818]));
convchan2 c_2_819 (.image, .kernel(kernels[819]), .conv_out(xor_out[819]));
convchan2 c_2_820 (.image, .kernel(kernels[820]), .conv_out(xor_out[820]));
convchan2 c_2_821 (.image, .kernel(kernels[821]), .conv_out(xor_out[821]));
convchan2 c_2_822 (.image, .kernel(kernels[822]), .conv_out(xor_out[822]));
convchan2 c_2_823 (.image, .kernel(kernels[823]), .conv_out(xor_out[823]));
convchan2 c_2_824 (.image, .kernel(kernels[824]), .conv_out(xor_out[824]));
convchan2 c_2_825 (.image, .kernel(kernels[825]), .conv_out(xor_out[825]));
convchan2 c_2_826 (.image, .kernel(kernels[826]), .conv_out(xor_out[826]));
convchan2 c_2_827 (.image, .kernel(kernels[827]), .conv_out(xor_out[827]));
convchan2 c_2_828 (.image, .kernel(kernels[828]), .conv_out(xor_out[828]));
convchan2 c_2_829 (.image, .kernel(kernels[829]), .conv_out(xor_out[829]));
convchan2 c_2_830 (.image, .kernel(kernels[830]), .conv_out(xor_out[830]));
convchan2 c_2_831 (.image, .kernel(kernels[831]), .conv_out(xor_out[831]));
convchan2 c_2_832 (.image, .kernel(kernels[832]), .conv_out(xor_out[832]));
convchan2 c_2_833 (.image, .kernel(kernels[833]), .conv_out(xor_out[833]));
convchan2 c_2_834 (.image, .kernel(kernels[834]), .conv_out(xor_out[834]));
convchan2 c_2_835 (.image, .kernel(kernels[835]), .conv_out(xor_out[835]));
convchan2 c_2_836 (.image, .kernel(kernels[836]), .conv_out(xor_out[836]));
convchan2 c_2_837 (.image, .kernel(kernels[837]), .conv_out(xor_out[837]));
convchan2 c_2_838 (.image, .kernel(kernels[838]), .conv_out(xor_out[838]));
convchan2 c_2_839 (.image, .kernel(kernels[839]), .conv_out(xor_out[839]));
convchan2 c_2_840 (.image, .kernel(kernels[840]), .conv_out(xor_out[840]));
convchan2 c_2_841 (.image, .kernel(kernels[841]), .conv_out(xor_out[841]));
convchan2 c_2_842 (.image, .kernel(kernels[842]), .conv_out(xor_out[842]));
convchan2 c_2_843 (.image, .kernel(kernels[843]), .conv_out(xor_out[843]));
convchan2 c_2_844 (.image, .kernel(kernels[844]), .conv_out(xor_out[844]));
convchan2 c_2_845 (.image, .kernel(kernels[845]), .conv_out(xor_out[845]));
convchan2 c_2_846 (.image, .kernel(kernels[846]), .conv_out(xor_out[846]));
convchan2 c_2_847 (.image, .kernel(kernels[847]), .conv_out(xor_out[847]));
convchan2 c_2_848 (.image, .kernel(kernels[848]), .conv_out(xor_out[848]));
convchan2 c_2_849 (.image, .kernel(kernels[849]), .conv_out(xor_out[849]));
convchan2 c_2_850 (.image, .kernel(kernels[850]), .conv_out(xor_out[850]));
convchan2 c_2_851 (.image, .kernel(kernels[851]), .conv_out(xor_out[851]));
convchan2 c_2_852 (.image, .kernel(kernels[852]), .conv_out(xor_out[852]));
convchan2 c_2_853 (.image, .kernel(kernels[853]), .conv_out(xor_out[853]));
convchan2 c_2_854 (.image, .kernel(kernels[854]), .conv_out(xor_out[854]));
convchan2 c_2_855 (.image, .kernel(kernels[855]), .conv_out(xor_out[855]));
convchan2 c_2_856 (.image, .kernel(kernels[856]), .conv_out(xor_out[856]));
convchan2 c_2_857 (.image, .kernel(kernels[857]), .conv_out(xor_out[857]));
convchan2 c_2_858 (.image, .kernel(kernels[858]), .conv_out(xor_out[858]));
convchan2 c_2_859 (.image, .kernel(kernels[859]), .conv_out(xor_out[859]));
convchan2 c_2_860 (.image, .kernel(kernels[860]), .conv_out(xor_out[860]));
convchan2 c_2_861 (.image, .kernel(kernels[861]), .conv_out(xor_out[861]));
convchan2 c_2_862 (.image, .kernel(kernels[862]), .conv_out(xor_out[862]));
convchan2 c_2_863 (.image, .kernel(kernels[863]), .conv_out(xor_out[863]));
convchan2 c_2_864 (.image, .kernel(kernels[864]), .conv_out(xor_out[864]));
convchan2 c_2_865 (.image, .kernel(kernels[865]), .conv_out(xor_out[865]));
convchan2 c_2_866 (.image, .kernel(kernels[866]), .conv_out(xor_out[866]));
convchan2 c_2_867 (.image, .kernel(kernels[867]), .conv_out(xor_out[867]));
convchan2 c_2_868 (.image, .kernel(kernels[868]), .conv_out(xor_out[868]));
convchan2 c_2_869 (.image, .kernel(kernels[869]), .conv_out(xor_out[869]));
convchan2 c_2_870 (.image, .kernel(kernels[870]), .conv_out(xor_out[870]));
convchan2 c_2_871 (.image, .kernel(kernels[871]), .conv_out(xor_out[871]));
convchan2 c_2_872 (.image, .kernel(kernels[872]), .conv_out(xor_out[872]));
convchan2 c_2_873 (.image, .kernel(kernels[873]), .conv_out(xor_out[873]));
convchan2 c_2_874 (.image, .kernel(kernels[874]), .conv_out(xor_out[874]));
convchan2 c_2_875 (.image, .kernel(kernels[875]), .conv_out(xor_out[875]));
convchan2 c_2_876 (.image, .kernel(kernels[876]), .conv_out(xor_out[876]));
convchan2 c_2_877 (.image, .kernel(kernels[877]), .conv_out(xor_out[877]));
convchan2 c_2_878 (.image, .kernel(kernels[878]), .conv_out(xor_out[878]));
convchan2 c_2_879 (.image, .kernel(kernels[879]), .conv_out(xor_out[879]));
convchan2 c_2_880 (.image, .kernel(kernels[880]), .conv_out(xor_out[880]));
convchan2 c_2_881 (.image, .kernel(kernels[881]), .conv_out(xor_out[881]));
convchan2 c_2_882 (.image, .kernel(kernels[882]), .conv_out(xor_out[882]));
convchan2 c_2_883 (.image, .kernel(kernels[883]), .conv_out(xor_out[883]));
convchan2 c_2_884 (.image, .kernel(kernels[884]), .conv_out(xor_out[884]));
convchan2 c_2_885 (.image, .kernel(kernels[885]), .conv_out(xor_out[885]));
convchan2 c_2_886 (.image, .kernel(kernels[886]), .conv_out(xor_out[886]));
convchan2 c_2_887 (.image, .kernel(kernels[887]), .conv_out(xor_out[887]));
convchan2 c_2_888 (.image, .kernel(kernels[888]), .conv_out(xor_out[888]));
convchan2 c_2_889 (.image, .kernel(kernels[889]), .conv_out(xor_out[889]));
convchan2 c_2_890 (.image, .kernel(kernels[890]), .conv_out(xor_out[890]));
convchan2 c_2_891 (.image, .kernel(kernels[891]), .conv_out(xor_out[891]));
convchan2 c_2_892 (.image, .kernel(kernels[892]), .conv_out(xor_out[892]));
convchan2 c_2_893 (.image, .kernel(kernels[893]), .conv_out(xor_out[893]));
convchan2 c_2_894 (.image, .kernel(kernels[894]), .conv_out(xor_out[894]));
convchan2 c_2_895 (.image, .kernel(kernels[895]), .conv_out(xor_out[895]));
convchan2 c_2_896 (.image, .kernel(kernels[896]), .conv_out(xor_out[896]));
convchan2 c_2_897 (.image, .kernel(kernels[897]), .conv_out(xor_out[897]));
convchan2 c_2_898 (.image, .kernel(kernels[898]), .conv_out(xor_out[898]));
convchan2 c_2_899 (.image, .kernel(kernels[899]), .conv_out(xor_out[899]));
convchan2 c_2_900 (.image, .kernel(kernels[900]), .conv_out(xor_out[900]));
convchan2 c_2_901 (.image, .kernel(kernels[901]), .conv_out(xor_out[901]));
convchan2 c_2_902 (.image, .kernel(kernels[902]), .conv_out(xor_out[902]));
convchan2 c_2_903 (.image, .kernel(kernels[903]), .conv_out(xor_out[903]));
convchan2 c_2_904 (.image, .kernel(kernels[904]), .conv_out(xor_out[904]));
convchan2 c_2_905 (.image, .kernel(kernels[905]), .conv_out(xor_out[905]));
convchan2 c_2_906 (.image, .kernel(kernels[906]), .conv_out(xor_out[906]));
convchan2 c_2_907 (.image, .kernel(kernels[907]), .conv_out(xor_out[907]));
convchan2 c_2_908 (.image, .kernel(kernels[908]), .conv_out(xor_out[908]));
convchan2 c_2_909 (.image, .kernel(kernels[909]), .conv_out(xor_out[909]));
convchan2 c_2_910 (.image, .kernel(kernels[910]), .conv_out(xor_out[910]));
convchan2 c_2_911 (.image, .kernel(kernels[911]), .conv_out(xor_out[911]));
convchan2 c_2_912 (.image, .kernel(kernels[912]), .conv_out(xor_out[912]));
convchan2 c_2_913 (.image, .kernel(kernels[913]), .conv_out(xor_out[913]));
convchan2 c_2_914 (.image, .kernel(kernels[914]), .conv_out(xor_out[914]));
convchan2 c_2_915 (.image, .kernel(kernels[915]), .conv_out(xor_out[915]));
convchan2 c_2_916 (.image, .kernel(kernels[916]), .conv_out(xor_out[916]));
convchan2 c_2_917 (.image, .kernel(kernels[917]), .conv_out(xor_out[917]));
convchan2 c_2_918 (.image, .kernel(kernels[918]), .conv_out(xor_out[918]));
convchan2 c_2_919 (.image, .kernel(kernels[919]), .conv_out(xor_out[919]));
convchan2 c_2_920 (.image, .kernel(kernels[920]), .conv_out(xor_out[920]));
convchan2 c_2_921 (.image, .kernel(kernels[921]), .conv_out(xor_out[921]));
convchan2 c_2_922 (.image, .kernel(kernels[922]), .conv_out(xor_out[922]));
convchan2 c_2_923 (.image, .kernel(kernels[923]), .conv_out(xor_out[923]));
convchan2 c_2_924 (.image, .kernel(kernels[924]), .conv_out(xor_out[924]));
convchan2 c_2_925 (.image, .kernel(kernels[925]), .conv_out(xor_out[925]));
convchan2 c_2_926 (.image, .kernel(kernels[926]), .conv_out(xor_out[926]));
convchan2 c_2_927 (.image, .kernel(kernels[927]), .conv_out(xor_out[927]));
convchan2 c_2_928 (.image, .kernel(kernels[928]), .conv_out(xor_out[928]));
convchan2 c_2_929 (.image, .kernel(kernels[929]), .conv_out(xor_out[929]));
convchan2 c_2_930 (.image, .kernel(kernels[930]), .conv_out(xor_out[930]));
convchan2 c_2_931 (.image, .kernel(kernels[931]), .conv_out(xor_out[931]));
convchan2 c_2_932 (.image, .kernel(kernels[932]), .conv_out(xor_out[932]));
convchan2 c_2_933 (.image, .kernel(kernels[933]), .conv_out(xor_out[933]));
convchan2 c_2_934 (.image, .kernel(kernels[934]), .conv_out(xor_out[934]));
convchan2 c_2_935 (.image, .kernel(kernels[935]), .conv_out(xor_out[935]));
convchan2 c_2_936 (.image, .kernel(kernels[936]), .conv_out(xor_out[936]));
convchan2 c_2_937 (.image, .kernel(kernels[937]), .conv_out(xor_out[937]));
convchan2 c_2_938 (.image, .kernel(kernels[938]), .conv_out(xor_out[938]));
convchan2 c_2_939 (.image, .kernel(kernels[939]), .conv_out(xor_out[939]));
convchan2 c_2_940 (.image, .kernel(kernels[940]), .conv_out(xor_out[940]));
convchan2 c_2_941 (.image, .kernel(kernels[941]), .conv_out(xor_out[941]));
convchan2 c_2_942 (.image, .kernel(kernels[942]), .conv_out(xor_out[942]));
convchan2 c_2_943 (.image, .kernel(kernels[943]), .conv_out(xor_out[943]));
convchan2 c_2_944 (.image, .kernel(kernels[944]), .conv_out(xor_out[944]));
convchan2 c_2_945 (.image, .kernel(kernels[945]), .conv_out(xor_out[945]));
convchan2 c_2_946 (.image, .kernel(kernels[946]), .conv_out(xor_out[946]));
convchan2 c_2_947 (.image, .kernel(kernels[947]), .conv_out(xor_out[947]));
convchan2 c_2_948 (.image, .kernel(kernels[948]), .conv_out(xor_out[948]));
convchan2 c_2_949 (.image, .kernel(kernels[949]), .conv_out(xor_out[949]));
convchan2 c_2_950 (.image, .kernel(kernels[950]), .conv_out(xor_out[950]));
convchan2 c_2_951 (.image, .kernel(kernels[951]), .conv_out(xor_out[951]));
convchan2 c_2_952 (.image, .kernel(kernels[952]), .conv_out(xor_out[952]));
convchan2 c_2_953 (.image, .kernel(kernels[953]), .conv_out(xor_out[953]));
convchan2 c_2_954 (.image, .kernel(kernels[954]), .conv_out(xor_out[954]));
convchan2 c_2_955 (.image, .kernel(kernels[955]), .conv_out(xor_out[955]));
convchan2 c_2_956 (.image, .kernel(kernels[956]), .conv_out(xor_out[956]));
convchan2 c_2_957 (.image, .kernel(kernels[957]), .conv_out(xor_out[957]));
convchan2 c_2_958 (.image, .kernel(kernels[958]), .conv_out(xor_out[958]));
convchan2 c_2_959 (.image, .kernel(kernels[959]), .conv_out(xor_out[959]));
convchan2 c_2_960 (.image, .kernel(kernels[960]), .conv_out(xor_out[960]));
convchan2 c_2_961 (.image, .kernel(kernels[961]), .conv_out(xor_out[961]));
convchan2 c_2_962 (.image, .kernel(kernels[962]), .conv_out(xor_out[962]));
convchan2 c_2_963 (.image, .kernel(kernels[963]), .conv_out(xor_out[963]));
convchan2 c_2_964 (.image, .kernel(kernels[964]), .conv_out(xor_out[964]));
convchan2 c_2_965 (.image, .kernel(kernels[965]), .conv_out(xor_out[965]));
convchan2 c_2_966 (.image, .kernel(kernels[966]), .conv_out(xor_out[966]));
convchan2 c_2_967 (.image, .kernel(kernels[967]), .conv_out(xor_out[967]));
convchan2 c_2_968 (.image, .kernel(kernels[968]), .conv_out(xor_out[968]));
convchan2 c_2_969 (.image, .kernel(kernels[969]), .conv_out(xor_out[969]));
convchan2 c_2_970 (.image, .kernel(kernels[970]), .conv_out(xor_out[970]));
convchan2 c_2_971 (.image, .kernel(kernels[971]), .conv_out(xor_out[971]));
convchan2 c_2_972 (.image, .kernel(kernels[972]), .conv_out(xor_out[972]));
convchan2 c_2_973 (.image, .kernel(kernels[973]), .conv_out(xor_out[973]));
convchan2 c_2_974 (.image, .kernel(kernels[974]), .conv_out(xor_out[974]));
convchan2 c_2_975 (.image, .kernel(kernels[975]), .conv_out(xor_out[975]));
convchan2 c_2_976 (.image, .kernel(kernels[976]), .conv_out(xor_out[976]));
convchan2 c_2_977 (.image, .kernel(kernels[977]), .conv_out(xor_out[977]));
convchan2 c_2_978 (.image, .kernel(kernels[978]), .conv_out(xor_out[978]));
convchan2 c_2_979 (.image, .kernel(kernels[979]), .conv_out(xor_out[979]));
convchan2 c_2_980 (.image, .kernel(kernels[980]), .conv_out(xor_out[980]));
convchan2 c_2_981 (.image, .kernel(kernels[981]), .conv_out(xor_out[981]));
convchan2 c_2_982 (.image, .kernel(kernels[982]), .conv_out(xor_out[982]));
convchan2 c_2_983 (.image, .kernel(kernels[983]), .conv_out(xor_out[983]));
convchan2 c_2_984 (.image, .kernel(kernels[984]), .conv_out(xor_out[984]));
convchan2 c_2_985 (.image, .kernel(kernels[985]), .conv_out(xor_out[985]));
convchan2 c_2_986 (.image, .kernel(kernels[986]), .conv_out(xor_out[986]));
convchan2 c_2_987 (.image, .kernel(kernels[987]), .conv_out(xor_out[987]));
convchan2 c_2_988 (.image, .kernel(kernels[988]), .conv_out(xor_out[988]));
convchan2 c_2_989 (.image, .kernel(kernels[989]), .conv_out(xor_out[989]));
convchan2 c_2_990 (.image, .kernel(kernels[990]), .conv_out(xor_out[990]));
convchan2 c_2_991 (.image, .kernel(kernels[991]), .conv_out(xor_out[991]));
convchan2 c_2_992 (.image, .kernel(kernels[992]), .conv_out(xor_out[992]));
convchan2 c_2_993 (.image, .kernel(kernels[993]), .conv_out(xor_out[993]));
convchan2 c_2_994 (.image, .kernel(kernels[994]), .conv_out(xor_out[994]));
convchan2 c_2_995 (.image, .kernel(kernels[995]), .conv_out(xor_out[995]));
convchan2 c_2_996 (.image, .kernel(kernels[996]), .conv_out(xor_out[996]));
convchan2 c_2_997 (.image, .kernel(kernels[997]), .conv_out(xor_out[997]));
convchan2 c_2_998 (.image, .kernel(kernels[998]), .conv_out(xor_out[998]));
convchan2 c_2_999 (.image, .kernel(kernels[999]), .conv_out(xor_out[999]));
convchan2 c_2_1000 (.image, .kernel(kernels[1000]), .conv_out(xor_out[1000]));
convchan2 c_2_1001 (.image, .kernel(kernels[1001]), .conv_out(xor_out[1001]));
convchan2 c_2_1002 (.image, .kernel(kernels[1002]), .conv_out(xor_out[1002]));
convchan2 c_2_1003 (.image, .kernel(kernels[1003]), .conv_out(xor_out[1003]));
convchan2 c_2_1004 (.image, .kernel(kernels[1004]), .conv_out(xor_out[1004]));
convchan2 c_2_1005 (.image, .kernel(kernels[1005]), .conv_out(xor_out[1005]));
convchan2 c_2_1006 (.image, .kernel(kernels[1006]), .conv_out(xor_out[1006]));
convchan2 c_2_1007 (.image, .kernel(kernels[1007]), .conv_out(xor_out[1007]));
convchan2 c_2_1008 (.image, .kernel(kernels[1008]), .conv_out(xor_out[1008]));
convchan2 c_2_1009 (.image, .kernel(kernels[1009]), .conv_out(xor_out[1009]));
convchan2 c_2_1010 (.image, .kernel(kernels[1010]), .conv_out(xor_out[1010]));
convchan2 c_2_1011 (.image, .kernel(kernels[1011]), .conv_out(xor_out[1011]));
convchan2 c_2_1012 (.image, .kernel(kernels[1012]), .conv_out(xor_out[1012]));
convchan2 c_2_1013 (.image, .kernel(kernels[1013]), .conv_out(xor_out[1013]));
convchan2 c_2_1014 (.image, .kernel(kernels[1014]), .conv_out(xor_out[1014]));
convchan2 c_2_1015 (.image, .kernel(kernels[1015]), .conv_out(xor_out[1015]));
convchan2 c_2_1016 (.image, .kernel(kernels[1016]), .conv_out(xor_out[1016]));
convchan2 c_2_1017 (.image, .kernel(kernels[1017]), .conv_out(xor_out[1017]));
convchan2 c_2_1018 (.image, .kernel(kernels[1018]), .conv_out(xor_out[1018]));
convchan2 c_2_1019 (.image, .kernel(kernels[1019]), .conv_out(xor_out[1019]));
convchan2 c_2_1020 (.image, .kernel(kernels[1020]), .conv_out(xor_out[1020]));
convchan2 c_2_1021 (.image, .kernel(kernels[1021]), .conv_out(xor_out[1021]));
convchan2 c_2_1022 (.image, .kernel(kernels[1022]), .conv_out(xor_out[1022]));
convchan2 c_2_1023 (.image, .kernel(kernels[1023]), .conv_out(xor_out[1023]));
convchan2 c_2_1024 (.image, .kernel(kernels[1024]), .conv_out(xor_out[1024]));
convchan2 c_2_1025 (.image, .kernel(kernels[1025]), .conv_out(xor_out[1025]));
convchan2 c_2_1026 (.image, .kernel(kernels[1026]), .conv_out(xor_out[1026]));
convchan2 c_2_1027 (.image, .kernel(kernels[1027]), .conv_out(xor_out[1027]));
convchan2 c_2_1028 (.image, .kernel(kernels[1028]), .conv_out(xor_out[1028]));
convchan2 c_2_1029 (.image, .kernel(kernels[1029]), .conv_out(xor_out[1029]));
convchan2 c_2_1030 (.image, .kernel(kernels[1030]), .conv_out(xor_out[1030]));
convchan2 c_2_1031 (.image, .kernel(kernels[1031]), .conv_out(xor_out[1031]));
convchan2 c_2_1032 (.image, .kernel(kernels[1032]), .conv_out(xor_out[1032]));
convchan2 c_2_1033 (.image, .kernel(kernels[1033]), .conv_out(xor_out[1033]));
convchan2 c_2_1034 (.image, .kernel(kernels[1034]), .conv_out(xor_out[1034]));
convchan2 c_2_1035 (.image, .kernel(kernels[1035]), .conv_out(xor_out[1035]));
convchan2 c_2_1036 (.image, .kernel(kernels[1036]), .conv_out(xor_out[1036]));
convchan2 c_2_1037 (.image, .kernel(kernels[1037]), .conv_out(xor_out[1037]));
convchan2 c_2_1038 (.image, .kernel(kernels[1038]), .conv_out(xor_out[1038]));
convchan2 c_2_1039 (.image, .kernel(kernels[1039]), .conv_out(xor_out[1039]));
convchan2 c_2_1040 (.image, .kernel(kernels[1040]), .conv_out(xor_out[1040]));
convchan2 c_2_1041 (.image, .kernel(kernels[1041]), .conv_out(xor_out[1041]));
convchan2 c_2_1042 (.image, .kernel(kernels[1042]), .conv_out(xor_out[1042]));
convchan2 c_2_1043 (.image, .kernel(kernels[1043]), .conv_out(xor_out[1043]));
convchan2 c_2_1044 (.image, .kernel(kernels[1044]), .conv_out(xor_out[1044]));
convchan2 c_2_1045 (.image, .kernel(kernels[1045]), .conv_out(xor_out[1045]));
convchan2 c_2_1046 (.image, .kernel(kernels[1046]), .conv_out(xor_out[1046]));
convchan2 c_2_1047 (.image, .kernel(kernels[1047]), .conv_out(xor_out[1047]));
convchan2 c_2_1048 (.image, .kernel(kernels[1048]), .conv_out(xor_out[1048]));
convchan2 c_2_1049 (.image, .kernel(kernels[1049]), .conv_out(xor_out[1049]));
convchan2 c_2_1050 (.image, .kernel(kernels[1050]), .conv_out(xor_out[1050]));
convchan2 c_2_1051 (.image, .kernel(kernels[1051]), .conv_out(xor_out[1051]));
convchan2 c_2_1052 (.image, .kernel(kernels[1052]), .conv_out(xor_out[1052]));
convchan2 c_2_1053 (.image, .kernel(kernels[1053]), .conv_out(xor_out[1053]));
convchan2 c_2_1054 (.image, .kernel(kernels[1054]), .conv_out(xor_out[1054]));
convchan2 c_2_1055 (.image, .kernel(kernels[1055]), .conv_out(xor_out[1055]));
convchan2 c_2_1056 (.image, .kernel(kernels[1056]), .conv_out(xor_out[1056]));
convchan2 c_2_1057 (.image, .kernel(kernels[1057]), .conv_out(xor_out[1057]));
convchan2 c_2_1058 (.image, .kernel(kernels[1058]), .conv_out(xor_out[1058]));
convchan2 c_2_1059 (.image, .kernel(kernels[1059]), .conv_out(xor_out[1059]));
convchan2 c_2_1060 (.image, .kernel(kernels[1060]), .conv_out(xor_out[1060]));
convchan2 c_2_1061 (.image, .kernel(kernels[1061]), .conv_out(xor_out[1061]));
convchan2 c_2_1062 (.image, .kernel(kernels[1062]), .conv_out(xor_out[1062]));
convchan2 c_2_1063 (.image, .kernel(kernels[1063]), .conv_out(xor_out[1063]));
convchan2 c_2_1064 (.image, .kernel(kernels[1064]), .conv_out(xor_out[1064]));
convchan2 c_2_1065 (.image, .kernel(kernels[1065]), .conv_out(xor_out[1065]));
convchan2 c_2_1066 (.image, .kernel(kernels[1066]), .conv_out(xor_out[1066]));
convchan2 c_2_1067 (.image, .kernel(kernels[1067]), .conv_out(xor_out[1067]));
convchan2 c_2_1068 (.image, .kernel(kernels[1068]), .conv_out(xor_out[1068]));
convchan2 c_2_1069 (.image, .kernel(kernels[1069]), .conv_out(xor_out[1069]));
convchan2 c_2_1070 (.image, .kernel(kernels[1070]), .conv_out(xor_out[1070]));
convchan2 c_2_1071 (.image, .kernel(kernels[1071]), .conv_out(xor_out[1071]));
convchan2 c_2_1072 (.image, .kernel(kernels[1072]), .conv_out(xor_out[1072]));
convchan2 c_2_1073 (.image, .kernel(kernels[1073]), .conv_out(xor_out[1073]));
convchan2 c_2_1074 (.image, .kernel(kernels[1074]), .conv_out(xor_out[1074]));
convchan2 c_2_1075 (.image, .kernel(kernels[1075]), .conv_out(xor_out[1075]));
convchan2 c_2_1076 (.image, .kernel(kernels[1076]), .conv_out(xor_out[1076]));
convchan2 c_2_1077 (.image, .kernel(kernels[1077]), .conv_out(xor_out[1077]));
convchan2 c_2_1078 (.image, .kernel(kernels[1078]), .conv_out(xor_out[1078]));
convchan2 c_2_1079 (.image, .kernel(kernels[1079]), .conv_out(xor_out[1079]));

accbin2 ab_2_0 (.accbin_in(xor_out[0:19]), .kernel_offset(kernel_offset[0]), .accbin_out(conv_one_out[0]));
accbin2 ab_2_1 (.accbin_in(xor_out[60:79]), .kernel_offset(kernel_offset[1]), .accbin_out(conv_one_out[1]));
accbin2 ab_2_2 (.accbin_in(xor_out[120:139]), .kernel_offset(kernel_offset[2]), .accbin_out(conv_one_out[2]));
accbin2 ab_2_3 (.accbin_in(xor_out[180:199]), .kernel_offset(kernel_offset[3]), .accbin_out(conv_one_out[3]));
accbin2 ab_2_4 (.accbin_in(xor_out[240:259]), .kernel_offset(kernel_offset[4]), .accbin_out(conv_one_out[4]));
accbin2 ab_2_5 (.accbin_in(xor_out[300:319]), .kernel_offset(kernel_offset[5]), .accbin_out(conv_one_out[5]));
accbin2 ab_2_6 (.accbin_in(xor_out[360:379]), .kernel_offset(kernel_offset[6]), .accbin_out(conv_one_out[6]));
accbin2 ab_2_7 (.accbin_in(xor_out[420:439]), .kernel_offset(kernel_offset[7]), .accbin_out(conv_one_out[7]));
accbin2 ab_2_8 (.accbin_in(xor_out[480:499]), .kernel_offset(kernel_offset[8]), .accbin_out(conv_one_out[8]));
accbin2 ab_2_9 (.accbin_in(xor_out[540:559]), .kernel_offset(kernel_offset[9]), .accbin_out(conv_one_out[9]));
accbin2 ab_2_10 (.accbin_in(xor_out[600:619]), .kernel_offset(kernel_offset[10]), .accbin_out(conv_one_out[10]));
accbin2 ab_2_11 (.accbin_in(xor_out[660:679]), .kernel_offset(kernel_offset[11]), .accbin_out(conv_one_out[11]));
accbin2 ab_2_12 (.accbin_in(xor_out[720:739]), .kernel_offset(kernel_offset[12]), .accbin_out(conv_one_out[12]));
accbin2 ab_2_13 (.accbin_in(xor_out[780:799]), .kernel_offset(kernel_offset[13]), .accbin_out(conv_one_out[13]));
accbin2 ab_2_14 (.accbin_in(xor_out[840:859]), .kernel_offset(kernel_offset[14]), .accbin_out(conv_one_out[14]));
accbin2 ab_2_15 (.accbin_in(xor_out[900:919]), .kernel_offset(kernel_offset[15]), .accbin_out(conv_one_out[15]));
accbin2 ab_2_16 (.accbin_in(xor_out[960:979]), .kernel_offset(kernel_offset[16]), .accbin_out(conv_one_out[16]));
accbin2 ab_2_17 (.accbin_in(xor_out[1020:1039]), .kernel_offset(kernel_offset[17]), .accbin_out(conv_one_out[17]));
accbin2 ab_2_18 (.accbin_in(xor_out[1080:1099]), .kernel_offset(kernel_offset[18]), .accbin_out(conv_one_out[18]));
accbin2 ab_2_19 (.accbin_in(xor_out[1140:1159]), .kernel_offset(kernel_offset[19]), .accbin_out(conv_one_out[19]));
accbin2 ab_2_20 (.accbin_in(xor_out[1200:1219]), .kernel_offset(kernel_offset[20]), .accbin_out(conv_one_out[20]));
accbin2 ab_2_21 (.accbin_in(xor_out[1260:1279]), .kernel_offset(kernel_offset[21]), .accbin_out(conv_one_out[21]));
accbin2 ab_2_22 (.accbin_in(xor_out[1320:1339]), .kernel_offset(kernel_offset[22]), .accbin_out(conv_one_out[22]));
accbin2 ab_2_23 (.accbin_in(xor_out[1380:1399]), .kernel_offset(kernel_offset[23]), .accbin_out(conv_one_out[23]));
accbin2 ab_2_24 (.accbin_in(xor_out[1440:1459]), .kernel_offset(kernel_offset[24]), .accbin_out(conv_one_out[24]));
accbin2 ab_2_25 (.accbin_in(xor_out[1500:1519]), .kernel_offset(kernel_offset[25]), .accbin_out(conv_one_out[25]));
accbin2 ab_2_26 (.accbin_in(xor_out[1560:1579]), .kernel_offset(kernel_offset[26]), .accbin_out(conv_one_out[26]));
accbin2 ab_2_27 (.accbin_in(xor_out[1620:1639]), .kernel_offset(kernel_offset[27]), .accbin_out(conv_one_out[27]));
accbin2 ab_2_28 (.accbin_in(xor_out[1680:1699]), .kernel_offset(kernel_offset[28]), .accbin_out(conv_one_out[28]));
accbin2 ab_2_29 (.accbin_in(xor_out[1740:1759]), .kernel_offset(kernel_offset[29]), .accbin_out(conv_one_out[29]));
accbin2 ab_2_30 (.accbin_in(xor_out[1800:1819]), .kernel_offset(kernel_offset[30]), .accbin_out(conv_one_out[30]));
accbin2 ab_2_31 (.accbin_in(xor_out[1860:1879]), .kernel_offset(kernel_offset[31]), .accbin_out(conv_one_out[31]));
accbin2 ab_2_32 (.accbin_in(xor_out[1920:1939]), .kernel_offset(kernel_offset[32]), .accbin_out(conv_one_out[32]));
accbin2 ab_2_33 (.accbin_in(xor_out[1980:1999]), .kernel_offset(kernel_offset[33]), .accbin_out(conv_one_out[33]));
accbin2 ab_2_34 (.accbin_in(xor_out[2040:2059]), .kernel_offset(kernel_offset[34]), .accbin_out(conv_one_out[34]));
accbin2 ab_2_35 (.accbin_in(xor_out[2100:2119]), .kernel_offset(kernel_offset[35]), .accbin_out(conv_one_out[35]));
accbin2 ab_2_36 (.accbin_in(xor_out[2160:2179]), .kernel_offset(kernel_offset[36]), .accbin_out(conv_one_out[36]));
accbin2 ab_2_37 (.accbin_in(xor_out[2220:2239]), .kernel_offset(kernel_offset[37]), .accbin_out(conv_one_out[37]));
accbin2 ab_2_38 (.accbin_in(xor_out[2280:2299]), .kernel_offset(kernel_offset[38]), .accbin_out(conv_one_out[38]));
accbin2 ab_2_39 (.accbin_in(xor_out[2340:2359]), .kernel_offset(kernel_offset[39]), .accbin_out(conv_one_out[39]));
accbin2 ab_2_40 (.accbin_in(xor_out[2400:2419]), .kernel_offset(kernel_offset[40]), .accbin_out(conv_one_out[40]));
accbin2 ab_2_41 (.accbin_in(xor_out[2460:2479]), .kernel_offset(kernel_offset[41]), .accbin_out(conv_one_out[41]));
accbin2 ab_2_42 (.accbin_in(xor_out[2520:2539]), .kernel_offset(kernel_offset[42]), .accbin_out(conv_one_out[42]));
accbin2 ab_2_43 (.accbin_in(xor_out[2580:2599]), .kernel_offset(kernel_offset[43]), .accbin_out(conv_one_out[43]));
accbin2 ab_2_44 (.accbin_in(xor_out[2640:2659]), .kernel_offset(kernel_offset[44]), .accbin_out(conv_one_out[44]));
accbin2 ab_2_45 (.accbin_in(xor_out[2700:2719]), .kernel_offset(kernel_offset[45]), .accbin_out(conv_one_out[45]));
accbin2 ab_2_46 (.accbin_in(xor_out[2760:2779]), .kernel_offset(kernel_offset[46]), .accbin_out(conv_one_out[46]));
accbin2 ab_2_47 (.accbin_in(xor_out[2820:2839]), .kernel_offset(kernel_offset[47]), .accbin_out(conv_one_out[47]));
accbin2 ab_2_48 (.accbin_in(xor_out[2880:2899]), .kernel_offset(kernel_offset[48]), .accbin_out(conv_one_out[48]));
accbin2 ab_2_49 (.accbin_in(xor_out[2940:2959]), .kernel_offset(kernel_offset[49]), .accbin_out(conv_one_out[49]));
accbin2 ab_2_50 (.accbin_in(xor_out[3000:3019]), .kernel_offset(kernel_offset[50]), .accbin_out(conv_one_out[50]));
accbin2 ab_2_51 (.accbin_in(xor_out[3060:3079]), .kernel_offset(kernel_offset[51]), .accbin_out(conv_one_out[51]));
accbin2 ab_2_52 (.accbin_in(xor_out[3120:3139]), .kernel_offset(kernel_offset[52]), .accbin_out(conv_one_out[52]));
accbin2 ab_2_53 (.accbin_in(xor_out[3180:3199]), .kernel_offset(kernel_offset[53]), .accbin_out(conv_one_out[53]));
accbin2 ab_2_54 (.accbin_in(xor_out[3240:3259]), .kernel_offset(kernel_offset[54]), .accbin_out(conv_one_out[54]));
accbin2 ab_2_55 (.accbin_in(xor_out[3300:3319]), .kernel_offset(kernel_offset[55]), .accbin_out(conv_one_out[55]));
accbin2 ab_2_56 (.accbin_in(xor_out[3360:3379]), .kernel_offset(kernel_offset[56]), .accbin_out(conv_one_out[56]));
accbin2 ab_2_57 (.accbin_in(xor_out[3420:3439]), .kernel_offset(kernel_offset[57]), .accbin_out(conv_one_out[57]));
accbin2 ab_2_58 (.accbin_in(xor_out[3480:3499]), .kernel_offset(kernel_offset[58]), .accbin_out(conv_one_out[58]));
accbin2 ab_2_59 (.accbin_in(xor_out[3540:3559]), .kernel_offset(kernel_offset[59]), .accbin_out(conv_one_out[59]));

endmodule