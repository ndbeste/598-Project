module conv2_120
    #( parameter bW = 8 )
    (
    input  logic [0:2*12*12    -1]    image         ,
    input  logic [0:2*60*5*5   -1]    kernels       ,
    output logic [0:2*60*8*8*bW-1]    xor_out 
    );

convchan2 c_2_0 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[0*5*5:1*5*5-1]), .o_out_fmap(xor_out[0*8*8*bW:1*8*8*bW-1]));
convchan2 c_2_1 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[1*5*5:2*5*5-1]), .o_out_fmap(xor_out[1*8*8*bW:2*8*8*bW-1]));
convchan2 c_2_2 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[2*5*5:3*5*5-1]), .o_out_fmap(xor_out[2*8*8*bW:3*8*8*bW-1]));
convchan2 c_2_3 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[3*5*5:4*5*5-1]), .o_out_fmap(xor_out[3*8*8*bW:4*8*8*bW-1]));
convchan2 c_2_4 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[4*5*5:5*5*5-1]), .o_out_fmap(xor_out[4*8*8*bW:5*8*8*bW-1]));
convchan2 c_2_5 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[5*5*5:6*5*5-1]), .o_out_fmap(xor_out[5*8*8*bW:6*8*8*bW-1]));
convchan2 c_2_6 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[6*5*5:7*5*5-1]), .o_out_fmap(xor_out[6*8*8*bW:7*8*8*bW-1]));
convchan2 c_2_7 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[7*5*5:8*5*5-1]), .o_out_fmap(xor_out[7*8*8*bW:8*8*8*bW-1]));
convchan2 c_2_8 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[8*5*5:9*5*5-1]), .o_out_fmap(xor_out[8*8*8*bW:9*8*8*bW-1]));
convchan2 c_2_9 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[9*5*5:10*5*5-1]), .o_out_fmap(xor_out[9*8*8*bW:10*8*8*bW-1]));
convchan2 c_2_10 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[10*5*5:11*5*5-1]), .o_out_fmap(xor_out[10*8*8*bW:11*8*8*bW-1]));
convchan2 c_2_11 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[11*5*5:12*5*5-1]), .o_out_fmap(xor_out[11*8*8*bW:12*8*8*bW-1]));
convchan2 c_2_12 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[12*5*5:13*5*5-1]), .o_out_fmap(xor_out[12*8*8*bW:13*8*8*bW-1]));
convchan2 c_2_13 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[13*5*5:14*5*5-1]), .o_out_fmap(xor_out[13*8*8*bW:14*8*8*bW-1]));
convchan2 c_2_14 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[14*5*5:15*5*5-1]), .o_out_fmap(xor_out[14*8*8*bW:15*8*8*bW-1]));
convchan2 c_2_15 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[15*5*5:16*5*5-1]), .o_out_fmap(xor_out[15*8*8*bW:16*8*8*bW-1]));
convchan2 c_2_16 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[16*5*5:17*5*5-1]), .o_out_fmap(xor_out[16*8*8*bW:17*8*8*bW-1]));
convchan2 c_2_17 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[17*5*5:18*5*5-1]), .o_out_fmap(xor_out[17*8*8*bW:18*8*8*bW-1]));
convchan2 c_2_18 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[18*5*5:19*5*5-1]), .o_out_fmap(xor_out[18*8*8*bW:19*8*8*bW-1]));
convchan2 c_2_19 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[19*5*5:20*5*5-1]), .o_out_fmap(xor_out[19*8*8*bW:20*8*8*bW-1]));
convchan2 c_2_20 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[20*5*5:21*5*5-1]), .o_out_fmap(xor_out[20*8*8*bW:21*8*8*bW-1]));
convchan2 c_2_21 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[21*5*5:22*5*5-1]), .o_out_fmap(xor_out[21*8*8*bW:22*8*8*bW-1]));
convchan2 c_2_22 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[22*5*5:23*5*5-1]), .o_out_fmap(xor_out[22*8*8*bW:23*8*8*bW-1]));
convchan2 c_2_23 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[23*5*5:24*5*5-1]), .o_out_fmap(xor_out[23*8*8*bW:24*8*8*bW-1]));
convchan2 c_2_24 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[24*5*5:25*5*5-1]), .o_out_fmap(xor_out[24*8*8*bW:25*8*8*bW-1]));
convchan2 c_2_25 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[25*5*5:26*5*5-1]), .o_out_fmap(xor_out[25*8*8*bW:26*8*8*bW-1]));
convchan2 c_2_26 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[26*5*5:27*5*5-1]), .o_out_fmap(xor_out[26*8*8*bW:27*8*8*bW-1]));
convchan2 c_2_27 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[27*5*5:28*5*5-1]), .o_out_fmap(xor_out[27*8*8*bW:28*8*8*bW-1]));
convchan2 c_2_28 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[28*5*5:29*5*5-1]), .o_out_fmap(xor_out[28*8*8*bW:29*8*8*bW-1]));
convchan2 c_2_29 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[29*5*5:30*5*5-1]), .o_out_fmap(xor_out[29*8*8*bW:30*8*8*bW-1]));
convchan2 c_2_30 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[30*5*5:31*5*5-1]), .o_out_fmap(xor_out[30*8*8*bW:31*8*8*bW-1]));
convchan2 c_2_31 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[31*5*5:32*5*5-1]), .o_out_fmap(xor_out[31*8*8*bW:32*8*8*bW-1]));
convchan2 c_2_32 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[32*5*5:33*5*5-1]), .o_out_fmap(xor_out[32*8*8*bW:33*8*8*bW-1]));
convchan2 c_2_33 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[33*5*5:34*5*5-1]), .o_out_fmap(xor_out[33*8*8*bW:34*8*8*bW-1]));
convchan2 c_2_34 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[34*5*5:35*5*5-1]), .o_out_fmap(xor_out[34*8*8*bW:35*8*8*bW-1]));
convchan2 c_2_35 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[35*5*5:36*5*5-1]), .o_out_fmap(xor_out[35*8*8*bW:36*8*8*bW-1]));
convchan2 c_2_36 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[36*5*5:37*5*5-1]), .o_out_fmap(xor_out[36*8*8*bW:37*8*8*bW-1]));
convchan2 c_2_37 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[37*5*5:38*5*5-1]), .o_out_fmap(xor_out[37*8*8*bW:38*8*8*bW-1]));
convchan2 c_2_38 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[38*5*5:39*5*5-1]), .o_out_fmap(xor_out[38*8*8*bW:39*8*8*bW-1]));
convchan2 c_2_39 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[39*5*5:40*5*5-1]), .o_out_fmap(xor_out[39*8*8*bW:40*8*8*bW-1]));
convchan2 c_2_40 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[40*5*5:41*5*5-1]), .o_out_fmap(xor_out[40*8*8*bW:41*8*8*bW-1]));
convchan2 c_2_41 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[41*5*5:42*5*5-1]), .o_out_fmap(xor_out[41*8*8*bW:42*8*8*bW-1]));
convchan2 c_2_42 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[42*5*5:43*5*5-1]), .o_out_fmap(xor_out[42*8*8*bW:43*8*8*bW-1]));
convchan2 c_2_43 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[43*5*5:44*5*5-1]), .o_out_fmap(xor_out[43*8*8*bW:44*8*8*bW-1]));
convchan2 c_2_44 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[44*5*5:45*5*5-1]), .o_out_fmap(xor_out[44*8*8*bW:45*8*8*bW-1]));
convchan2 c_2_45 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[45*5*5:46*5*5-1]), .o_out_fmap(xor_out[45*8*8*bW:46*8*8*bW-1]));
convchan2 c_2_46 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[46*5*5:47*5*5-1]), .o_out_fmap(xor_out[46*8*8*bW:47*8*8*bW-1]));
convchan2 c_2_47 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[47*5*5:48*5*5-1]), .o_out_fmap(xor_out[47*8*8*bW:48*8*8*bW-1]));
convchan2 c_2_48 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[48*5*5:49*5*5-1]), .o_out_fmap(xor_out[48*8*8*bW:49*8*8*bW-1]));
convchan2 c_2_49 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[49*5*5:50*5*5-1]), .o_out_fmap(xor_out[49*8*8*bW:50*8*8*bW-1]));
convchan2 c_2_50 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[50*5*5:51*5*5-1]), .o_out_fmap(xor_out[50*8*8*bW:51*8*8*bW-1]));
convchan2 c_2_51 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[51*5*5:52*5*5-1]), .o_out_fmap(xor_out[51*8*8*bW:52*8*8*bW-1]));
convchan2 c_2_52 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[52*5*5:53*5*5-1]), .o_out_fmap(xor_out[52*8*8*bW:53*8*8*bW-1]));
convchan2 c_2_53 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[53*5*5:54*5*5-1]), .o_out_fmap(xor_out[53*8*8*bW:54*8*8*bW-1]));
convchan2 c_2_54 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[54*5*5:55*5*5-1]), .o_out_fmap(xor_out[54*8*8*bW:55*8*8*bW-1]));
convchan2 c_2_55 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[55*5*5:56*5*5-1]), .o_out_fmap(xor_out[55*8*8*bW:56*8*8*bW-1]));
convchan2 c_2_56 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[56*5*5:57*5*5-1]), .o_out_fmap(xor_out[56*8*8*bW:57*8*8*bW-1]));
convchan2 c_2_57 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[57*5*5:58*5*5-1]), .o_out_fmap(xor_out[57*8*8*bW:58*8*8*bW-1]));
convchan2 c_2_58 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[58*5*5:59*5*5-1]), .o_out_fmap(xor_out[58*8*8*bW:59*8*8*bW-1]));
convchan2 c_2_59 (.i_image(image[0*12*12:1*12*12-1]), .i_kernel(kernels[59*5*5:60*5*5-1]), .o_out_fmap(xor_out[59*8*8*bW:60*8*8*bW-1]));
convchan2 c_2_60 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[60*5*5:61*5*5-1]), .o_out_fmap(xor_out[60*8*8*bW:61*8*8*bW-1]));
convchan2 c_2_61 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[61*5*5:62*5*5-1]), .o_out_fmap(xor_out[61*8*8*bW:62*8*8*bW-1]));
convchan2 c_2_62 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[62*5*5:63*5*5-1]), .o_out_fmap(xor_out[62*8*8*bW:63*8*8*bW-1]));
convchan2 c_2_63 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[63*5*5:64*5*5-1]), .o_out_fmap(xor_out[63*8*8*bW:64*8*8*bW-1]));
convchan2 c_2_64 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[64*5*5:65*5*5-1]), .o_out_fmap(xor_out[64*8*8*bW:65*8*8*bW-1]));
convchan2 c_2_65 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[65*5*5:66*5*5-1]), .o_out_fmap(xor_out[65*8*8*bW:66*8*8*bW-1]));
convchan2 c_2_66 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[66*5*5:67*5*5-1]), .o_out_fmap(xor_out[66*8*8*bW:67*8*8*bW-1]));
convchan2 c_2_67 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[67*5*5:68*5*5-1]), .o_out_fmap(xor_out[67*8*8*bW:68*8*8*bW-1]));
convchan2 c_2_68 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[68*5*5:69*5*5-1]), .o_out_fmap(xor_out[68*8*8*bW:69*8*8*bW-1]));
convchan2 c_2_69 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[69*5*5:70*5*5-1]), .o_out_fmap(xor_out[69*8*8*bW:70*8*8*bW-1]));
convchan2 c_2_70 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[70*5*5:71*5*5-1]), .o_out_fmap(xor_out[70*8*8*bW:71*8*8*bW-1]));
convchan2 c_2_71 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[71*5*5:72*5*5-1]), .o_out_fmap(xor_out[71*8*8*bW:72*8*8*bW-1]));
convchan2 c_2_72 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[72*5*5:73*5*5-1]), .o_out_fmap(xor_out[72*8*8*bW:73*8*8*bW-1]));
convchan2 c_2_73 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[73*5*5:74*5*5-1]), .o_out_fmap(xor_out[73*8*8*bW:74*8*8*bW-1]));
convchan2 c_2_74 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[74*5*5:75*5*5-1]), .o_out_fmap(xor_out[74*8*8*bW:75*8*8*bW-1]));
convchan2 c_2_75 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[75*5*5:76*5*5-1]), .o_out_fmap(xor_out[75*8*8*bW:76*8*8*bW-1]));
convchan2 c_2_76 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[76*5*5:77*5*5-1]), .o_out_fmap(xor_out[76*8*8*bW:77*8*8*bW-1]));
convchan2 c_2_77 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[77*5*5:78*5*5-1]), .o_out_fmap(xor_out[77*8*8*bW:78*8*8*bW-1]));
convchan2 c_2_78 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[78*5*5:79*5*5-1]), .o_out_fmap(xor_out[78*8*8*bW:79*8*8*bW-1]));
convchan2 c_2_79 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[79*5*5:80*5*5-1]), .o_out_fmap(xor_out[79*8*8*bW:80*8*8*bW-1]));
convchan2 c_2_80 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[80*5*5:81*5*5-1]), .o_out_fmap(xor_out[80*8*8*bW:81*8*8*bW-1]));
convchan2 c_2_81 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[81*5*5:82*5*5-1]), .o_out_fmap(xor_out[81*8*8*bW:82*8*8*bW-1]));
convchan2 c_2_82 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[82*5*5:83*5*5-1]), .o_out_fmap(xor_out[82*8*8*bW:83*8*8*bW-1]));
convchan2 c_2_83 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[83*5*5:84*5*5-1]), .o_out_fmap(xor_out[83*8*8*bW:84*8*8*bW-1]));
convchan2 c_2_84 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[84*5*5:85*5*5-1]), .o_out_fmap(xor_out[84*8*8*bW:85*8*8*bW-1]));
convchan2 c_2_85 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[85*5*5:86*5*5-1]), .o_out_fmap(xor_out[85*8*8*bW:86*8*8*bW-1]));
convchan2 c_2_86 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[86*5*5:87*5*5-1]), .o_out_fmap(xor_out[86*8*8*bW:87*8*8*bW-1]));
convchan2 c_2_87 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[87*5*5:88*5*5-1]), .o_out_fmap(xor_out[87*8*8*bW:88*8*8*bW-1]));
convchan2 c_2_88 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[88*5*5:89*5*5-1]), .o_out_fmap(xor_out[88*8*8*bW:89*8*8*bW-1]));
convchan2 c_2_89 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[89*5*5:90*5*5-1]), .o_out_fmap(xor_out[89*8*8*bW:90*8*8*bW-1]));
convchan2 c_2_90 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[90*5*5:91*5*5-1]), .o_out_fmap(xor_out[90*8*8*bW:91*8*8*bW-1]));
convchan2 c_2_91 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[91*5*5:92*5*5-1]), .o_out_fmap(xor_out[91*8*8*bW:92*8*8*bW-1]));
convchan2 c_2_92 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[92*5*5:93*5*5-1]), .o_out_fmap(xor_out[92*8*8*bW:93*8*8*bW-1]));
convchan2 c_2_93 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[93*5*5:94*5*5-1]), .o_out_fmap(xor_out[93*8*8*bW:94*8*8*bW-1]));
convchan2 c_2_94 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[94*5*5:95*5*5-1]), .o_out_fmap(xor_out[94*8*8*bW:95*8*8*bW-1]));
convchan2 c_2_95 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[95*5*5:96*5*5-1]), .o_out_fmap(xor_out[95*8*8*bW:96*8*8*bW-1]));
convchan2 c_2_96 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[96*5*5:97*5*5-1]), .o_out_fmap(xor_out[96*8*8*bW:97*8*8*bW-1]));
convchan2 c_2_97 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[97*5*5:98*5*5-1]), .o_out_fmap(xor_out[97*8*8*bW:98*8*8*bW-1]));
convchan2 c_2_98 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[98*5*5:99*5*5-1]), .o_out_fmap(xor_out[98*8*8*bW:99*8*8*bW-1]));
convchan2 c_2_99 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[99*5*5:100*5*5-1]), .o_out_fmap(xor_out[99*8*8*bW:100*8*8*bW-1]));
convchan2 c_2_100 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[100*5*5:101*5*5-1]), .o_out_fmap(xor_out[100*8*8*bW:101*8*8*bW-1]));
convchan2 c_2_101 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[101*5*5:102*5*5-1]), .o_out_fmap(xor_out[101*8*8*bW:102*8*8*bW-1]));
convchan2 c_2_102 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[102*5*5:103*5*5-1]), .o_out_fmap(xor_out[102*8*8*bW:103*8*8*bW-1]));
convchan2 c_2_103 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[103*5*5:104*5*5-1]), .o_out_fmap(xor_out[103*8*8*bW:104*8*8*bW-1]));
convchan2 c_2_104 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[104*5*5:105*5*5-1]), .o_out_fmap(xor_out[104*8*8*bW:105*8*8*bW-1]));
convchan2 c_2_105 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[105*5*5:106*5*5-1]), .o_out_fmap(xor_out[105*8*8*bW:106*8*8*bW-1]));
convchan2 c_2_106 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[106*5*5:107*5*5-1]), .o_out_fmap(xor_out[106*8*8*bW:107*8*8*bW-1]));
convchan2 c_2_107 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[107*5*5:108*5*5-1]), .o_out_fmap(xor_out[107*8*8*bW:108*8*8*bW-1]));
convchan2 c_2_108 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[108*5*5:109*5*5-1]), .o_out_fmap(xor_out[108*8*8*bW:109*8*8*bW-1]));
convchan2 c_2_109 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[109*5*5:110*5*5-1]), .o_out_fmap(xor_out[109*8*8*bW:110*8*8*bW-1]));
convchan2 c_2_110 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[110*5*5:111*5*5-1]), .o_out_fmap(xor_out[110*8*8*bW:111*8*8*bW-1]));
convchan2 c_2_111 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[111*5*5:112*5*5-1]), .o_out_fmap(xor_out[111*8*8*bW:112*8*8*bW-1]));
convchan2 c_2_112 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[112*5*5:113*5*5-1]), .o_out_fmap(xor_out[112*8*8*bW:113*8*8*bW-1]));
convchan2 c_2_113 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[113*5*5:114*5*5-1]), .o_out_fmap(xor_out[113*8*8*bW:114*8*8*bW-1]));
convchan2 c_2_114 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[114*5*5:115*5*5-1]), .o_out_fmap(xor_out[114*8*8*bW:115*8*8*bW-1]));
convchan2 c_2_115 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[115*5*5:116*5*5-1]), .o_out_fmap(xor_out[115*8*8*bW:116*8*8*bW-1]));
convchan2 c_2_116 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[116*5*5:117*5*5-1]), .o_out_fmap(xor_out[116*8*8*bW:117*8*8*bW-1]));
convchan2 c_2_117 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[117*5*5:118*5*5-1]), .o_out_fmap(xor_out[117*8*8*bW:118*8*8*bW-1]));
convchan2 c_2_118 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[118*5*5:119*5*5-1]), .o_out_fmap(xor_out[118*8*8*bW:119*8*8*bW-1]));
convchan2 c_2_119 (.i_image(image[1*12*12:2*12*12-1]), .i_kernel(kernels[119*5*5:120*5*5-1]), .o_out_fmap(xor_out[119*8*8*bW:120*8*8*bW-1]));

endmodule