module accbin1
    #( parameter bW = 8 )
    (
    input  logic [bW-1:0] accbin_in      [0:4][0:23][0:23],
    input  logic [bW-1:0] kernel_offset,
    output logic          accbin_out          [0:23][0:23]
    );

logic [bW-1:0]    sum_out [0:23][0:23];

assign sum_out[0][0] = accbin_in[0][0][0] + accbin_in[1][0][0] + accbin_in[2][0][0] + accbin_in[3][0][0] + accbin_in[4][0][0];
assign sum_out[0][1] = accbin_in[0][0][1] + accbin_in[1][0][1] + accbin_in[2][0][1] + accbin_in[3][0][1] + accbin_in[4][0][1];
assign sum_out[0][2] = accbin_in[0][0][2] + accbin_in[1][0][2] + accbin_in[2][0][2] + accbin_in[3][0][2] + accbin_in[4][0][2];
assign sum_out[0][3] = accbin_in[0][0][3] + accbin_in[1][0][3] + accbin_in[2][0][3] + accbin_in[3][0][3] + accbin_in[4][0][3];
assign sum_out[0][4] = accbin_in[0][0][4] + accbin_in[1][0][4] + accbin_in[2][0][4] + accbin_in[3][0][4] + accbin_in[4][0][4];
assign sum_out[0][5] = accbin_in[0][0][5] + accbin_in[1][0][5] + accbin_in[2][0][5] + accbin_in[3][0][5] + accbin_in[4][0][5];
assign sum_out[0][6] = accbin_in[0][0][6] + accbin_in[1][0][6] + accbin_in[2][0][6] + accbin_in[3][0][6] + accbin_in[4][0][6];
assign sum_out[0][7] = accbin_in[0][0][7] + accbin_in[1][0][7] + accbin_in[2][0][7] + accbin_in[3][0][7] + accbin_in[4][0][7];
assign sum_out[0][8] = accbin_in[0][0][8] + accbin_in[1][0][8] + accbin_in[2][0][8] + accbin_in[3][0][8] + accbin_in[4][0][8];
assign sum_out[0][9] = accbin_in[0][0][9] + accbin_in[1][0][9] + accbin_in[2][0][9] + accbin_in[3][0][9] + accbin_in[4][0][9];
assign sum_out[0][10] = accbin_in[0][0][10] + accbin_in[1][0][10] + accbin_in[2][0][10] + accbin_in[3][0][10] + accbin_in[4][0][10];
assign sum_out[0][11] = accbin_in[0][0][11] + accbin_in[1][0][11] + accbin_in[2][0][11] + accbin_in[3][0][11] + accbin_in[4][0][11];
assign sum_out[0][12] = accbin_in[0][0][12] + accbin_in[1][0][12] + accbin_in[2][0][12] + accbin_in[3][0][12] + accbin_in[4][0][12];
assign sum_out[0][13] = accbin_in[0][0][13] + accbin_in[1][0][13] + accbin_in[2][0][13] + accbin_in[3][0][13] + accbin_in[4][0][13];
assign sum_out[0][14] = accbin_in[0][0][14] + accbin_in[1][0][14] + accbin_in[2][0][14] + accbin_in[3][0][14] + accbin_in[4][0][14];
assign sum_out[0][15] = accbin_in[0][0][15] + accbin_in[1][0][15] + accbin_in[2][0][15] + accbin_in[3][0][15] + accbin_in[4][0][15];
assign sum_out[0][16] = accbin_in[0][0][16] + accbin_in[1][0][16] + accbin_in[2][0][16] + accbin_in[3][0][16] + accbin_in[4][0][16];
assign sum_out[0][17] = accbin_in[0][0][17] + accbin_in[1][0][17] + accbin_in[2][0][17] + accbin_in[3][0][17] + accbin_in[4][0][17];
assign sum_out[0][18] = accbin_in[0][0][18] + accbin_in[1][0][18] + accbin_in[2][0][18] + accbin_in[3][0][18] + accbin_in[4][0][18];
assign sum_out[0][19] = accbin_in[0][0][19] + accbin_in[1][0][19] + accbin_in[2][0][19] + accbin_in[3][0][19] + accbin_in[4][0][19];
assign sum_out[0][20] = accbin_in[0][0][20] + accbin_in[1][0][20] + accbin_in[2][0][20] + accbin_in[3][0][20] + accbin_in[4][0][20];
assign sum_out[0][21] = accbin_in[0][0][21] + accbin_in[1][0][21] + accbin_in[2][0][21] + accbin_in[3][0][21] + accbin_in[4][0][21];
assign sum_out[0][22] = accbin_in[0][0][22] + accbin_in[1][0][22] + accbin_in[2][0][22] + accbin_in[3][0][22] + accbin_in[4][0][22];
assign sum_out[0][23] = accbin_in[0][0][23] + accbin_in[1][0][23] + accbin_in[2][0][23] + accbin_in[3][0][23] + accbin_in[4][0][23];
assign sum_out[1][0] = accbin_in[0][1][0] + accbin_in[1][1][0] + accbin_in[2][1][0] + accbin_in[3][1][0] + accbin_in[4][1][0];
assign sum_out[1][1] = accbin_in[0][1][1] + accbin_in[1][1][1] + accbin_in[2][1][1] + accbin_in[3][1][1] + accbin_in[4][1][1];
assign sum_out[1][2] = accbin_in[0][1][2] + accbin_in[1][1][2] + accbin_in[2][1][2] + accbin_in[3][1][2] + accbin_in[4][1][2];
assign sum_out[1][3] = accbin_in[0][1][3] + accbin_in[1][1][3] + accbin_in[2][1][3] + accbin_in[3][1][3] + accbin_in[4][1][3];
assign sum_out[1][4] = accbin_in[0][1][4] + accbin_in[1][1][4] + accbin_in[2][1][4] + accbin_in[3][1][4] + accbin_in[4][1][4];
assign sum_out[1][5] = accbin_in[0][1][5] + accbin_in[1][1][5] + accbin_in[2][1][5] + accbin_in[3][1][5] + accbin_in[4][1][5];
assign sum_out[1][6] = accbin_in[0][1][6] + accbin_in[1][1][6] + accbin_in[2][1][6] + accbin_in[3][1][6] + accbin_in[4][1][6];
assign sum_out[1][7] = accbin_in[0][1][7] + accbin_in[1][1][7] + accbin_in[2][1][7] + accbin_in[3][1][7] + accbin_in[4][1][7];
assign sum_out[1][8] = accbin_in[0][1][8] + accbin_in[1][1][8] + accbin_in[2][1][8] + accbin_in[3][1][8] + accbin_in[4][1][8];
assign sum_out[1][9] = accbin_in[0][1][9] + accbin_in[1][1][9] + accbin_in[2][1][9] + accbin_in[3][1][9] + accbin_in[4][1][9];
assign sum_out[1][10] = accbin_in[0][1][10] + accbin_in[1][1][10] + accbin_in[2][1][10] + accbin_in[3][1][10] + accbin_in[4][1][10];
assign sum_out[1][11] = accbin_in[0][1][11] + accbin_in[1][1][11] + accbin_in[2][1][11] + accbin_in[3][1][11] + accbin_in[4][1][11];
assign sum_out[1][12] = accbin_in[0][1][12] + accbin_in[1][1][12] + accbin_in[2][1][12] + accbin_in[3][1][12] + accbin_in[4][1][12];
assign sum_out[1][13] = accbin_in[0][1][13] + accbin_in[1][1][13] + accbin_in[2][1][13] + accbin_in[3][1][13] + accbin_in[4][1][13];
assign sum_out[1][14] = accbin_in[0][1][14] + accbin_in[1][1][14] + accbin_in[2][1][14] + accbin_in[3][1][14] + accbin_in[4][1][14];
assign sum_out[1][15] = accbin_in[0][1][15] + accbin_in[1][1][15] + accbin_in[2][1][15] + accbin_in[3][1][15] + accbin_in[4][1][15];
assign sum_out[1][16] = accbin_in[0][1][16] + accbin_in[1][1][16] + accbin_in[2][1][16] + accbin_in[3][1][16] + accbin_in[4][1][16];
assign sum_out[1][17] = accbin_in[0][1][17] + accbin_in[1][1][17] + accbin_in[2][1][17] + accbin_in[3][1][17] + accbin_in[4][1][17];
assign sum_out[1][18] = accbin_in[0][1][18] + accbin_in[1][1][18] + accbin_in[2][1][18] + accbin_in[3][1][18] + accbin_in[4][1][18];
assign sum_out[1][19] = accbin_in[0][1][19] + accbin_in[1][1][19] + accbin_in[2][1][19] + accbin_in[3][1][19] + accbin_in[4][1][19];
assign sum_out[1][20] = accbin_in[0][1][20] + accbin_in[1][1][20] + accbin_in[2][1][20] + accbin_in[3][1][20] + accbin_in[4][1][20];
assign sum_out[1][21] = accbin_in[0][1][21] + accbin_in[1][1][21] + accbin_in[2][1][21] + accbin_in[3][1][21] + accbin_in[4][1][21];
assign sum_out[1][22] = accbin_in[0][1][22] + accbin_in[1][1][22] + accbin_in[2][1][22] + accbin_in[3][1][22] + accbin_in[4][1][22];
assign sum_out[1][23] = accbin_in[0][1][23] + accbin_in[1][1][23] + accbin_in[2][1][23] + accbin_in[3][1][23] + accbin_in[4][1][23];
assign sum_out[2][0] = accbin_in[0][2][0] + accbin_in[1][2][0] + accbin_in[2][2][0] + accbin_in[3][2][0] + accbin_in[4][2][0];
assign sum_out[2][1] = accbin_in[0][2][1] + accbin_in[1][2][1] + accbin_in[2][2][1] + accbin_in[3][2][1] + accbin_in[4][2][1];
assign sum_out[2][2] = accbin_in[0][2][2] + accbin_in[1][2][2] + accbin_in[2][2][2] + accbin_in[3][2][2] + accbin_in[4][2][2];
assign sum_out[2][3] = accbin_in[0][2][3] + accbin_in[1][2][3] + accbin_in[2][2][3] + accbin_in[3][2][3] + accbin_in[4][2][3];
assign sum_out[2][4] = accbin_in[0][2][4] + accbin_in[1][2][4] + accbin_in[2][2][4] + accbin_in[3][2][4] + accbin_in[4][2][4];
assign sum_out[2][5] = accbin_in[0][2][5] + accbin_in[1][2][5] + accbin_in[2][2][5] + accbin_in[3][2][5] + accbin_in[4][2][5];
assign sum_out[2][6] = accbin_in[0][2][6] + accbin_in[1][2][6] + accbin_in[2][2][6] + accbin_in[3][2][6] + accbin_in[4][2][6];
assign sum_out[2][7] = accbin_in[0][2][7] + accbin_in[1][2][7] + accbin_in[2][2][7] + accbin_in[3][2][7] + accbin_in[4][2][7];
assign sum_out[2][8] = accbin_in[0][2][8] + accbin_in[1][2][8] + accbin_in[2][2][8] + accbin_in[3][2][8] + accbin_in[4][2][8];
assign sum_out[2][9] = accbin_in[0][2][9] + accbin_in[1][2][9] + accbin_in[2][2][9] + accbin_in[3][2][9] + accbin_in[4][2][9];
assign sum_out[2][10] = accbin_in[0][2][10] + accbin_in[1][2][10] + accbin_in[2][2][10] + accbin_in[3][2][10] + accbin_in[4][2][10];
assign sum_out[2][11] = accbin_in[0][2][11] + accbin_in[1][2][11] + accbin_in[2][2][11] + accbin_in[3][2][11] + accbin_in[4][2][11];
assign sum_out[2][12] = accbin_in[0][2][12] + accbin_in[1][2][12] + accbin_in[2][2][12] + accbin_in[3][2][12] + accbin_in[4][2][12];
assign sum_out[2][13] = accbin_in[0][2][13] + accbin_in[1][2][13] + accbin_in[2][2][13] + accbin_in[3][2][13] + accbin_in[4][2][13];
assign sum_out[2][14] = accbin_in[0][2][14] + accbin_in[1][2][14] + accbin_in[2][2][14] + accbin_in[3][2][14] + accbin_in[4][2][14];
assign sum_out[2][15] = accbin_in[0][2][15] + accbin_in[1][2][15] + accbin_in[2][2][15] + accbin_in[3][2][15] + accbin_in[4][2][15];
assign sum_out[2][16] = accbin_in[0][2][16] + accbin_in[1][2][16] + accbin_in[2][2][16] + accbin_in[3][2][16] + accbin_in[4][2][16];
assign sum_out[2][17] = accbin_in[0][2][17] + accbin_in[1][2][17] + accbin_in[2][2][17] + accbin_in[3][2][17] + accbin_in[4][2][17];
assign sum_out[2][18] = accbin_in[0][2][18] + accbin_in[1][2][18] + accbin_in[2][2][18] + accbin_in[3][2][18] + accbin_in[4][2][18];
assign sum_out[2][19] = accbin_in[0][2][19] + accbin_in[1][2][19] + accbin_in[2][2][19] + accbin_in[3][2][19] + accbin_in[4][2][19];
assign sum_out[2][20] = accbin_in[0][2][20] + accbin_in[1][2][20] + accbin_in[2][2][20] + accbin_in[3][2][20] + accbin_in[4][2][20];
assign sum_out[2][21] = accbin_in[0][2][21] + accbin_in[1][2][21] + accbin_in[2][2][21] + accbin_in[3][2][21] + accbin_in[4][2][21];
assign sum_out[2][22] = accbin_in[0][2][22] + accbin_in[1][2][22] + accbin_in[2][2][22] + accbin_in[3][2][22] + accbin_in[4][2][22];
assign sum_out[2][23] = accbin_in[0][2][23] + accbin_in[1][2][23] + accbin_in[2][2][23] + accbin_in[3][2][23] + accbin_in[4][2][23];
assign sum_out[3][0] = accbin_in[0][3][0] + accbin_in[1][3][0] + accbin_in[2][3][0] + accbin_in[3][3][0] + accbin_in[4][3][0];
assign sum_out[3][1] = accbin_in[0][3][1] + accbin_in[1][3][1] + accbin_in[2][3][1] + accbin_in[3][3][1] + accbin_in[4][3][1];
assign sum_out[3][2] = accbin_in[0][3][2] + accbin_in[1][3][2] + accbin_in[2][3][2] + accbin_in[3][3][2] + accbin_in[4][3][2];
assign sum_out[3][3] = accbin_in[0][3][3] + accbin_in[1][3][3] + accbin_in[2][3][3] + accbin_in[3][3][3] + accbin_in[4][3][3];
assign sum_out[3][4] = accbin_in[0][3][4] + accbin_in[1][3][4] + accbin_in[2][3][4] + accbin_in[3][3][4] + accbin_in[4][3][4];
assign sum_out[3][5] = accbin_in[0][3][5] + accbin_in[1][3][5] + accbin_in[2][3][5] + accbin_in[3][3][5] + accbin_in[4][3][5];
assign sum_out[3][6] = accbin_in[0][3][6] + accbin_in[1][3][6] + accbin_in[2][3][6] + accbin_in[3][3][6] + accbin_in[4][3][6];
assign sum_out[3][7] = accbin_in[0][3][7] + accbin_in[1][3][7] + accbin_in[2][3][7] + accbin_in[3][3][7] + accbin_in[4][3][7];
assign sum_out[3][8] = accbin_in[0][3][8] + accbin_in[1][3][8] + accbin_in[2][3][8] + accbin_in[3][3][8] + accbin_in[4][3][8];
assign sum_out[3][9] = accbin_in[0][3][9] + accbin_in[1][3][9] + accbin_in[2][3][9] + accbin_in[3][3][9] + accbin_in[4][3][9];
assign sum_out[3][10] = accbin_in[0][3][10] + accbin_in[1][3][10] + accbin_in[2][3][10] + accbin_in[3][3][10] + accbin_in[4][3][10];
assign sum_out[3][11] = accbin_in[0][3][11] + accbin_in[1][3][11] + accbin_in[2][3][11] + accbin_in[3][3][11] + accbin_in[4][3][11];
assign sum_out[3][12] = accbin_in[0][3][12] + accbin_in[1][3][12] + accbin_in[2][3][12] + accbin_in[3][3][12] + accbin_in[4][3][12];
assign sum_out[3][13] = accbin_in[0][3][13] + accbin_in[1][3][13] + accbin_in[2][3][13] + accbin_in[3][3][13] + accbin_in[4][3][13];
assign sum_out[3][14] = accbin_in[0][3][14] + accbin_in[1][3][14] + accbin_in[2][3][14] + accbin_in[3][3][14] + accbin_in[4][3][14];
assign sum_out[3][15] = accbin_in[0][3][15] + accbin_in[1][3][15] + accbin_in[2][3][15] + accbin_in[3][3][15] + accbin_in[4][3][15];
assign sum_out[3][16] = accbin_in[0][3][16] + accbin_in[1][3][16] + accbin_in[2][3][16] + accbin_in[3][3][16] + accbin_in[4][3][16];
assign sum_out[3][17] = accbin_in[0][3][17] + accbin_in[1][3][17] + accbin_in[2][3][17] + accbin_in[3][3][17] + accbin_in[4][3][17];
assign sum_out[3][18] = accbin_in[0][3][18] + accbin_in[1][3][18] + accbin_in[2][3][18] + accbin_in[3][3][18] + accbin_in[4][3][18];
assign sum_out[3][19] = accbin_in[0][3][19] + accbin_in[1][3][19] + accbin_in[2][3][19] + accbin_in[3][3][19] + accbin_in[4][3][19];
assign sum_out[3][20] = accbin_in[0][3][20] + accbin_in[1][3][20] + accbin_in[2][3][20] + accbin_in[3][3][20] + accbin_in[4][3][20];
assign sum_out[3][21] = accbin_in[0][3][21] + accbin_in[1][3][21] + accbin_in[2][3][21] + accbin_in[3][3][21] + accbin_in[4][3][21];
assign sum_out[3][22] = accbin_in[0][3][22] + accbin_in[1][3][22] + accbin_in[2][3][22] + accbin_in[3][3][22] + accbin_in[4][3][22];
assign sum_out[3][23] = accbin_in[0][3][23] + accbin_in[1][3][23] + accbin_in[2][3][23] + accbin_in[3][3][23] + accbin_in[4][3][23];
assign sum_out[4][0] = accbin_in[0][4][0] + accbin_in[1][4][0] + accbin_in[2][4][0] + accbin_in[3][4][0] + accbin_in[4][4][0];
assign sum_out[4][1] = accbin_in[0][4][1] + accbin_in[1][4][1] + accbin_in[2][4][1] + accbin_in[3][4][1] + accbin_in[4][4][1];
assign sum_out[4][2] = accbin_in[0][4][2] + accbin_in[1][4][2] + accbin_in[2][4][2] + accbin_in[3][4][2] + accbin_in[4][4][2];
assign sum_out[4][3] = accbin_in[0][4][3] + accbin_in[1][4][3] + accbin_in[2][4][3] + accbin_in[3][4][3] + accbin_in[4][4][3];
assign sum_out[4][4] = accbin_in[0][4][4] + accbin_in[1][4][4] + accbin_in[2][4][4] + accbin_in[3][4][4] + accbin_in[4][4][4];
assign sum_out[4][5] = accbin_in[0][4][5] + accbin_in[1][4][5] + accbin_in[2][4][5] + accbin_in[3][4][5] + accbin_in[4][4][5];
assign sum_out[4][6] = accbin_in[0][4][6] + accbin_in[1][4][6] + accbin_in[2][4][6] + accbin_in[3][4][6] + accbin_in[4][4][6];
assign sum_out[4][7] = accbin_in[0][4][7] + accbin_in[1][4][7] + accbin_in[2][4][7] + accbin_in[3][4][7] + accbin_in[4][4][7];
assign sum_out[4][8] = accbin_in[0][4][8] + accbin_in[1][4][8] + accbin_in[2][4][8] + accbin_in[3][4][8] + accbin_in[4][4][8];
assign sum_out[4][9] = accbin_in[0][4][9] + accbin_in[1][4][9] + accbin_in[2][4][9] + accbin_in[3][4][9] + accbin_in[4][4][9];
assign sum_out[4][10] = accbin_in[0][4][10] + accbin_in[1][4][10] + accbin_in[2][4][10] + accbin_in[3][4][10] + accbin_in[4][4][10];
assign sum_out[4][11] = accbin_in[0][4][11] + accbin_in[1][4][11] + accbin_in[2][4][11] + accbin_in[3][4][11] + accbin_in[4][4][11];
assign sum_out[4][12] = accbin_in[0][4][12] + accbin_in[1][4][12] + accbin_in[2][4][12] + accbin_in[3][4][12] + accbin_in[4][4][12];
assign sum_out[4][13] = accbin_in[0][4][13] + accbin_in[1][4][13] + accbin_in[2][4][13] + accbin_in[3][4][13] + accbin_in[4][4][13];
assign sum_out[4][14] = accbin_in[0][4][14] + accbin_in[1][4][14] + accbin_in[2][4][14] + accbin_in[3][4][14] + accbin_in[4][4][14];
assign sum_out[4][15] = accbin_in[0][4][15] + accbin_in[1][4][15] + accbin_in[2][4][15] + accbin_in[3][4][15] + accbin_in[4][4][15];
assign sum_out[4][16] = accbin_in[0][4][16] + accbin_in[1][4][16] + accbin_in[2][4][16] + accbin_in[3][4][16] + accbin_in[4][4][16];
assign sum_out[4][17] = accbin_in[0][4][17] + accbin_in[1][4][17] + accbin_in[2][4][17] + accbin_in[3][4][17] + accbin_in[4][4][17];
assign sum_out[4][18] = accbin_in[0][4][18] + accbin_in[1][4][18] + accbin_in[2][4][18] + accbin_in[3][4][18] + accbin_in[4][4][18];
assign sum_out[4][19] = accbin_in[0][4][19] + accbin_in[1][4][19] + accbin_in[2][4][19] + accbin_in[3][4][19] + accbin_in[4][4][19];
assign sum_out[4][20] = accbin_in[0][4][20] + accbin_in[1][4][20] + accbin_in[2][4][20] + accbin_in[3][4][20] + accbin_in[4][4][20];
assign sum_out[4][21] = accbin_in[0][4][21] + accbin_in[1][4][21] + accbin_in[2][4][21] + accbin_in[3][4][21] + accbin_in[4][4][21];
assign sum_out[4][22] = accbin_in[0][4][22] + accbin_in[1][4][22] + accbin_in[2][4][22] + accbin_in[3][4][22] + accbin_in[4][4][22];
assign sum_out[4][23] = accbin_in[0][4][23] + accbin_in[1][4][23] + accbin_in[2][4][23] + accbin_in[3][4][23] + accbin_in[4][4][23];
assign sum_out[5][0] = accbin_in[0][5][0] + accbin_in[1][5][0] + accbin_in[2][5][0] + accbin_in[3][5][0] + accbin_in[4][5][0];
assign sum_out[5][1] = accbin_in[0][5][1] + accbin_in[1][5][1] + accbin_in[2][5][1] + accbin_in[3][5][1] + accbin_in[4][5][1];
assign sum_out[5][2] = accbin_in[0][5][2] + accbin_in[1][5][2] + accbin_in[2][5][2] + accbin_in[3][5][2] + accbin_in[4][5][2];
assign sum_out[5][3] = accbin_in[0][5][3] + accbin_in[1][5][3] + accbin_in[2][5][3] + accbin_in[3][5][3] + accbin_in[4][5][3];
assign sum_out[5][4] = accbin_in[0][5][4] + accbin_in[1][5][4] + accbin_in[2][5][4] + accbin_in[3][5][4] + accbin_in[4][5][4];
assign sum_out[5][5] = accbin_in[0][5][5] + accbin_in[1][5][5] + accbin_in[2][5][5] + accbin_in[3][5][5] + accbin_in[4][5][5];
assign sum_out[5][6] = accbin_in[0][5][6] + accbin_in[1][5][6] + accbin_in[2][5][6] + accbin_in[3][5][6] + accbin_in[4][5][6];
assign sum_out[5][7] = accbin_in[0][5][7] + accbin_in[1][5][7] + accbin_in[2][5][7] + accbin_in[3][5][7] + accbin_in[4][5][7];
assign sum_out[5][8] = accbin_in[0][5][8] + accbin_in[1][5][8] + accbin_in[2][5][8] + accbin_in[3][5][8] + accbin_in[4][5][8];
assign sum_out[5][9] = accbin_in[0][5][9] + accbin_in[1][5][9] + accbin_in[2][5][9] + accbin_in[3][5][9] + accbin_in[4][5][9];
assign sum_out[5][10] = accbin_in[0][5][10] + accbin_in[1][5][10] + accbin_in[2][5][10] + accbin_in[3][5][10] + accbin_in[4][5][10];
assign sum_out[5][11] = accbin_in[0][5][11] + accbin_in[1][5][11] + accbin_in[2][5][11] + accbin_in[3][5][11] + accbin_in[4][5][11];
assign sum_out[5][12] = accbin_in[0][5][12] + accbin_in[1][5][12] + accbin_in[2][5][12] + accbin_in[3][5][12] + accbin_in[4][5][12];
assign sum_out[5][13] = accbin_in[0][5][13] + accbin_in[1][5][13] + accbin_in[2][5][13] + accbin_in[3][5][13] + accbin_in[4][5][13];
assign sum_out[5][14] = accbin_in[0][5][14] + accbin_in[1][5][14] + accbin_in[2][5][14] + accbin_in[3][5][14] + accbin_in[4][5][14];
assign sum_out[5][15] = accbin_in[0][5][15] + accbin_in[1][5][15] + accbin_in[2][5][15] + accbin_in[3][5][15] + accbin_in[4][5][15];
assign sum_out[5][16] = accbin_in[0][5][16] + accbin_in[1][5][16] + accbin_in[2][5][16] + accbin_in[3][5][16] + accbin_in[4][5][16];
assign sum_out[5][17] = accbin_in[0][5][17] + accbin_in[1][5][17] + accbin_in[2][5][17] + accbin_in[3][5][17] + accbin_in[4][5][17];
assign sum_out[5][18] = accbin_in[0][5][18] + accbin_in[1][5][18] + accbin_in[2][5][18] + accbin_in[3][5][18] + accbin_in[4][5][18];
assign sum_out[5][19] = accbin_in[0][5][19] + accbin_in[1][5][19] + accbin_in[2][5][19] + accbin_in[3][5][19] + accbin_in[4][5][19];
assign sum_out[5][20] = accbin_in[0][5][20] + accbin_in[1][5][20] + accbin_in[2][5][20] + accbin_in[3][5][20] + accbin_in[4][5][20];
assign sum_out[5][21] = accbin_in[0][5][21] + accbin_in[1][5][21] + accbin_in[2][5][21] + accbin_in[3][5][21] + accbin_in[4][5][21];
assign sum_out[5][22] = accbin_in[0][5][22] + accbin_in[1][5][22] + accbin_in[2][5][22] + accbin_in[3][5][22] + accbin_in[4][5][22];
assign sum_out[5][23] = accbin_in[0][5][23] + accbin_in[1][5][23] + accbin_in[2][5][23] + accbin_in[3][5][23] + accbin_in[4][5][23];
assign sum_out[6][0] = accbin_in[0][6][0] + accbin_in[1][6][0] + accbin_in[2][6][0] + accbin_in[3][6][0] + accbin_in[4][6][0];
assign sum_out[6][1] = accbin_in[0][6][1] + accbin_in[1][6][1] + accbin_in[2][6][1] + accbin_in[3][6][1] + accbin_in[4][6][1];
assign sum_out[6][2] = accbin_in[0][6][2] + accbin_in[1][6][2] + accbin_in[2][6][2] + accbin_in[3][6][2] + accbin_in[4][6][2];
assign sum_out[6][3] = accbin_in[0][6][3] + accbin_in[1][6][3] + accbin_in[2][6][3] + accbin_in[3][6][3] + accbin_in[4][6][3];
assign sum_out[6][4] = accbin_in[0][6][4] + accbin_in[1][6][4] + accbin_in[2][6][4] + accbin_in[3][6][4] + accbin_in[4][6][4];
assign sum_out[6][5] = accbin_in[0][6][5] + accbin_in[1][6][5] + accbin_in[2][6][5] + accbin_in[3][6][5] + accbin_in[4][6][5];
assign sum_out[6][6] = accbin_in[0][6][6] + accbin_in[1][6][6] + accbin_in[2][6][6] + accbin_in[3][6][6] + accbin_in[4][6][6];
assign sum_out[6][7] = accbin_in[0][6][7] + accbin_in[1][6][7] + accbin_in[2][6][7] + accbin_in[3][6][7] + accbin_in[4][6][7];
assign sum_out[6][8] = accbin_in[0][6][8] + accbin_in[1][6][8] + accbin_in[2][6][8] + accbin_in[3][6][8] + accbin_in[4][6][8];
assign sum_out[6][9] = accbin_in[0][6][9] + accbin_in[1][6][9] + accbin_in[2][6][9] + accbin_in[3][6][9] + accbin_in[4][6][9];
assign sum_out[6][10] = accbin_in[0][6][10] + accbin_in[1][6][10] + accbin_in[2][6][10] + accbin_in[3][6][10] + accbin_in[4][6][10];
assign sum_out[6][11] = accbin_in[0][6][11] + accbin_in[1][6][11] + accbin_in[2][6][11] + accbin_in[3][6][11] + accbin_in[4][6][11];
assign sum_out[6][12] = accbin_in[0][6][12] + accbin_in[1][6][12] + accbin_in[2][6][12] + accbin_in[3][6][12] + accbin_in[4][6][12];
assign sum_out[6][13] = accbin_in[0][6][13] + accbin_in[1][6][13] + accbin_in[2][6][13] + accbin_in[3][6][13] + accbin_in[4][6][13];
assign sum_out[6][14] = accbin_in[0][6][14] + accbin_in[1][6][14] + accbin_in[2][6][14] + accbin_in[3][6][14] + accbin_in[4][6][14];
assign sum_out[6][15] = accbin_in[0][6][15] + accbin_in[1][6][15] + accbin_in[2][6][15] + accbin_in[3][6][15] + accbin_in[4][6][15];
assign sum_out[6][16] = accbin_in[0][6][16] + accbin_in[1][6][16] + accbin_in[2][6][16] + accbin_in[3][6][16] + accbin_in[4][6][16];
assign sum_out[6][17] = accbin_in[0][6][17] + accbin_in[1][6][17] + accbin_in[2][6][17] + accbin_in[3][6][17] + accbin_in[4][6][17];
assign sum_out[6][18] = accbin_in[0][6][18] + accbin_in[1][6][18] + accbin_in[2][6][18] + accbin_in[3][6][18] + accbin_in[4][6][18];
assign sum_out[6][19] = accbin_in[0][6][19] + accbin_in[1][6][19] + accbin_in[2][6][19] + accbin_in[3][6][19] + accbin_in[4][6][19];
assign sum_out[6][20] = accbin_in[0][6][20] + accbin_in[1][6][20] + accbin_in[2][6][20] + accbin_in[3][6][20] + accbin_in[4][6][20];
assign sum_out[6][21] = accbin_in[0][6][21] + accbin_in[1][6][21] + accbin_in[2][6][21] + accbin_in[3][6][21] + accbin_in[4][6][21];
assign sum_out[6][22] = accbin_in[0][6][22] + accbin_in[1][6][22] + accbin_in[2][6][22] + accbin_in[3][6][22] + accbin_in[4][6][22];
assign sum_out[6][23] = accbin_in[0][6][23] + accbin_in[1][6][23] + accbin_in[2][6][23] + accbin_in[3][6][23] + accbin_in[4][6][23];
assign sum_out[7][0] = accbin_in[0][7][0] + accbin_in[1][7][0] + accbin_in[2][7][0] + accbin_in[3][7][0] + accbin_in[4][7][0];
assign sum_out[7][1] = accbin_in[0][7][1] + accbin_in[1][7][1] + accbin_in[2][7][1] + accbin_in[3][7][1] + accbin_in[4][7][1];
assign sum_out[7][2] = accbin_in[0][7][2] + accbin_in[1][7][2] + accbin_in[2][7][2] + accbin_in[3][7][2] + accbin_in[4][7][2];
assign sum_out[7][3] = accbin_in[0][7][3] + accbin_in[1][7][3] + accbin_in[2][7][3] + accbin_in[3][7][3] + accbin_in[4][7][3];
assign sum_out[7][4] = accbin_in[0][7][4] + accbin_in[1][7][4] + accbin_in[2][7][4] + accbin_in[3][7][4] + accbin_in[4][7][4];
assign sum_out[7][5] = accbin_in[0][7][5] + accbin_in[1][7][5] + accbin_in[2][7][5] + accbin_in[3][7][5] + accbin_in[4][7][5];
assign sum_out[7][6] = accbin_in[0][7][6] + accbin_in[1][7][6] + accbin_in[2][7][6] + accbin_in[3][7][6] + accbin_in[4][7][6];
assign sum_out[7][7] = accbin_in[0][7][7] + accbin_in[1][7][7] + accbin_in[2][7][7] + accbin_in[3][7][7] + accbin_in[4][7][7];
assign sum_out[7][8] = accbin_in[0][7][8] + accbin_in[1][7][8] + accbin_in[2][7][8] + accbin_in[3][7][8] + accbin_in[4][7][8];
assign sum_out[7][9] = accbin_in[0][7][9] + accbin_in[1][7][9] + accbin_in[2][7][9] + accbin_in[3][7][9] + accbin_in[4][7][9];
assign sum_out[7][10] = accbin_in[0][7][10] + accbin_in[1][7][10] + accbin_in[2][7][10] + accbin_in[3][7][10] + accbin_in[4][7][10];
assign sum_out[7][11] = accbin_in[0][7][11] + accbin_in[1][7][11] + accbin_in[2][7][11] + accbin_in[3][7][11] + accbin_in[4][7][11];
assign sum_out[7][12] = accbin_in[0][7][12] + accbin_in[1][7][12] + accbin_in[2][7][12] + accbin_in[3][7][12] + accbin_in[4][7][12];
assign sum_out[7][13] = accbin_in[0][7][13] + accbin_in[1][7][13] + accbin_in[2][7][13] + accbin_in[3][7][13] + accbin_in[4][7][13];
assign sum_out[7][14] = accbin_in[0][7][14] + accbin_in[1][7][14] + accbin_in[2][7][14] + accbin_in[3][7][14] + accbin_in[4][7][14];
assign sum_out[7][15] = accbin_in[0][7][15] + accbin_in[1][7][15] + accbin_in[2][7][15] + accbin_in[3][7][15] + accbin_in[4][7][15];
assign sum_out[7][16] = accbin_in[0][7][16] + accbin_in[1][7][16] + accbin_in[2][7][16] + accbin_in[3][7][16] + accbin_in[4][7][16];
assign sum_out[7][17] = accbin_in[0][7][17] + accbin_in[1][7][17] + accbin_in[2][7][17] + accbin_in[3][7][17] + accbin_in[4][7][17];
assign sum_out[7][18] = accbin_in[0][7][18] + accbin_in[1][7][18] + accbin_in[2][7][18] + accbin_in[3][7][18] + accbin_in[4][7][18];
assign sum_out[7][19] = accbin_in[0][7][19] + accbin_in[1][7][19] + accbin_in[2][7][19] + accbin_in[3][7][19] + accbin_in[4][7][19];
assign sum_out[7][20] = accbin_in[0][7][20] + accbin_in[1][7][20] + accbin_in[2][7][20] + accbin_in[3][7][20] + accbin_in[4][7][20];
assign sum_out[7][21] = accbin_in[0][7][21] + accbin_in[1][7][21] + accbin_in[2][7][21] + accbin_in[3][7][21] + accbin_in[4][7][21];
assign sum_out[7][22] = accbin_in[0][7][22] + accbin_in[1][7][22] + accbin_in[2][7][22] + accbin_in[3][7][22] + accbin_in[4][7][22];
assign sum_out[7][23] = accbin_in[0][7][23] + accbin_in[1][7][23] + accbin_in[2][7][23] + accbin_in[3][7][23] + accbin_in[4][7][23];
assign sum_out[8][0] = accbin_in[0][8][0] + accbin_in[1][8][0] + accbin_in[2][8][0] + accbin_in[3][8][0] + accbin_in[4][8][0];
assign sum_out[8][1] = accbin_in[0][8][1] + accbin_in[1][8][1] + accbin_in[2][8][1] + accbin_in[3][8][1] + accbin_in[4][8][1];
assign sum_out[8][2] = accbin_in[0][8][2] + accbin_in[1][8][2] + accbin_in[2][8][2] + accbin_in[3][8][2] + accbin_in[4][8][2];
assign sum_out[8][3] = accbin_in[0][8][3] + accbin_in[1][8][3] + accbin_in[2][8][3] + accbin_in[3][8][3] + accbin_in[4][8][3];
assign sum_out[8][4] = accbin_in[0][8][4] + accbin_in[1][8][4] + accbin_in[2][8][4] + accbin_in[3][8][4] + accbin_in[4][8][4];
assign sum_out[8][5] = accbin_in[0][8][5] + accbin_in[1][8][5] + accbin_in[2][8][5] + accbin_in[3][8][5] + accbin_in[4][8][5];
assign sum_out[8][6] = accbin_in[0][8][6] + accbin_in[1][8][6] + accbin_in[2][8][6] + accbin_in[3][8][6] + accbin_in[4][8][6];
assign sum_out[8][7] = accbin_in[0][8][7] + accbin_in[1][8][7] + accbin_in[2][8][7] + accbin_in[3][8][7] + accbin_in[4][8][7];
assign sum_out[8][8] = accbin_in[0][8][8] + accbin_in[1][8][8] + accbin_in[2][8][8] + accbin_in[3][8][8] + accbin_in[4][8][8];
assign sum_out[8][9] = accbin_in[0][8][9] + accbin_in[1][8][9] + accbin_in[2][8][9] + accbin_in[3][8][9] + accbin_in[4][8][9];
assign sum_out[8][10] = accbin_in[0][8][10] + accbin_in[1][8][10] + accbin_in[2][8][10] + accbin_in[3][8][10] + accbin_in[4][8][10];
assign sum_out[8][11] = accbin_in[0][8][11] + accbin_in[1][8][11] + accbin_in[2][8][11] + accbin_in[3][8][11] + accbin_in[4][8][11];
assign sum_out[8][12] = accbin_in[0][8][12] + accbin_in[1][8][12] + accbin_in[2][8][12] + accbin_in[3][8][12] + accbin_in[4][8][12];
assign sum_out[8][13] = accbin_in[0][8][13] + accbin_in[1][8][13] + accbin_in[2][8][13] + accbin_in[3][8][13] + accbin_in[4][8][13];
assign sum_out[8][14] = accbin_in[0][8][14] + accbin_in[1][8][14] + accbin_in[2][8][14] + accbin_in[3][8][14] + accbin_in[4][8][14];
assign sum_out[8][15] = accbin_in[0][8][15] + accbin_in[1][8][15] + accbin_in[2][8][15] + accbin_in[3][8][15] + accbin_in[4][8][15];
assign sum_out[8][16] = accbin_in[0][8][16] + accbin_in[1][8][16] + accbin_in[2][8][16] + accbin_in[3][8][16] + accbin_in[4][8][16];
assign sum_out[8][17] = accbin_in[0][8][17] + accbin_in[1][8][17] + accbin_in[2][8][17] + accbin_in[3][8][17] + accbin_in[4][8][17];
assign sum_out[8][18] = accbin_in[0][8][18] + accbin_in[1][8][18] + accbin_in[2][8][18] + accbin_in[3][8][18] + accbin_in[4][8][18];
assign sum_out[8][19] = accbin_in[0][8][19] + accbin_in[1][8][19] + accbin_in[2][8][19] + accbin_in[3][8][19] + accbin_in[4][8][19];
assign sum_out[8][20] = accbin_in[0][8][20] + accbin_in[1][8][20] + accbin_in[2][8][20] + accbin_in[3][8][20] + accbin_in[4][8][20];
assign sum_out[8][21] = accbin_in[0][8][21] + accbin_in[1][8][21] + accbin_in[2][8][21] + accbin_in[3][8][21] + accbin_in[4][8][21];
assign sum_out[8][22] = accbin_in[0][8][22] + accbin_in[1][8][22] + accbin_in[2][8][22] + accbin_in[3][8][22] + accbin_in[4][8][22];
assign sum_out[8][23] = accbin_in[0][8][23] + accbin_in[1][8][23] + accbin_in[2][8][23] + accbin_in[3][8][23] + accbin_in[4][8][23];
assign sum_out[9][0] = accbin_in[0][9][0] + accbin_in[1][9][0] + accbin_in[2][9][0] + accbin_in[3][9][0] + accbin_in[4][9][0];
assign sum_out[9][1] = accbin_in[0][9][1] + accbin_in[1][9][1] + accbin_in[2][9][1] + accbin_in[3][9][1] + accbin_in[4][9][1];
assign sum_out[9][2] = accbin_in[0][9][2] + accbin_in[1][9][2] + accbin_in[2][9][2] + accbin_in[3][9][2] + accbin_in[4][9][2];
assign sum_out[9][3] = accbin_in[0][9][3] + accbin_in[1][9][3] + accbin_in[2][9][3] + accbin_in[3][9][3] + accbin_in[4][9][3];
assign sum_out[9][4] = accbin_in[0][9][4] + accbin_in[1][9][4] + accbin_in[2][9][4] + accbin_in[3][9][4] + accbin_in[4][9][4];
assign sum_out[9][5] = accbin_in[0][9][5] + accbin_in[1][9][5] + accbin_in[2][9][5] + accbin_in[3][9][5] + accbin_in[4][9][5];
assign sum_out[9][6] = accbin_in[0][9][6] + accbin_in[1][9][6] + accbin_in[2][9][6] + accbin_in[3][9][6] + accbin_in[4][9][6];
assign sum_out[9][7] = accbin_in[0][9][7] + accbin_in[1][9][7] + accbin_in[2][9][7] + accbin_in[3][9][7] + accbin_in[4][9][7];
assign sum_out[9][8] = accbin_in[0][9][8] + accbin_in[1][9][8] + accbin_in[2][9][8] + accbin_in[3][9][8] + accbin_in[4][9][8];
assign sum_out[9][9] = accbin_in[0][9][9] + accbin_in[1][9][9] + accbin_in[2][9][9] + accbin_in[3][9][9] + accbin_in[4][9][9];
assign sum_out[9][10] = accbin_in[0][9][10] + accbin_in[1][9][10] + accbin_in[2][9][10] + accbin_in[3][9][10] + accbin_in[4][9][10];
assign sum_out[9][11] = accbin_in[0][9][11] + accbin_in[1][9][11] + accbin_in[2][9][11] + accbin_in[3][9][11] + accbin_in[4][9][11];
assign sum_out[9][12] = accbin_in[0][9][12] + accbin_in[1][9][12] + accbin_in[2][9][12] + accbin_in[3][9][12] + accbin_in[4][9][12];
assign sum_out[9][13] = accbin_in[0][9][13] + accbin_in[1][9][13] + accbin_in[2][9][13] + accbin_in[3][9][13] + accbin_in[4][9][13];
assign sum_out[9][14] = accbin_in[0][9][14] + accbin_in[1][9][14] + accbin_in[2][9][14] + accbin_in[3][9][14] + accbin_in[4][9][14];
assign sum_out[9][15] = accbin_in[0][9][15] + accbin_in[1][9][15] + accbin_in[2][9][15] + accbin_in[3][9][15] + accbin_in[4][9][15];
assign sum_out[9][16] = accbin_in[0][9][16] + accbin_in[1][9][16] + accbin_in[2][9][16] + accbin_in[3][9][16] + accbin_in[4][9][16];
assign sum_out[9][17] = accbin_in[0][9][17] + accbin_in[1][9][17] + accbin_in[2][9][17] + accbin_in[3][9][17] + accbin_in[4][9][17];
assign sum_out[9][18] = accbin_in[0][9][18] + accbin_in[1][9][18] + accbin_in[2][9][18] + accbin_in[3][9][18] + accbin_in[4][9][18];
assign sum_out[9][19] = accbin_in[0][9][19] + accbin_in[1][9][19] + accbin_in[2][9][19] + accbin_in[3][9][19] + accbin_in[4][9][19];
assign sum_out[9][20] = accbin_in[0][9][20] + accbin_in[1][9][20] + accbin_in[2][9][20] + accbin_in[3][9][20] + accbin_in[4][9][20];
assign sum_out[9][21] = accbin_in[0][9][21] + accbin_in[1][9][21] + accbin_in[2][9][21] + accbin_in[3][9][21] + accbin_in[4][9][21];
assign sum_out[9][22] = accbin_in[0][9][22] + accbin_in[1][9][22] + accbin_in[2][9][22] + accbin_in[3][9][22] + accbin_in[4][9][22];
assign sum_out[9][23] = accbin_in[0][9][23] + accbin_in[1][9][23] + accbin_in[2][9][23] + accbin_in[3][9][23] + accbin_in[4][9][23];
assign sum_out[10][0] = accbin_in[0][10][0] + accbin_in[1][10][0] + accbin_in[2][10][0] + accbin_in[3][10][0] + accbin_in[4][10][0];
assign sum_out[10][1] = accbin_in[0][10][1] + accbin_in[1][10][1] + accbin_in[2][10][1] + accbin_in[3][10][1] + accbin_in[4][10][1];
assign sum_out[10][2] = accbin_in[0][10][2] + accbin_in[1][10][2] + accbin_in[2][10][2] + accbin_in[3][10][2] + accbin_in[4][10][2];
assign sum_out[10][3] = accbin_in[0][10][3] + accbin_in[1][10][3] + accbin_in[2][10][3] + accbin_in[3][10][3] + accbin_in[4][10][3];
assign sum_out[10][4] = accbin_in[0][10][4] + accbin_in[1][10][4] + accbin_in[2][10][4] + accbin_in[3][10][4] + accbin_in[4][10][4];
assign sum_out[10][5] = accbin_in[0][10][5] + accbin_in[1][10][5] + accbin_in[2][10][5] + accbin_in[3][10][5] + accbin_in[4][10][5];
assign sum_out[10][6] = accbin_in[0][10][6] + accbin_in[1][10][6] + accbin_in[2][10][6] + accbin_in[3][10][6] + accbin_in[4][10][6];
assign sum_out[10][7] = accbin_in[0][10][7] + accbin_in[1][10][7] + accbin_in[2][10][7] + accbin_in[3][10][7] + accbin_in[4][10][7];
assign sum_out[10][8] = accbin_in[0][10][8] + accbin_in[1][10][8] + accbin_in[2][10][8] + accbin_in[3][10][8] + accbin_in[4][10][8];
assign sum_out[10][9] = accbin_in[0][10][9] + accbin_in[1][10][9] + accbin_in[2][10][9] + accbin_in[3][10][9] + accbin_in[4][10][9];
assign sum_out[10][10] = accbin_in[0][10][10] + accbin_in[1][10][10] + accbin_in[2][10][10] + accbin_in[3][10][10] + accbin_in[4][10][10];
assign sum_out[10][11] = accbin_in[0][10][11] + accbin_in[1][10][11] + accbin_in[2][10][11] + accbin_in[3][10][11] + accbin_in[4][10][11];
assign sum_out[10][12] = accbin_in[0][10][12] + accbin_in[1][10][12] + accbin_in[2][10][12] + accbin_in[3][10][12] + accbin_in[4][10][12];
assign sum_out[10][13] = accbin_in[0][10][13] + accbin_in[1][10][13] + accbin_in[2][10][13] + accbin_in[3][10][13] + accbin_in[4][10][13];
assign sum_out[10][14] = accbin_in[0][10][14] + accbin_in[1][10][14] + accbin_in[2][10][14] + accbin_in[3][10][14] + accbin_in[4][10][14];
assign sum_out[10][15] = accbin_in[0][10][15] + accbin_in[1][10][15] + accbin_in[2][10][15] + accbin_in[3][10][15] + accbin_in[4][10][15];
assign sum_out[10][16] = accbin_in[0][10][16] + accbin_in[1][10][16] + accbin_in[2][10][16] + accbin_in[3][10][16] + accbin_in[4][10][16];
assign sum_out[10][17] = accbin_in[0][10][17] + accbin_in[1][10][17] + accbin_in[2][10][17] + accbin_in[3][10][17] + accbin_in[4][10][17];
assign sum_out[10][18] = accbin_in[0][10][18] + accbin_in[1][10][18] + accbin_in[2][10][18] + accbin_in[3][10][18] + accbin_in[4][10][18];
assign sum_out[10][19] = accbin_in[0][10][19] + accbin_in[1][10][19] + accbin_in[2][10][19] + accbin_in[3][10][19] + accbin_in[4][10][19];
assign sum_out[10][20] = accbin_in[0][10][20] + accbin_in[1][10][20] + accbin_in[2][10][20] + accbin_in[3][10][20] + accbin_in[4][10][20];
assign sum_out[10][21] = accbin_in[0][10][21] + accbin_in[1][10][21] + accbin_in[2][10][21] + accbin_in[3][10][21] + accbin_in[4][10][21];
assign sum_out[10][22] = accbin_in[0][10][22] + accbin_in[1][10][22] + accbin_in[2][10][22] + accbin_in[3][10][22] + accbin_in[4][10][22];
assign sum_out[10][23] = accbin_in[0][10][23] + accbin_in[1][10][23] + accbin_in[2][10][23] + accbin_in[3][10][23] + accbin_in[4][10][23];
assign sum_out[11][0] = accbin_in[0][11][0] + accbin_in[1][11][0] + accbin_in[2][11][0] + accbin_in[3][11][0] + accbin_in[4][11][0];
assign sum_out[11][1] = accbin_in[0][11][1] + accbin_in[1][11][1] + accbin_in[2][11][1] + accbin_in[3][11][1] + accbin_in[4][11][1];
assign sum_out[11][2] = accbin_in[0][11][2] + accbin_in[1][11][2] + accbin_in[2][11][2] + accbin_in[3][11][2] + accbin_in[4][11][2];
assign sum_out[11][3] = accbin_in[0][11][3] + accbin_in[1][11][3] + accbin_in[2][11][3] + accbin_in[3][11][3] + accbin_in[4][11][3];
assign sum_out[11][4] = accbin_in[0][11][4] + accbin_in[1][11][4] + accbin_in[2][11][4] + accbin_in[3][11][4] + accbin_in[4][11][4];
assign sum_out[11][5] = accbin_in[0][11][5] + accbin_in[1][11][5] + accbin_in[2][11][5] + accbin_in[3][11][5] + accbin_in[4][11][5];
assign sum_out[11][6] = accbin_in[0][11][6] + accbin_in[1][11][6] + accbin_in[2][11][6] + accbin_in[3][11][6] + accbin_in[4][11][6];
assign sum_out[11][7] = accbin_in[0][11][7] + accbin_in[1][11][7] + accbin_in[2][11][7] + accbin_in[3][11][7] + accbin_in[4][11][7];
assign sum_out[11][8] = accbin_in[0][11][8] + accbin_in[1][11][8] + accbin_in[2][11][8] + accbin_in[3][11][8] + accbin_in[4][11][8];
assign sum_out[11][9] = accbin_in[0][11][9] + accbin_in[1][11][9] + accbin_in[2][11][9] + accbin_in[3][11][9] + accbin_in[4][11][9];
assign sum_out[11][10] = accbin_in[0][11][10] + accbin_in[1][11][10] + accbin_in[2][11][10] + accbin_in[3][11][10] + accbin_in[4][11][10];
assign sum_out[11][11] = accbin_in[0][11][11] + accbin_in[1][11][11] + accbin_in[2][11][11] + accbin_in[3][11][11] + accbin_in[4][11][11];
assign sum_out[11][12] = accbin_in[0][11][12] + accbin_in[1][11][12] + accbin_in[2][11][12] + accbin_in[3][11][12] + accbin_in[4][11][12];
assign sum_out[11][13] = accbin_in[0][11][13] + accbin_in[1][11][13] + accbin_in[2][11][13] + accbin_in[3][11][13] + accbin_in[4][11][13];
assign sum_out[11][14] = accbin_in[0][11][14] + accbin_in[1][11][14] + accbin_in[2][11][14] + accbin_in[3][11][14] + accbin_in[4][11][14];
assign sum_out[11][15] = accbin_in[0][11][15] + accbin_in[1][11][15] + accbin_in[2][11][15] + accbin_in[3][11][15] + accbin_in[4][11][15];
assign sum_out[11][16] = accbin_in[0][11][16] + accbin_in[1][11][16] + accbin_in[2][11][16] + accbin_in[3][11][16] + accbin_in[4][11][16];
assign sum_out[11][17] = accbin_in[0][11][17] + accbin_in[1][11][17] + accbin_in[2][11][17] + accbin_in[3][11][17] + accbin_in[4][11][17];
assign sum_out[11][18] = accbin_in[0][11][18] + accbin_in[1][11][18] + accbin_in[2][11][18] + accbin_in[3][11][18] + accbin_in[4][11][18];
assign sum_out[11][19] = accbin_in[0][11][19] + accbin_in[1][11][19] + accbin_in[2][11][19] + accbin_in[3][11][19] + accbin_in[4][11][19];
assign sum_out[11][20] = accbin_in[0][11][20] + accbin_in[1][11][20] + accbin_in[2][11][20] + accbin_in[3][11][20] + accbin_in[4][11][20];
assign sum_out[11][21] = accbin_in[0][11][21] + accbin_in[1][11][21] + accbin_in[2][11][21] + accbin_in[3][11][21] + accbin_in[4][11][21];
assign sum_out[11][22] = accbin_in[0][11][22] + accbin_in[1][11][22] + accbin_in[2][11][22] + accbin_in[3][11][22] + accbin_in[4][11][22];
assign sum_out[11][23] = accbin_in[0][11][23] + accbin_in[1][11][23] + accbin_in[2][11][23] + accbin_in[3][11][23] + accbin_in[4][11][23];
assign sum_out[12][0] = accbin_in[0][12][0] + accbin_in[1][12][0] + accbin_in[2][12][0] + accbin_in[3][12][0] + accbin_in[4][12][0];
assign sum_out[12][1] = accbin_in[0][12][1] + accbin_in[1][12][1] + accbin_in[2][12][1] + accbin_in[3][12][1] + accbin_in[4][12][1];
assign sum_out[12][2] = accbin_in[0][12][2] + accbin_in[1][12][2] + accbin_in[2][12][2] + accbin_in[3][12][2] + accbin_in[4][12][2];
assign sum_out[12][3] = accbin_in[0][12][3] + accbin_in[1][12][3] + accbin_in[2][12][3] + accbin_in[3][12][3] + accbin_in[4][12][3];
assign sum_out[12][4] = accbin_in[0][12][4] + accbin_in[1][12][4] + accbin_in[2][12][4] + accbin_in[3][12][4] + accbin_in[4][12][4];
assign sum_out[12][5] = accbin_in[0][12][5] + accbin_in[1][12][5] + accbin_in[2][12][5] + accbin_in[3][12][5] + accbin_in[4][12][5];
assign sum_out[12][6] = accbin_in[0][12][6] + accbin_in[1][12][6] + accbin_in[2][12][6] + accbin_in[3][12][6] + accbin_in[4][12][6];
assign sum_out[12][7] = accbin_in[0][12][7] + accbin_in[1][12][7] + accbin_in[2][12][7] + accbin_in[3][12][7] + accbin_in[4][12][7];
assign sum_out[12][8] = accbin_in[0][12][8] + accbin_in[1][12][8] + accbin_in[2][12][8] + accbin_in[3][12][8] + accbin_in[4][12][8];
assign sum_out[12][9] = accbin_in[0][12][9] + accbin_in[1][12][9] + accbin_in[2][12][9] + accbin_in[3][12][9] + accbin_in[4][12][9];
assign sum_out[12][10] = accbin_in[0][12][10] + accbin_in[1][12][10] + accbin_in[2][12][10] + accbin_in[3][12][10] + accbin_in[4][12][10];
assign sum_out[12][11] = accbin_in[0][12][11] + accbin_in[1][12][11] + accbin_in[2][12][11] + accbin_in[3][12][11] + accbin_in[4][12][11];
assign sum_out[12][12] = accbin_in[0][12][12] + accbin_in[1][12][12] + accbin_in[2][12][12] + accbin_in[3][12][12] + accbin_in[4][12][12];
assign sum_out[12][13] = accbin_in[0][12][13] + accbin_in[1][12][13] + accbin_in[2][12][13] + accbin_in[3][12][13] + accbin_in[4][12][13];
assign sum_out[12][14] = accbin_in[0][12][14] + accbin_in[1][12][14] + accbin_in[2][12][14] + accbin_in[3][12][14] + accbin_in[4][12][14];
assign sum_out[12][15] = accbin_in[0][12][15] + accbin_in[1][12][15] + accbin_in[2][12][15] + accbin_in[3][12][15] + accbin_in[4][12][15];
assign sum_out[12][16] = accbin_in[0][12][16] + accbin_in[1][12][16] + accbin_in[2][12][16] + accbin_in[3][12][16] + accbin_in[4][12][16];
assign sum_out[12][17] = accbin_in[0][12][17] + accbin_in[1][12][17] + accbin_in[2][12][17] + accbin_in[3][12][17] + accbin_in[4][12][17];
assign sum_out[12][18] = accbin_in[0][12][18] + accbin_in[1][12][18] + accbin_in[2][12][18] + accbin_in[3][12][18] + accbin_in[4][12][18];
assign sum_out[12][19] = accbin_in[0][12][19] + accbin_in[1][12][19] + accbin_in[2][12][19] + accbin_in[3][12][19] + accbin_in[4][12][19];
assign sum_out[12][20] = accbin_in[0][12][20] + accbin_in[1][12][20] + accbin_in[2][12][20] + accbin_in[3][12][20] + accbin_in[4][12][20];
assign sum_out[12][21] = accbin_in[0][12][21] + accbin_in[1][12][21] + accbin_in[2][12][21] + accbin_in[3][12][21] + accbin_in[4][12][21];
assign sum_out[12][22] = accbin_in[0][12][22] + accbin_in[1][12][22] + accbin_in[2][12][22] + accbin_in[3][12][22] + accbin_in[4][12][22];
assign sum_out[12][23] = accbin_in[0][12][23] + accbin_in[1][12][23] + accbin_in[2][12][23] + accbin_in[3][12][23] + accbin_in[4][12][23];
assign sum_out[13][0] = accbin_in[0][13][0] + accbin_in[1][13][0] + accbin_in[2][13][0] + accbin_in[3][13][0] + accbin_in[4][13][0];
assign sum_out[13][1] = accbin_in[0][13][1] + accbin_in[1][13][1] + accbin_in[2][13][1] + accbin_in[3][13][1] + accbin_in[4][13][1];
assign sum_out[13][2] = accbin_in[0][13][2] + accbin_in[1][13][2] + accbin_in[2][13][2] + accbin_in[3][13][2] + accbin_in[4][13][2];
assign sum_out[13][3] = accbin_in[0][13][3] + accbin_in[1][13][3] + accbin_in[2][13][3] + accbin_in[3][13][3] + accbin_in[4][13][3];
assign sum_out[13][4] = accbin_in[0][13][4] + accbin_in[1][13][4] + accbin_in[2][13][4] + accbin_in[3][13][4] + accbin_in[4][13][4];
assign sum_out[13][5] = accbin_in[0][13][5] + accbin_in[1][13][5] + accbin_in[2][13][5] + accbin_in[3][13][5] + accbin_in[4][13][5];
assign sum_out[13][6] = accbin_in[0][13][6] + accbin_in[1][13][6] + accbin_in[2][13][6] + accbin_in[3][13][6] + accbin_in[4][13][6];
assign sum_out[13][7] = accbin_in[0][13][7] + accbin_in[1][13][7] + accbin_in[2][13][7] + accbin_in[3][13][7] + accbin_in[4][13][7];
assign sum_out[13][8] = accbin_in[0][13][8] + accbin_in[1][13][8] + accbin_in[2][13][8] + accbin_in[3][13][8] + accbin_in[4][13][8];
assign sum_out[13][9] = accbin_in[0][13][9] + accbin_in[1][13][9] + accbin_in[2][13][9] + accbin_in[3][13][9] + accbin_in[4][13][9];
assign sum_out[13][10] = accbin_in[0][13][10] + accbin_in[1][13][10] + accbin_in[2][13][10] + accbin_in[3][13][10] + accbin_in[4][13][10];
assign sum_out[13][11] = accbin_in[0][13][11] + accbin_in[1][13][11] + accbin_in[2][13][11] + accbin_in[3][13][11] + accbin_in[4][13][11];
assign sum_out[13][12] = accbin_in[0][13][12] + accbin_in[1][13][12] + accbin_in[2][13][12] + accbin_in[3][13][12] + accbin_in[4][13][12];
assign sum_out[13][13] = accbin_in[0][13][13] + accbin_in[1][13][13] + accbin_in[2][13][13] + accbin_in[3][13][13] + accbin_in[4][13][13];
assign sum_out[13][14] = accbin_in[0][13][14] + accbin_in[1][13][14] + accbin_in[2][13][14] + accbin_in[3][13][14] + accbin_in[4][13][14];
assign sum_out[13][15] = accbin_in[0][13][15] + accbin_in[1][13][15] + accbin_in[2][13][15] + accbin_in[3][13][15] + accbin_in[4][13][15];
assign sum_out[13][16] = accbin_in[0][13][16] + accbin_in[1][13][16] + accbin_in[2][13][16] + accbin_in[3][13][16] + accbin_in[4][13][16];
assign sum_out[13][17] = accbin_in[0][13][17] + accbin_in[1][13][17] + accbin_in[2][13][17] + accbin_in[3][13][17] + accbin_in[4][13][17];
assign sum_out[13][18] = accbin_in[0][13][18] + accbin_in[1][13][18] + accbin_in[2][13][18] + accbin_in[3][13][18] + accbin_in[4][13][18];
assign sum_out[13][19] = accbin_in[0][13][19] + accbin_in[1][13][19] + accbin_in[2][13][19] + accbin_in[3][13][19] + accbin_in[4][13][19];
assign sum_out[13][20] = accbin_in[0][13][20] + accbin_in[1][13][20] + accbin_in[2][13][20] + accbin_in[3][13][20] + accbin_in[4][13][20];
assign sum_out[13][21] = accbin_in[0][13][21] + accbin_in[1][13][21] + accbin_in[2][13][21] + accbin_in[3][13][21] + accbin_in[4][13][21];
assign sum_out[13][22] = accbin_in[0][13][22] + accbin_in[1][13][22] + accbin_in[2][13][22] + accbin_in[3][13][22] + accbin_in[4][13][22];
assign sum_out[13][23] = accbin_in[0][13][23] + accbin_in[1][13][23] + accbin_in[2][13][23] + accbin_in[3][13][23] + accbin_in[4][13][23];
assign sum_out[14][0] = accbin_in[0][14][0] + accbin_in[1][14][0] + accbin_in[2][14][0] + accbin_in[3][14][0] + accbin_in[4][14][0];
assign sum_out[14][1] = accbin_in[0][14][1] + accbin_in[1][14][1] + accbin_in[2][14][1] + accbin_in[3][14][1] + accbin_in[4][14][1];
assign sum_out[14][2] = accbin_in[0][14][2] + accbin_in[1][14][2] + accbin_in[2][14][2] + accbin_in[3][14][2] + accbin_in[4][14][2];
assign sum_out[14][3] = accbin_in[0][14][3] + accbin_in[1][14][3] + accbin_in[2][14][3] + accbin_in[3][14][3] + accbin_in[4][14][3];
assign sum_out[14][4] = accbin_in[0][14][4] + accbin_in[1][14][4] + accbin_in[2][14][4] + accbin_in[3][14][4] + accbin_in[4][14][4];
assign sum_out[14][5] = accbin_in[0][14][5] + accbin_in[1][14][5] + accbin_in[2][14][5] + accbin_in[3][14][5] + accbin_in[4][14][5];
assign sum_out[14][6] = accbin_in[0][14][6] + accbin_in[1][14][6] + accbin_in[2][14][6] + accbin_in[3][14][6] + accbin_in[4][14][6];
assign sum_out[14][7] = accbin_in[0][14][7] + accbin_in[1][14][7] + accbin_in[2][14][7] + accbin_in[3][14][7] + accbin_in[4][14][7];
assign sum_out[14][8] = accbin_in[0][14][8] + accbin_in[1][14][8] + accbin_in[2][14][8] + accbin_in[3][14][8] + accbin_in[4][14][8];
assign sum_out[14][9] = accbin_in[0][14][9] + accbin_in[1][14][9] + accbin_in[2][14][9] + accbin_in[3][14][9] + accbin_in[4][14][9];
assign sum_out[14][10] = accbin_in[0][14][10] + accbin_in[1][14][10] + accbin_in[2][14][10] + accbin_in[3][14][10] + accbin_in[4][14][10];
assign sum_out[14][11] = accbin_in[0][14][11] + accbin_in[1][14][11] + accbin_in[2][14][11] + accbin_in[3][14][11] + accbin_in[4][14][11];
assign sum_out[14][12] = accbin_in[0][14][12] + accbin_in[1][14][12] + accbin_in[2][14][12] + accbin_in[3][14][12] + accbin_in[4][14][12];
assign sum_out[14][13] = accbin_in[0][14][13] + accbin_in[1][14][13] + accbin_in[2][14][13] + accbin_in[3][14][13] + accbin_in[4][14][13];
assign sum_out[14][14] = accbin_in[0][14][14] + accbin_in[1][14][14] + accbin_in[2][14][14] + accbin_in[3][14][14] + accbin_in[4][14][14];
assign sum_out[14][15] = accbin_in[0][14][15] + accbin_in[1][14][15] + accbin_in[2][14][15] + accbin_in[3][14][15] + accbin_in[4][14][15];
assign sum_out[14][16] = accbin_in[0][14][16] + accbin_in[1][14][16] + accbin_in[2][14][16] + accbin_in[3][14][16] + accbin_in[4][14][16];
assign sum_out[14][17] = accbin_in[0][14][17] + accbin_in[1][14][17] + accbin_in[2][14][17] + accbin_in[3][14][17] + accbin_in[4][14][17];
assign sum_out[14][18] = accbin_in[0][14][18] + accbin_in[1][14][18] + accbin_in[2][14][18] + accbin_in[3][14][18] + accbin_in[4][14][18];
assign sum_out[14][19] = accbin_in[0][14][19] + accbin_in[1][14][19] + accbin_in[2][14][19] + accbin_in[3][14][19] + accbin_in[4][14][19];
assign sum_out[14][20] = accbin_in[0][14][20] + accbin_in[1][14][20] + accbin_in[2][14][20] + accbin_in[3][14][20] + accbin_in[4][14][20];
assign sum_out[14][21] = accbin_in[0][14][21] + accbin_in[1][14][21] + accbin_in[2][14][21] + accbin_in[3][14][21] + accbin_in[4][14][21];
assign sum_out[14][22] = accbin_in[0][14][22] + accbin_in[1][14][22] + accbin_in[2][14][22] + accbin_in[3][14][22] + accbin_in[4][14][22];
assign sum_out[14][23] = accbin_in[0][14][23] + accbin_in[1][14][23] + accbin_in[2][14][23] + accbin_in[3][14][23] + accbin_in[4][14][23];
assign sum_out[15][0] = accbin_in[0][15][0] + accbin_in[1][15][0] + accbin_in[2][15][0] + accbin_in[3][15][0] + accbin_in[4][15][0];
assign sum_out[15][1] = accbin_in[0][15][1] + accbin_in[1][15][1] + accbin_in[2][15][1] + accbin_in[3][15][1] + accbin_in[4][15][1];
assign sum_out[15][2] = accbin_in[0][15][2] + accbin_in[1][15][2] + accbin_in[2][15][2] + accbin_in[3][15][2] + accbin_in[4][15][2];
assign sum_out[15][3] = accbin_in[0][15][3] + accbin_in[1][15][3] + accbin_in[2][15][3] + accbin_in[3][15][3] + accbin_in[4][15][3];
assign sum_out[15][4] = accbin_in[0][15][4] + accbin_in[1][15][4] + accbin_in[2][15][4] + accbin_in[3][15][4] + accbin_in[4][15][4];
assign sum_out[15][5] = accbin_in[0][15][5] + accbin_in[1][15][5] + accbin_in[2][15][5] + accbin_in[3][15][5] + accbin_in[4][15][5];
assign sum_out[15][6] = accbin_in[0][15][6] + accbin_in[1][15][6] + accbin_in[2][15][6] + accbin_in[3][15][6] + accbin_in[4][15][6];
assign sum_out[15][7] = accbin_in[0][15][7] + accbin_in[1][15][7] + accbin_in[2][15][7] + accbin_in[3][15][7] + accbin_in[4][15][7];
assign sum_out[15][8] = accbin_in[0][15][8] + accbin_in[1][15][8] + accbin_in[2][15][8] + accbin_in[3][15][8] + accbin_in[4][15][8];
assign sum_out[15][9] = accbin_in[0][15][9] + accbin_in[1][15][9] + accbin_in[2][15][9] + accbin_in[3][15][9] + accbin_in[4][15][9];
assign sum_out[15][10] = accbin_in[0][15][10] + accbin_in[1][15][10] + accbin_in[2][15][10] + accbin_in[3][15][10] + accbin_in[4][15][10];
assign sum_out[15][11] = accbin_in[0][15][11] + accbin_in[1][15][11] + accbin_in[2][15][11] + accbin_in[3][15][11] + accbin_in[4][15][11];
assign sum_out[15][12] = accbin_in[0][15][12] + accbin_in[1][15][12] + accbin_in[2][15][12] + accbin_in[3][15][12] + accbin_in[4][15][12];
assign sum_out[15][13] = accbin_in[0][15][13] + accbin_in[1][15][13] + accbin_in[2][15][13] + accbin_in[3][15][13] + accbin_in[4][15][13];
assign sum_out[15][14] = accbin_in[0][15][14] + accbin_in[1][15][14] + accbin_in[2][15][14] + accbin_in[3][15][14] + accbin_in[4][15][14];
assign sum_out[15][15] = accbin_in[0][15][15] + accbin_in[1][15][15] + accbin_in[2][15][15] + accbin_in[3][15][15] + accbin_in[4][15][15];
assign sum_out[15][16] = accbin_in[0][15][16] + accbin_in[1][15][16] + accbin_in[2][15][16] + accbin_in[3][15][16] + accbin_in[4][15][16];
assign sum_out[15][17] = accbin_in[0][15][17] + accbin_in[1][15][17] + accbin_in[2][15][17] + accbin_in[3][15][17] + accbin_in[4][15][17];
assign sum_out[15][18] = accbin_in[0][15][18] + accbin_in[1][15][18] + accbin_in[2][15][18] + accbin_in[3][15][18] + accbin_in[4][15][18];
assign sum_out[15][19] = accbin_in[0][15][19] + accbin_in[1][15][19] + accbin_in[2][15][19] + accbin_in[3][15][19] + accbin_in[4][15][19];
assign sum_out[15][20] = accbin_in[0][15][20] + accbin_in[1][15][20] + accbin_in[2][15][20] + accbin_in[3][15][20] + accbin_in[4][15][20];
assign sum_out[15][21] = accbin_in[0][15][21] + accbin_in[1][15][21] + accbin_in[2][15][21] + accbin_in[3][15][21] + accbin_in[4][15][21];
assign sum_out[15][22] = accbin_in[0][15][22] + accbin_in[1][15][22] + accbin_in[2][15][22] + accbin_in[3][15][22] + accbin_in[4][15][22];
assign sum_out[15][23] = accbin_in[0][15][23] + accbin_in[1][15][23] + accbin_in[2][15][23] + accbin_in[3][15][23] + accbin_in[4][15][23];
assign sum_out[16][0] = accbin_in[0][16][0] + accbin_in[1][16][0] + accbin_in[2][16][0] + accbin_in[3][16][0] + accbin_in[4][16][0];
assign sum_out[16][1] = accbin_in[0][16][1] + accbin_in[1][16][1] + accbin_in[2][16][1] + accbin_in[3][16][1] + accbin_in[4][16][1];
assign sum_out[16][2] = accbin_in[0][16][2] + accbin_in[1][16][2] + accbin_in[2][16][2] + accbin_in[3][16][2] + accbin_in[4][16][2];
assign sum_out[16][3] = accbin_in[0][16][3] + accbin_in[1][16][3] + accbin_in[2][16][3] + accbin_in[3][16][3] + accbin_in[4][16][3];
assign sum_out[16][4] = accbin_in[0][16][4] + accbin_in[1][16][4] + accbin_in[2][16][4] + accbin_in[3][16][4] + accbin_in[4][16][4];
assign sum_out[16][5] = accbin_in[0][16][5] + accbin_in[1][16][5] + accbin_in[2][16][5] + accbin_in[3][16][5] + accbin_in[4][16][5];
assign sum_out[16][6] = accbin_in[0][16][6] + accbin_in[1][16][6] + accbin_in[2][16][6] + accbin_in[3][16][6] + accbin_in[4][16][6];
assign sum_out[16][7] = accbin_in[0][16][7] + accbin_in[1][16][7] + accbin_in[2][16][7] + accbin_in[3][16][7] + accbin_in[4][16][7];
assign sum_out[16][8] = accbin_in[0][16][8] + accbin_in[1][16][8] + accbin_in[2][16][8] + accbin_in[3][16][8] + accbin_in[4][16][8];
assign sum_out[16][9] = accbin_in[0][16][9] + accbin_in[1][16][9] + accbin_in[2][16][9] + accbin_in[3][16][9] + accbin_in[4][16][9];
assign sum_out[16][10] = accbin_in[0][16][10] + accbin_in[1][16][10] + accbin_in[2][16][10] + accbin_in[3][16][10] + accbin_in[4][16][10];
assign sum_out[16][11] = accbin_in[0][16][11] + accbin_in[1][16][11] + accbin_in[2][16][11] + accbin_in[3][16][11] + accbin_in[4][16][11];
assign sum_out[16][12] = accbin_in[0][16][12] + accbin_in[1][16][12] + accbin_in[2][16][12] + accbin_in[3][16][12] + accbin_in[4][16][12];
assign sum_out[16][13] = accbin_in[0][16][13] + accbin_in[1][16][13] + accbin_in[2][16][13] + accbin_in[3][16][13] + accbin_in[4][16][13];
assign sum_out[16][14] = accbin_in[0][16][14] + accbin_in[1][16][14] + accbin_in[2][16][14] + accbin_in[3][16][14] + accbin_in[4][16][14];
assign sum_out[16][15] = accbin_in[0][16][15] + accbin_in[1][16][15] + accbin_in[2][16][15] + accbin_in[3][16][15] + accbin_in[4][16][15];
assign sum_out[16][16] = accbin_in[0][16][16] + accbin_in[1][16][16] + accbin_in[2][16][16] + accbin_in[3][16][16] + accbin_in[4][16][16];
assign sum_out[16][17] = accbin_in[0][16][17] + accbin_in[1][16][17] + accbin_in[2][16][17] + accbin_in[3][16][17] + accbin_in[4][16][17];
assign sum_out[16][18] = accbin_in[0][16][18] + accbin_in[1][16][18] + accbin_in[2][16][18] + accbin_in[3][16][18] + accbin_in[4][16][18];
assign sum_out[16][19] = accbin_in[0][16][19] + accbin_in[1][16][19] + accbin_in[2][16][19] + accbin_in[3][16][19] + accbin_in[4][16][19];
assign sum_out[16][20] = accbin_in[0][16][20] + accbin_in[1][16][20] + accbin_in[2][16][20] + accbin_in[3][16][20] + accbin_in[4][16][20];
assign sum_out[16][21] = accbin_in[0][16][21] + accbin_in[1][16][21] + accbin_in[2][16][21] + accbin_in[3][16][21] + accbin_in[4][16][21];
assign sum_out[16][22] = accbin_in[0][16][22] + accbin_in[1][16][22] + accbin_in[2][16][22] + accbin_in[3][16][22] + accbin_in[4][16][22];
assign sum_out[16][23] = accbin_in[0][16][23] + accbin_in[1][16][23] + accbin_in[2][16][23] + accbin_in[3][16][23] + accbin_in[4][16][23];
assign sum_out[17][0] = accbin_in[0][17][0] + accbin_in[1][17][0] + accbin_in[2][17][0] + accbin_in[3][17][0] + accbin_in[4][17][0];
assign sum_out[17][1] = accbin_in[0][17][1] + accbin_in[1][17][1] + accbin_in[2][17][1] + accbin_in[3][17][1] + accbin_in[4][17][1];
assign sum_out[17][2] = accbin_in[0][17][2] + accbin_in[1][17][2] + accbin_in[2][17][2] + accbin_in[3][17][2] + accbin_in[4][17][2];
assign sum_out[17][3] = accbin_in[0][17][3] + accbin_in[1][17][3] + accbin_in[2][17][3] + accbin_in[3][17][3] + accbin_in[4][17][3];
assign sum_out[17][4] = accbin_in[0][17][4] + accbin_in[1][17][4] + accbin_in[2][17][4] + accbin_in[3][17][4] + accbin_in[4][17][4];
assign sum_out[17][5] = accbin_in[0][17][5] + accbin_in[1][17][5] + accbin_in[2][17][5] + accbin_in[3][17][5] + accbin_in[4][17][5];
assign sum_out[17][6] = accbin_in[0][17][6] + accbin_in[1][17][6] + accbin_in[2][17][6] + accbin_in[3][17][6] + accbin_in[4][17][6];
assign sum_out[17][7] = accbin_in[0][17][7] + accbin_in[1][17][7] + accbin_in[2][17][7] + accbin_in[3][17][7] + accbin_in[4][17][7];
assign sum_out[17][8] = accbin_in[0][17][8] + accbin_in[1][17][8] + accbin_in[2][17][8] + accbin_in[3][17][8] + accbin_in[4][17][8];
assign sum_out[17][9] = accbin_in[0][17][9] + accbin_in[1][17][9] + accbin_in[2][17][9] + accbin_in[3][17][9] + accbin_in[4][17][9];
assign sum_out[17][10] = accbin_in[0][17][10] + accbin_in[1][17][10] + accbin_in[2][17][10] + accbin_in[3][17][10] + accbin_in[4][17][10];
assign sum_out[17][11] = accbin_in[0][17][11] + accbin_in[1][17][11] + accbin_in[2][17][11] + accbin_in[3][17][11] + accbin_in[4][17][11];
assign sum_out[17][12] = accbin_in[0][17][12] + accbin_in[1][17][12] + accbin_in[2][17][12] + accbin_in[3][17][12] + accbin_in[4][17][12];
assign sum_out[17][13] = accbin_in[0][17][13] + accbin_in[1][17][13] + accbin_in[2][17][13] + accbin_in[3][17][13] + accbin_in[4][17][13];
assign sum_out[17][14] = accbin_in[0][17][14] + accbin_in[1][17][14] + accbin_in[2][17][14] + accbin_in[3][17][14] + accbin_in[4][17][14];
assign sum_out[17][15] = accbin_in[0][17][15] + accbin_in[1][17][15] + accbin_in[2][17][15] + accbin_in[3][17][15] + accbin_in[4][17][15];
assign sum_out[17][16] = accbin_in[0][17][16] + accbin_in[1][17][16] + accbin_in[2][17][16] + accbin_in[3][17][16] + accbin_in[4][17][16];
assign sum_out[17][17] = accbin_in[0][17][17] + accbin_in[1][17][17] + accbin_in[2][17][17] + accbin_in[3][17][17] + accbin_in[4][17][17];
assign sum_out[17][18] = accbin_in[0][17][18] + accbin_in[1][17][18] + accbin_in[2][17][18] + accbin_in[3][17][18] + accbin_in[4][17][18];
assign sum_out[17][19] = accbin_in[0][17][19] + accbin_in[1][17][19] + accbin_in[2][17][19] + accbin_in[3][17][19] + accbin_in[4][17][19];
assign sum_out[17][20] = accbin_in[0][17][20] + accbin_in[1][17][20] + accbin_in[2][17][20] + accbin_in[3][17][20] + accbin_in[4][17][20];
assign sum_out[17][21] = accbin_in[0][17][21] + accbin_in[1][17][21] + accbin_in[2][17][21] + accbin_in[3][17][21] + accbin_in[4][17][21];
assign sum_out[17][22] = accbin_in[0][17][22] + accbin_in[1][17][22] + accbin_in[2][17][22] + accbin_in[3][17][22] + accbin_in[4][17][22];
assign sum_out[17][23] = accbin_in[0][17][23] + accbin_in[1][17][23] + accbin_in[2][17][23] + accbin_in[3][17][23] + accbin_in[4][17][23];
assign sum_out[18][0] = accbin_in[0][18][0] + accbin_in[1][18][0] + accbin_in[2][18][0] + accbin_in[3][18][0] + accbin_in[4][18][0];
assign sum_out[18][1] = accbin_in[0][18][1] + accbin_in[1][18][1] + accbin_in[2][18][1] + accbin_in[3][18][1] + accbin_in[4][18][1];
assign sum_out[18][2] = accbin_in[0][18][2] + accbin_in[1][18][2] + accbin_in[2][18][2] + accbin_in[3][18][2] + accbin_in[4][18][2];
assign sum_out[18][3] = accbin_in[0][18][3] + accbin_in[1][18][3] + accbin_in[2][18][3] + accbin_in[3][18][3] + accbin_in[4][18][3];
assign sum_out[18][4] = accbin_in[0][18][4] + accbin_in[1][18][4] + accbin_in[2][18][4] + accbin_in[3][18][4] + accbin_in[4][18][4];
assign sum_out[18][5] = accbin_in[0][18][5] + accbin_in[1][18][5] + accbin_in[2][18][5] + accbin_in[3][18][5] + accbin_in[4][18][5];
assign sum_out[18][6] = accbin_in[0][18][6] + accbin_in[1][18][6] + accbin_in[2][18][6] + accbin_in[3][18][6] + accbin_in[4][18][6];
assign sum_out[18][7] = accbin_in[0][18][7] + accbin_in[1][18][7] + accbin_in[2][18][7] + accbin_in[3][18][7] + accbin_in[4][18][7];
assign sum_out[18][8] = accbin_in[0][18][8] + accbin_in[1][18][8] + accbin_in[2][18][8] + accbin_in[3][18][8] + accbin_in[4][18][8];
assign sum_out[18][9] = accbin_in[0][18][9] + accbin_in[1][18][9] + accbin_in[2][18][9] + accbin_in[3][18][9] + accbin_in[4][18][9];
assign sum_out[18][10] = accbin_in[0][18][10] + accbin_in[1][18][10] + accbin_in[2][18][10] + accbin_in[3][18][10] + accbin_in[4][18][10];
assign sum_out[18][11] = accbin_in[0][18][11] + accbin_in[1][18][11] + accbin_in[2][18][11] + accbin_in[3][18][11] + accbin_in[4][18][11];
assign sum_out[18][12] = accbin_in[0][18][12] + accbin_in[1][18][12] + accbin_in[2][18][12] + accbin_in[3][18][12] + accbin_in[4][18][12];
assign sum_out[18][13] = accbin_in[0][18][13] + accbin_in[1][18][13] + accbin_in[2][18][13] + accbin_in[3][18][13] + accbin_in[4][18][13];
assign sum_out[18][14] = accbin_in[0][18][14] + accbin_in[1][18][14] + accbin_in[2][18][14] + accbin_in[3][18][14] + accbin_in[4][18][14];
assign sum_out[18][15] = accbin_in[0][18][15] + accbin_in[1][18][15] + accbin_in[2][18][15] + accbin_in[3][18][15] + accbin_in[4][18][15];
assign sum_out[18][16] = accbin_in[0][18][16] + accbin_in[1][18][16] + accbin_in[2][18][16] + accbin_in[3][18][16] + accbin_in[4][18][16];
assign sum_out[18][17] = accbin_in[0][18][17] + accbin_in[1][18][17] + accbin_in[2][18][17] + accbin_in[3][18][17] + accbin_in[4][18][17];
assign sum_out[18][18] = accbin_in[0][18][18] + accbin_in[1][18][18] + accbin_in[2][18][18] + accbin_in[3][18][18] + accbin_in[4][18][18];
assign sum_out[18][19] = accbin_in[0][18][19] + accbin_in[1][18][19] + accbin_in[2][18][19] + accbin_in[3][18][19] + accbin_in[4][18][19];
assign sum_out[18][20] = accbin_in[0][18][20] + accbin_in[1][18][20] + accbin_in[2][18][20] + accbin_in[3][18][20] + accbin_in[4][18][20];
assign sum_out[18][21] = accbin_in[0][18][21] + accbin_in[1][18][21] + accbin_in[2][18][21] + accbin_in[3][18][21] + accbin_in[4][18][21];
assign sum_out[18][22] = accbin_in[0][18][22] + accbin_in[1][18][22] + accbin_in[2][18][22] + accbin_in[3][18][22] + accbin_in[4][18][22];
assign sum_out[18][23] = accbin_in[0][18][23] + accbin_in[1][18][23] + accbin_in[2][18][23] + accbin_in[3][18][23] + accbin_in[4][18][23];
assign sum_out[19][0] = accbin_in[0][19][0] + accbin_in[1][19][0] + accbin_in[2][19][0] + accbin_in[3][19][0] + accbin_in[4][19][0];
assign sum_out[19][1] = accbin_in[0][19][1] + accbin_in[1][19][1] + accbin_in[2][19][1] + accbin_in[3][19][1] + accbin_in[4][19][1];
assign sum_out[19][2] = accbin_in[0][19][2] + accbin_in[1][19][2] + accbin_in[2][19][2] + accbin_in[3][19][2] + accbin_in[4][19][2];
assign sum_out[19][3] = accbin_in[0][19][3] + accbin_in[1][19][3] + accbin_in[2][19][3] + accbin_in[3][19][3] + accbin_in[4][19][3];
assign sum_out[19][4] = accbin_in[0][19][4] + accbin_in[1][19][4] + accbin_in[2][19][4] + accbin_in[3][19][4] + accbin_in[4][19][4];
assign sum_out[19][5] = accbin_in[0][19][5] + accbin_in[1][19][5] + accbin_in[2][19][5] + accbin_in[3][19][5] + accbin_in[4][19][5];
assign sum_out[19][6] = accbin_in[0][19][6] + accbin_in[1][19][6] + accbin_in[2][19][6] + accbin_in[3][19][6] + accbin_in[4][19][6];
assign sum_out[19][7] = accbin_in[0][19][7] + accbin_in[1][19][7] + accbin_in[2][19][7] + accbin_in[3][19][7] + accbin_in[4][19][7];
assign sum_out[19][8] = accbin_in[0][19][8] + accbin_in[1][19][8] + accbin_in[2][19][8] + accbin_in[3][19][8] + accbin_in[4][19][8];
assign sum_out[19][9] = accbin_in[0][19][9] + accbin_in[1][19][9] + accbin_in[2][19][9] + accbin_in[3][19][9] + accbin_in[4][19][9];
assign sum_out[19][10] = accbin_in[0][19][10] + accbin_in[1][19][10] + accbin_in[2][19][10] + accbin_in[3][19][10] + accbin_in[4][19][10];
assign sum_out[19][11] = accbin_in[0][19][11] + accbin_in[1][19][11] + accbin_in[2][19][11] + accbin_in[3][19][11] + accbin_in[4][19][11];
assign sum_out[19][12] = accbin_in[0][19][12] + accbin_in[1][19][12] + accbin_in[2][19][12] + accbin_in[3][19][12] + accbin_in[4][19][12];
assign sum_out[19][13] = accbin_in[0][19][13] + accbin_in[1][19][13] + accbin_in[2][19][13] + accbin_in[3][19][13] + accbin_in[4][19][13];
assign sum_out[19][14] = accbin_in[0][19][14] + accbin_in[1][19][14] + accbin_in[2][19][14] + accbin_in[3][19][14] + accbin_in[4][19][14];
assign sum_out[19][15] = accbin_in[0][19][15] + accbin_in[1][19][15] + accbin_in[2][19][15] + accbin_in[3][19][15] + accbin_in[4][19][15];
assign sum_out[19][16] = accbin_in[0][19][16] + accbin_in[1][19][16] + accbin_in[2][19][16] + accbin_in[3][19][16] + accbin_in[4][19][16];
assign sum_out[19][17] = accbin_in[0][19][17] + accbin_in[1][19][17] + accbin_in[2][19][17] + accbin_in[3][19][17] + accbin_in[4][19][17];
assign sum_out[19][18] = accbin_in[0][19][18] + accbin_in[1][19][18] + accbin_in[2][19][18] + accbin_in[3][19][18] + accbin_in[4][19][18];
assign sum_out[19][19] = accbin_in[0][19][19] + accbin_in[1][19][19] + accbin_in[2][19][19] + accbin_in[3][19][19] + accbin_in[4][19][19];
assign sum_out[19][20] = accbin_in[0][19][20] + accbin_in[1][19][20] + accbin_in[2][19][20] + accbin_in[3][19][20] + accbin_in[4][19][20];
assign sum_out[19][21] = accbin_in[0][19][21] + accbin_in[1][19][21] + accbin_in[2][19][21] + accbin_in[3][19][21] + accbin_in[4][19][21];
assign sum_out[19][22] = accbin_in[0][19][22] + accbin_in[1][19][22] + accbin_in[2][19][22] + accbin_in[3][19][22] + accbin_in[4][19][22];
assign sum_out[19][23] = accbin_in[0][19][23] + accbin_in[1][19][23] + accbin_in[2][19][23] + accbin_in[3][19][23] + accbin_in[4][19][23];
assign sum_out[20][0] = accbin_in[0][20][0] + accbin_in[1][20][0] + accbin_in[2][20][0] + accbin_in[3][20][0] + accbin_in[4][20][0];
assign sum_out[20][1] = accbin_in[0][20][1] + accbin_in[1][20][1] + accbin_in[2][20][1] + accbin_in[3][20][1] + accbin_in[4][20][1];
assign sum_out[20][2] = accbin_in[0][20][2] + accbin_in[1][20][2] + accbin_in[2][20][2] + accbin_in[3][20][2] + accbin_in[4][20][2];
assign sum_out[20][3] = accbin_in[0][20][3] + accbin_in[1][20][3] + accbin_in[2][20][3] + accbin_in[3][20][3] + accbin_in[4][20][3];
assign sum_out[20][4] = accbin_in[0][20][4] + accbin_in[1][20][4] + accbin_in[2][20][4] + accbin_in[3][20][4] + accbin_in[4][20][4];
assign sum_out[20][5] = accbin_in[0][20][5] + accbin_in[1][20][5] + accbin_in[2][20][5] + accbin_in[3][20][5] + accbin_in[4][20][5];
assign sum_out[20][6] = accbin_in[0][20][6] + accbin_in[1][20][6] + accbin_in[2][20][6] + accbin_in[3][20][6] + accbin_in[4][20][6];
assign sum_out[20][7] = accbin_in[0][20][7] + accbin_in[1][20][7] + accbin_in[2][20][7] + accbin_in[3][20][7] + accbin_in[4][20][7];
assign sum_out[20][8] = accbin_in[0][20][8] + accbin_in[1][20][8] + accbin_in[2][20][8] + accbin_in[3][20][8] + accbin_in[4][20][8];
assign sum_out[20][9] = accbin_in[0][20][9] + accbin_in[1][20][9] + accbin_in[2][20][9] + accbin_in[3][20][9] + accbin_in[4][20][9];
assign sum_out[20][10] = accbin_in[0][20][10] + accbin_in[1][20][10] + accbin_in[2][20][10] + accbin_in[3][20][10] + accbin_in[4][20][10];
assign sum_out[20][11] = accbin_in[0][20][11] + accbin_in[1][20][11] + accbin_in[2][20][11] + accbin_in[3][20][11] + accbin_in[4][20][11];
assign sum_out[20][12] = accbin_in[0][20][12] + accbin_in[1][20][12] + accbin_in[2][20][12] + accbin_in[3][20][12] + accbin_in[4][20][12];
assign sum_out[20][13] = accbin_in[0][20][13] + accbin_in[1][20][13] + accbin_in[2][20][13] + accbin_in[3][20][13] + accbin_in[4][20][13];
assign sum_out[20][14] = accbin_in[0][20][14] + accbin_in[1][20][14] + accbin_in[2][20][14] + accbin_in[3][20][14] + accbin_in[4][20][14];
assign sum_out[20][15] = accbin_in[0][20][15] + accbin_in[1][20][15] + accbin_in[2][20][15] + accbin_in[3][20][15] + accbin_in[4][20][15];
assign sum_out[20][16] = accbin_in[0][20][16] + accbin_in[1][20][16] + accbin_in[2][20][16] + accbin_in[3][20][16] + accbin_in[4][20][16];
assign sum_out[20][17] = accbin_in[0][20][17] + accbin_in[1][20][17] + accbin_in[2][20][17] + accbin_in[3][20][17] + accbin_in[4][20][17];
assign sum_out[20][18] = accbin_in[0][20][18] + accbin_in[1][20][18] + accbin_in[2][20][18] + accbin_in[3][20][18] + accbin_in[4][20][18];
assign sum_out[20][19] = accbin_in[0][20][19] + accbin_in[1][20][19] + accbin_in[2][20][19] + accbin_in[3][20][19] + accbin_in[4][20][19];
assign sum_out[20][20] = accbin_in[0][20][20] + accbin_in[1][20][20] + accbin_in[2][20][20] + accbin_in[3][20][20] + accbin_in[4][20][20];
assign sum_out[20][21] = accbin_in[0][20][21] + accbin_in[1][20][21] + accbin_in[2][20][21] + accbin_in[3][20][21] + accbin_in[4][20][21];
assign sum_out[20][22] = accbin_in[0][20][22] + accbin_in[1][20][22] + accbin_in[2][20][22] + accbin_in[3][20][22] + accbin_in[4][20][22];
assign sum_out[20][23] = accbin_in[0][20][23] + accbin_in[1][20][23] + accbin_in[2][20][23] + accbin_in[3][20][23] + accbin_in[4][20][23];
assign sum_out[21][0] = accbin_in[0][21][0] + accbin_in[1][21][0] + accbin_in[2][21][0] + accbin_in[3][21][0] + accbin_in[4][21][0];
assign sum_out[21][1] = accbin_in[0][21][1] + accbin_in[1][21][1] + accbin_in[2][21][1] + accbin_in[3][21][1] + accbin_in[4][21][1];
assign sum_out[21][2] = accbin_in[0][21][2] + accbin_in[1][21][2] + accbin_in[2][21][2] + accbin_in[3][21][2] + accbin_in[4][21][2];
assign sum_out[21][3] = accbin_in[0][21][3] + accbin_in[1][21][3] + accbin_in[2][21][3] + accbin_in[3][21][3] + accbin_in[4][21][3];
assign sum_out[21][4] = accbin_in[0][21][4] + accbin_in[1][21][4] + accbin_in[2][21][4] + accbin_in[3][21][4] + accbin_in[4][21][4];
assign sum_out[21][5] = accbin_in[0][21][5] + accbin_in[1][21][5] + accbin_in[2][21][5] + accbin_in[3][21][5] + accbin_in[4][21][5];
assign sum_out[21][6] = accbin_in[0][21][6] + accbin_in[1][21][6] + accbin_in[2][21][6] + accbin_in[3][21][6] + accbin_in[4][21][6];
assign sum_out[21][7] = accbin_in[0][21][7] + accbin_in[1][21][7] + accbin_in[2][21][7] + accbin_in[3][21][7] + accbin_in[4][21][7];
assign sum_out[21][8] = accbin_in[0][21][8] + accbin_in[1][21][8] + accbin_in[2][21][8] + accbin_in[3][21][8] + accbin_in[4][21][8];
assign sum_out[21][9] = accbin_in[0][21][9] + accbin_in[1][21][9] + accbin_in[2][21][9] + accbin_in[3][21][9] + accbin_in[4][21][9];
assign sum_out[21][10] = accbin_in[0][21][10] + accbin_in[1][21][10] + accbin_in[2][21][10] + accbin_in[3][21][10] + accbin_in[4][21][10];
assign sum_out[21][11] = accbin_in[0][21][11] + accbin_in[1][21][11] + accbin_in[2][21][11] + accbin_in[3][21][11] + accbin_in[4][21][11];
assign sum_out[21][12] = accbin_in[0][21][12] + accbin_in[1][21][12] + accbin_in[2][21][12] + accbin_in[3][21][12] + accbin_in[4][21][12];
assign sum_out[21][13] = accbin_in[0][21][13] + accbin_in[1][21][13] + accbin_in[2][21][13] + accbin_in[3][21][13] + accbin_in[4][21][13];
assign sum_out[21][14] = accbin_in[0][21][14] + accbin_in[1][21][14] + accbin_in[2][21][14] + accbin_in[3][21][14] + accbin_in[4][21][14];
assign sum_out[21][15] = accbin_in[0][21][15] + accbin_in[1][21][15] + accbin_in[2][21][15] + accbin_in[3][21][15] + accbin_in[4][21][15];
assign sum_out[21][16] = accbin_in[0][21][16] + accbin_in[1][21][16] + accbin_in[2][21][16] + accbin_in[3][21][16] + accbin_in[4][21][16];
assign sum_out[21][17] = accbin_in[0][21][17] + accbin_in[1][21][17] + accbin_in[2][21][17] + accbin_in[3][21][17] + accbin_in[4][21][17];
assign sum_out[21][18] = accbin_in[0][21][18] + accbin_in[1][21][18] + accbin_in[2][21][18] + accbin_in[3][21][18] + accbin_in[4][21][18];
assign sum_out[21][19] = accbin_in[0][21][19] + accbin_in[1][21][19] + accbin_in[2][21][19] + accbin_in[3][21][19] + accbin_in[4][21][19];
assign sum_out[21][20] = accbin_in[0][21][20] + accbin_in[1][21][20] + accbin_in[2][21][20] + accbin_in[3][21][20] + accbin_in[4][21][20];
assign sum_out[21][21] = accbin_in[0][21][21] + accbin_in[1][21][21] + accbin_in[2][21][21] + accbin_in[3][21][21] + accbin_in[4][21][21];
assign sum_out[21][22] = accbin_in[0][21][22] + accbin_in[1][21][22] + accbin_in[2][21][22] + accbin_in[3][21][22] + accbin_in[4][21][22];
assign sum_out[21][23] = accbin_in[0][21][23] + accbin_in[1][21][23] + accbin_in[2][21][23] + accbin_in[3][21][23] + accbin_in[4][21][23];
assign sum_out[22][0] = accbin_in[0][22][0] + accbin_in[1][22][0] + accbin_in[2][22][0] + accbin_in[3][22][0] + accbin_in[4][22][0];
assign sum_out[22][1] = accbin_in[0][22][1] + accbin_in[1][22][1] + accbin_in[2][22][1] + accbin_in[3][22][1] + accbin_in[4][22][1];
assign sum_out[22][2] = accbin_in[0][22][2] + accbin_in[1][22][2] + accbin_in[2][22][2] + accbin_in[3][22][2] + accbin_in[4][22][2];
assign sum_out[22][3] = accbin_in[0][22][3] + accbin_in[1][22][3] + accbin_in[2][22][3] + accbin_in[3][22][3] + accbin_in[4][22][3];
assign sum_out[22][4] = accbin_in[0][22][4] + accbin_in[1][22][4] + accbin_in[2][22][4] + accbin_in[3][22][4] + accbin_in[4][22][4];
assign sum_out[22][5] = accbin_in[0][22][5] + accbin_in[1][22][5] + accbin_in[2][22][5] + accbin_in[3][22][5] + accbin_in[4][22][5];
assign sum_out[22][6] = accbin_in[0][22][6] + accbin_in[1][22][6] + accbin_in[2][22][6] + accbin_in[3][22][6] + accbin_in[4][22][6];
assign sum_out[22][7] = accbin_in[0][22][7] + accbin_in[1][22][7] + accbin_in[2][22][7] + accbin_in[3][22][7] + accbin_in[4][22][7];
assign sum_out[22][8] = accbin_in[0][22][8] + accbin_in[1][22][8] + accbin_in[2][22][8] + accbin_in[3][22][8] + accbin_in[4][22][8];
assign sum_out[22][9] = accbin_in[0][22][9] + accbin_in[1][22][9] + accbin_in[2][22][9] + accbin_in[3][22][9] + accbin_in[4][22][9];
assign sum_out[22][10] = accbin_in[0][22][10] + accbin_in[1][22][10] + accbin_in[2][22][10] + accbin_in[3][22][10] + accbin_in[4][22][10];
assign sum_out[22][11] = accbin_in[0][22][11] + accbin_in[1][22][11] + accbin_in[2][22][11] + accbin_in[3][22][11] + accbin_in[4][22][11];
assign sum_out[22][12] = accbin_in[0][22][12] + accbin_in[1][22][12] + accbin_in[2][22][12] + accbin_in[3][22][12] + accbin_in[4][22][12];
assign sum_out[22][13] = accbin_in[0][22][13] + accbin_in[1][22][13] + accbin_in[2][22][13] + accbin_in[3][22][13] + accbin_in[4][22][13];
assign sum_out[22][14] = accbin_in[0][22][14] + accbin_in[1][22][14] + accbin_in[2][22][14] + accbin_in[3][22][14] + accbin_in[4][22][14];
assign sum_out[22][15] = accbin_in[0][22][15] + accbin_in[1][22][15] + accbin_in[2][22][15] + accbin_in[3][22][15] + accbin_in[4][22][15];
assign sum_out[22][16] = accbin_in[0][22][16] + accbin_in[1][22][16] + accbin_in[2][22][16] + accbin_in[3][22][16] + accbin_in[4][22][16];
assign sum_out[22][17] = accbin_in[0][22][17] + accbin_in[1][22][17] + accbin_in[2][22][17] + accbin_in[3][22][17] + accbin_in[4][22][17];
assign sum_out[22][18] = accbin_in[0][22][18] + accbin_in[1][22][18] + accbin_in[2][22][18] + accbin_in[3][22][18] + accbin_in[4][22][18];
assign sum_out[22][19] = accbin_in[0][22][19] + accbin_in[1][22][19] + accbin_in[2][22][19] + accbin_in[3][22][19] + accbin_in[4][22][19];
assign sum_out[22][20] = accbin_in[0][22][20] + accbin_in[1][22][20] + accbin_in[2][22][20] + accbin_in[3][22][20] + accbin_in[4][22][20];
assign sum_out[22][21] = accbin_in[0][22][21] + accbin_in[1][22][21] + accbin_in[2][22][21] + accbin_in[3][22][21] + accbin_in[4][22][21];
assign sum_out[22][22] = accbin_in[0][22][22] + accbin_in[1][22][22] + accbin_in[2][22][22] + accbin_in[3][22][22] + accbin_in[4][22][22];
assign sum_out[22][23] = accbin_in[0][22][23] + accbin_in[1][22][23] + accbin_in[2][22][23] + accbin_in[3][22][23] + accbin_in[4][22][23];
assign sum_out[23][0] = accbin_in[0][23][0] + accbin_in[1][23][0] + accbin_in[2][23][0] + accbin_in[3][23][0] + accbin_in[4][23][0];
assign sum_out[23][1] = accbin_in[0][23][1] + accbin_in[1][23][1] + accbin_in[2][23][1] + accbin_in[3][23][1] + accbin_in[4][23][1];
assign sum_out[23][2] = accbin_in[0][23][2] + accbin_in[1][23][2] + accbin_in[2][23][2] + accbin_in[3][23][2] + accbin_in[4][23][2];
assign sum_out[23][3] = accbin_in[0][23][3] + accbin_in[1][23][3] + accbin_in[2][23][3] + accbin_in[3][23][3] + accbin_in[4][23][3];
assign sum_out[23][4] = accbin_in[0][23][4] + accbin_in[1][23][4] + accbin_in[2][23][4] + accbin_in[3][23][4] + accbin_in[4][23][4];
assign sum_out[23][5] = accbin_in[0][23][5] + accbin_in[1][23][5] + accbin_in[2][23][5] + accbin_in[3][23][5] + accbin_in[4][23][5];
assign sum_out[23][6] = accbin_in[0][23][6] + accbin_in[1][23][6] + accbin_in[2][23][6] + accbin_in[3][23][6] + accbin_in[4][23][6];
assign sum_out[23][7] = accbin_in[0][23][7] + accbin_in[1][23][7] + accbin_in[2][23][7] + accbin_in[3][23][7] + accbin_in[4][23][7];
assign sum_out[23][8] = accbin_in[0][23][8] + accbin_in[1][23][8] + accbin_in[2][23][8] + accbin_in[3][23][8] + accbin_in[4][23][8];
assign sum_out[23][9] = accbin_in[0][23][9] + accbin_in[1][23][9] + accbin_in[2][23][9] + accbin_in[3][23][9] + accbin_in[4][23][9];
assign sum_out[23][10] = accbin_in[0][23][10] + accbin_in[1][23][10] + accbin_in[2][23][10] + accbin_in[3][23][10] + accbin_in[4][23][10];
assign sum_out[23][11] = accbin_in[0][23][11] + accbin_in[1][23][11] + accbin_in[2][23][11] + accbin_in[3][23][11] + accbin_in[4][23][11];
assign sum_out[23][12] = accbin_in[0][23][12] + accbin_in[1][23][12] + accbin_in[2][23][12] + accbin_in[3][23][12] + accbin_in[4][23][12];
assign sum_out[23][13] = accbin_in[0][23][13] + accbin_in[1][23][13] + accbin_in[2][23][13] + accbin_in[3][23][13] + accbin_in[4][23][13];
assign sum_out[23][14] = accbin_in[0][23][14] + accbin_in[1][23][14] + accbin_in[2][23][14] + accbin_in[3][23][14] + accbin_in[4][23][14];
assign sum_out[23][15] = accbin_in[0][23][15] + accbin_in[1][23][15] + accbin_in[2][23][15] + accbin_in[3][23][15] + accbin_in[4][23][15];
assign sum_out[23][16] = accbin_in[0][23][16] + accbin_in[1][23][16] + accbin_in[2][23][16] + accbin_in[3][23][16] + accbin_in[4][23][16];
assign sum_out[23][17] = accbin_in[0][23][17] + accbin_in[1][23][17] + accbin_in[2][23][17] + accbin_in[3][23][17] + accbin_in[4][23][17];
assign sum_out[23][18] = accbin_in[0][23][18] + accbin_in[1][23][18] + accbin_in[2][23][18] + accbin_in[3][23][18] + accbin_in[4][23][18];
assign sum_out[23][19] = accbin_in[0][23][19] + accbin_in[1][23][19] + accbin_in[2][23][19] + accbin_in[3][23][19] + accbin_in[4][23][19];
assign sum_out[23][20] = accbin_in[0][23][20] + accbin_in[1][23][20] + accbin_in[2][23][20] + accbin_in[3][23][20] + accbin_in[4][23][20];
assign sum_out[23][21] = accbin_in[0][23][21] + accbin_in[1][23][21] + accbin_in[2][23][21] + accbin_in[3][23][21] + accbin_in[4][23][21];
assign sum_out[23][22] = accbin_in[0][23][22] + accbin_in[1][23][22] + accbin_in[2][23][22] + accbin_in[3][23][22] + accbin_in[4][23][22];
assign sum_out[23][23] = accbin_in[0][23][23] + accbin_in[1][23][23] + accbin_in[2][23][23] + accbin_in[3][23][23] + accbin_in[4][23][23];

assign accbin_out[0][0] = (sum_out[0][0] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[0][1] = (sum_out[0][1] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[0][2] = (sum_out[0][2] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[0][3] = (sum_out[0][3] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[0][4] = (sum_out[0][4] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[0][5] = (sum_out[0][5] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[0][6] = (sum_out[0][6] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[0][7] = (sum_out[0][7] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[0][8] = (sum_out[0][8] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[0][9] = (sum_out[0][9] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[0][10] = (sum_out[0][10] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[0][11] = (sum_out[0][11] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[0][12] = (sum_out[0][12] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[0][13] = (sum_out[0][13] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[0][14] = (sum_out[0][14] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[0][15] = (sum_out[0][15] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[0][16] = (sum_out[0][16] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[0][17] = (sum_out[0][17] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[0][18] = (sum_out[0][18] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[0][19] = (sum_out[0][19] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[0][20] = (sum_out[0][20] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[0][21] = (sum_out[0][21] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[0][22] = (sum_out[0][22] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[0][23] = (sum_out[0][23] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[1][0] = (sum_out[1][0] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[1][1] = (sum_out[1][1] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[1][2] = (sum_out[1][2] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[1][3] = (sum_out[1][3] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[1][4] = (sum_out[1][4] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[1][5] = (sum_out[1][5] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[1][6] = (sum_out[1][6] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[1][7] = (sum_out[1][7] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[1][8] = (sum_out[1][8] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[1][9] = (sum_out[1][9] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[1][10] = (sum_out[1][10] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[1][11] = (sum_out[1][11] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[1][12] = (sum_out[1][12] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[1][13] = (sum_out[1][13] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[1][14] = (sum_out[1][14] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[1][15] = (sum_out[1][15] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[1][16] = (sum_out[1][16] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[1][17] = (sum_out[1][17] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[1][18] = (sum_out[1][18] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[1][19] = (sum_out[1][19] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[1][20] = (sum_out[1][20] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[1][21] = (sum_out[1][21] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[1][22] = (sum_out[1][22] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[1][23] = (sum_out[1][23] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[2][0] = (sum_out[2][0] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[2][1] = (sum_out[2][1] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[2][2] = (sum_out[2][2] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[2][3] = (sum_out[2][3] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[2][4] = (sum_out[2][4] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[2][5] = (sum_out[2][5] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[2][6] = (sum_out[2][6] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[2][7] = (sum_out[2][7] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[2][8] = (sum_out[2][8] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[2][9] = (sum_out[2][9] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[2][10] = (sum_out[2][10] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[2][11] = (sum_out[2][11] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[2][12] = (sum_out[2][12] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[2][13] = (sum_out[2][13] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[2][14] = (sum_out[2][14] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[2][15] = (sum_out[2][15] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[2][16] = (sum_out[2][16] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[2][17] = (sum_out[2][17] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[2][18] = (sum_out[2][18] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[2][19] = (sum_out[2][19] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[2][20] = (sum_out[2][20] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[2][21] = (sum_out[2][21] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[2][22] = (sum_out[2][22] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[2][23] = (sum_out[2][23] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[3][0] = (sum_out[3][0] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[3][1] = (sum_out[3][1] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[3][2] = (sum_out[3][2] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[3][3] = (sum_out[3][3] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[3][4] = (sum_out[3][4] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[3][5] = (sum_out[3][5] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[3][6] = (sum_out[3][6] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[3][7] = (sum_out[3][7] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[3][8] = (sum_out[3][8] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[3][9] = (sum_out[3][9] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[3][10] = (sum_out[3][10] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[3][11] = (sum_out[3][11] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[3][12] = (sum_out[3][12] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[3][13] = (sum_out[3][13] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[3][14] = (sum_out[3][14] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[3][15] = (sum_out[3][15] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[3][16] = (sum_out[3][16] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[3][17] = (sum_out[3][17] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[3][18] = (sum_out[3][18] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[3][19] = (sum_out[3][19] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[3][20] = (sum_out[3][20] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[3][21] = (sum_out[3][21] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[3][22] = (sum_out[3][22] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[3][23] = (sum_out[3][23] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[4][0] = (sum_out[4][0] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[4][1] = (sum_out[4][1] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[4][2] = (sum_out[4][2] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[4][3] = (sum_out[4][3] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[4][4] = (sum_out[4][4] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[4][5] = (sum_out[4][5] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[4][6] = (sum_out[4][6] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[4][7] = (sum_out[4][7] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[4][8] = (sum_out[4][8] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[4][9] = (sum_out[4][9] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[4][10] = (sum_out[4][10] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[4][11] = (sum_out[4][11] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[4][12] = (sum_out[4][12] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[4][13] = (sum_out[4][13] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[4][14] = (sum_out[4][14] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[4][15] = (sum_out[4][15] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[4][16] = (sum_out[4][16] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[4][17] = (sum_out[4][17] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[4][18] = (sum_out[4][18] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[4][19] = (sum_out[4][19] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[4][20] = (sum_out[4][20] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[4][21] = (sum_out[4][21] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[4][22] = (sum_out[4][22] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[4][23] = (sum_out[4][23] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[5][0] = (sum_out[5][0] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[5][1] = (sum_out[5][1] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[5][2] = (sum_out[5][2] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[5][3] = (sum_out[5][3] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[5][4] = (sum_out[5][4] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[5][5] = (sum_out[5][5] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[5][6] = (sum_out[5][6] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[5][7] = (sum_out[5][7] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[5][8] = (sum_out[5][8] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[5][9] = (sum_out[5][9] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[5][10] = (sum_out[5][10] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[5][11] = (sum_out[5][11] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[5][12] = (sum_out[5][12] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[5][13] = (sum_out[5][13] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[5][14] = (sum_out[5][14] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[5][15] = (sum_out[5][15] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[5][16] = (sum_out[5][16] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[5][17] = (sum_out[5][17] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[5][18] = (sum_out[5][18] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[5][19] = (sum_out[5][19] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[5][20] = (sum_out[5][20] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[5][21] = (sum_out[5][21] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[5][22] = (sum_out[5][22] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[5][23] = (sum_out[5][23] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[6][0] = (sum_out[6][0] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[6][1] = (sum_out[6][1] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[6][2] = (sum_out[6][2] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[6][3] = (sum_out[6][3] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[6][4] = (sum_out[6][4] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[6][5] = (sum_out[6][5] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[6][6] = (sum_out[6][6] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[6][7] = (sum_out[6][7] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[6][8] = (sum_out[6][8] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[6][9] = (sum_out[6][9] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[6][10] = (sum_out[6][10] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[6][11] = (sum_out[6][11] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[6][12] = (sum_out[6][12] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[6][13] = (sum_out[6][13] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[6][14] = (sum_out[6][14] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[6][15] = (sum_out[6][15] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[6][16] = (sum_out[6][16] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[6][17] = (sum_out[6][17] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[6][18] = (sum_out[6][18] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[6][19] = (sum_out[6][19] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[6][20] = (sum_out[6][20] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[6][21] = (sum_out[6][21] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[6][22] = (sum_out[6][22] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[6][23] = (sum_out[6][23] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[7][0] = (sum_out[7][0] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[7][1] = (sum_out[7][1] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[7][2] = (sum_out[7][2] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[7][3] = (sum_out[7][3] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[7][4] = (sum_out[7][4] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[7][5] = (sum_out[7][5] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[7][6] = (sum_out[7][6] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[7][7] = (sum_out[7][7] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[7][8] = (sum_out[7][8] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[7][9] = (sum_out[7][9] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[7][10] = (sum_out[7][10] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[7][11] = (sum_out[7][11] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[7][12] = (sum_out[7][12] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[7][13] = (sum_out[7][13] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[7][14] = (sum_out[7][14] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[7][15] = (sum_out[7][15] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[7][16] = (sum_out[7][16] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[7][17] = (sum_out[7][17] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[7][18] = (sum_out[7][18] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[7][19] = (sum_out[7][19] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[7][20] = (sum_out[7][20] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[7][21] = (sum_out[7][21] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[7][22] = (sum_out[7][22] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[7][23] = (sum_out[7][23] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[8][0] = (sum_out[8][0] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[8][1] = (sum_out[8][1] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[8][2] = (sum_out[8][2] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[8][3] = (sum_out[8][3] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[8][4] = (sum_out[8][4] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[8][5] = (sum_out[8][5] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[8][6] = (sum_out[8][6] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[8][7] = (sum_out[8][7] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[8][8] = (sum_out[8][8] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[8][9] = (sum_out[8][9] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[8][10] = (sum_out[8][10] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[8][11] = (sum_out[8][11] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[8][12] = (sum_out[8][12] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[8][13] = (sum_out[8][13] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[8][14] = (sum_out[8][14] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[8][15] = (sum_out[8][15] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[8][16] = (sum_out[8][16] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[8][17] = (sum_out[8][17] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[8][18] = (sum_out[8][18] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[8][19] = (sum_out[8][19] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[8][20] = (sum_out[8][20] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[8][21] = (sum_out[8][21] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[8][22] = (sum_out[8][22] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[8][23] = (sum_out[8][23] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[9][0] = (sum_out[9][0] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[9][1] = (sum_out[9][1] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[9][2] = (sum_out[9][2] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[9][3] = (sum_out[9][3] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[9][4] = (sum_out[9][4] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[9][5] = (sum_out[9][5] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[9][6] = (sum_out[9][6] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[9][7] = (sum_out[9][7] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[9][8] = (sum_out[9][8] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[9][9] = (sum_out[9][9] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[9][10] = (sum_out[9][10] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[9][11] = (sum_out[9][11] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[9][12] = (sum_out[9][12] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[9][13] = (sum_out[9][13] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[9][14] = (sum_out[9][14] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[9][15] = (sum_out[9][15] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[9][16] = (sum_out[9][16] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[9][17] = (sum_out[9][17] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[9][18] = (sum_out[9][18] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[9][19] = (sum_out[9][19] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[9][20] = (sum_out[9][20] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[9][21] = (sum_out[9][21] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[9][22] = (sum_out[9][22] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[9][23] = (sum_out[9][23] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[10][0] = (sum_out[10][0] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[10][1] = (sum_out[10][1] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[10][2] = (sum_out[10][2] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[10][3] = (sum_out[10][3] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[10][4] = (sum_out[10][4] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[10][5] = (sum_out[10][5] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[10][6] = (sum_out[10][6] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[10][7] = (sum_out[10][7] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[10][8] = (sum_out[10][8] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[10][9] = (sum_out[10][9] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[10][10] = (sum_out[10][10] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[10][11] = (sum_out[10][11] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[10][12] = (sum_out[10][12] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[10][13] = (sum_out[10][13] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[10][14] = (sum_out[10][14] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[10][15] = (sum_out[10][15] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[10][16] = (sum_out[10][16] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[10][17] = (sum_out[10][17] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[10][18] = (sum_out[10][18] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[10][19] = (sum_out[10][19] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[10][20] = (sum_out[10][20] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[10][21] = (sum_out[10][21] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[10][22] = (sum_out[10][22] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[10][23] = (sum_out[10][23] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[11][0] = (sum_out[11][0] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[11][1] = (sum_out[11][1] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[11][2] = (sum_out[11][2] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[11][3] = (sum_out[11][3] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[11][4] = (sum_out[11][4] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[11][5] = (sum_out[11][5] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[11][6] = (sum_out[11][6] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[11][7] = (sum_out[11][7] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[11][8] = (sum_out[11][8] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[11][9] = (sum_out[11][9] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[11][10] = (sum_out[11][10] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[11][11] = (sum_out[11][11] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[11][12] = (sum_out[11][12] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[11][13] = (sum_out[11][13] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[11][14] = (sum_out[11][14] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[11][15] = (sum_out[11][15] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[11][16] = (sum_out[11][16] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[11][17] = (sum_out[11][17] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[11][18] = (sum_out[11][18] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[11][19] = (sum_out[11][19] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[11][20] = (sum_out[11][20] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[11][21] = (sum_out[11][21] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[11][22] = (sum_out[11][22] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[11][23] = (sum_out[11][23] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[12][0] = (sum_out[12][0] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[12][1] = (sum_out[12][1] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[12][2] = (sum_out[12][2] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[12][3] = (sum_out[12][3] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[12][4] = (sum_out[12][4] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[12][5] = (sum_out[12][5] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[12][6] = (sum_out[12][6] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[12][7] = (sum_out[12][7] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[12][8] = (sum_out[12][8] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[12][9] = (sum_out[12][9] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[12][10] = (sum_out[12][10] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[12][11] = (sum_out[12][11] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[12][12] = (sum_out[12][12] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[12][13] = (sum_out[12][13] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[12][14] = (sum_out[12][14] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[12][15] = (sum_out[12][15] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[12][16] = (sum_out[12][16] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[12][17] = (sum_out[12][17] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[12][18] = (sum_out[12][18] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[12][19] = (sum_out[12][19] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[12][20] = (sum_out[12][20] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[12][21] = (sum_out[12][21] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[12][22] = (sum_out[12][22] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[12][23] = (sum_out[12][23] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[13][0] = (sum_out[13][0] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[13][1] = (sum_out[13][1] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[13][2] = (sum_out[13][2] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[13][3] = (sum_out[13][3] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[13][4] = (sum_out[13][4] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[13][5] = (sum_out[13][5] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[13][6] = (sum_out[13][6] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[13][7] = (sum_out[13][7] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[13][8] = (sum_out[13][8] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[13][9] = (sum_out[13][9] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[13][10] = (sum_out[13][10] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[13][11] = (sum_out[13][11] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[13][12] = (sum_out[13][12] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[13][13] = (sum_out[13][13] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[13][14] = (sum_out[13][14] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[13][15] = (sum_out[13][15] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[13][16] = (sum_out[13][16] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[13][17] = (sum_out[13][17] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[13][18] = (sum_out[13][18] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[13][19] = (sum_out[13][19] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[13][20] = (sum_out[13][20] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[13][21] = (sum_out[13][21] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[13][22] = (sum_out[13][22] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[13][23] = (sum_out[13][23] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[14][0] = (sum_out[14][0] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[14][1] = (sum_out[14][1] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[14][2] = (sum_out[14][2] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[14][3] = (sum_out[14][3] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[14][4] = (sum_out[14][4] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[14][5] = (sum_out[14][5] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[14][6] = (sum_out[14][6] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[14][7] = (sum_out[14][7] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[14][8] = (sum_out[14][8] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[14][9] = (sum_out[14][9] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[14][10] = (sum_out[14][10] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[14][11] = (sum_out[14][11] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[14][12] = (sum_out[14][12] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[14][13] = (sum_out[14][13] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[14][14] = (sum_out[14][14] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[14][15] = (sum_out[14][15] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[14][16] = (sum_out[14][16] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[14][17] = (sum_out[14][17] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[14][18] = (sum_out[14][18] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[14][19] = (sum_out[14][19] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[14][20] = (sum_out[14][20] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[14][21] = (sum_out[14][21] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[14][22] = (sum_out[14][22] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[14][23] = (sum_out[14][23] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[15][0] = (sum_out[15][0] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[15][1] = (sum_out[15][1] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[15][2] = (sum_out[15][2] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[15][3] = (sum_out[15][3] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[15][4] = (sum_out[15][4] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[15][5] = (sum_out[15][5] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[15][6] = (sum_out[15][6] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[15][7] = (sum_out[15][7] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[15][8] = (sum_out[15][8] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[15][9] = (sum_out[15][9] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[15][10] = (sum_out[15][10] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[15][11] = (sum_out[15][11] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[15][12] = (sum_out[15][12] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[15][13] = (sum_out[15][13] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[15][14] = (sum_out[15][14] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[15][15] = (sum_out[15][15] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[15][16] = (sum_out[15][16] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[15][17] = (sum_out[15][17] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[15][18] = (sum_out[15][18] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[15][19] = (sum_out[15][19] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[15][20] = (sum_out[15][20] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[15][21] = (sum_out[15][21] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[15][22] = (sum_out[15][22] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[15][23] = (sum_out[15][23] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[16][0] = (sum_out[16][0] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[16][1] = (sum_out[16][1] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[16][2] = (sum_out[16][2] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[16][3] = (sum_out[16][3] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[16][4] = (sum_out[16][4] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[16][5] = (sum_out[16][5] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[16][6] = (sum_out[16][6] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[16][7] = (sum_out[16][7] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[16][8] = (sum_out[16][8] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[16][9] = (sum_out[16][9] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[16][10] = (sum_out[16][10] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[16][11] = (sum_out[16][11] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[16][12] = (sum_out[16][12] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[16][13] = (sum_out[16][13] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[16][14] = (sum_out[16][14] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[16][15] = (sum_out[16][15] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[16][16] = (sum_out[16][16] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[16][17] = (sum_out[16][17] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[16][18] = (sum_out[16][18] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[16][19] = (sum_out[16][19] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[16][20] = (sum_out[16][20] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[16][21] = (sum_out[16][21] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[16][22] = (sum_out[16][22] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[16][23] = (sum_out[16][23] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[17][0] = (sum_out[17][0] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[17][1] = (sum_out[17][1] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[17][2] = (sum_out[17][2] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[17][3] = (sum_out[17][3] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[17][4] = (sum_out[17][4] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[17][5] = (sum_out[17][5] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[17][6] = (sum_out[17][6] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[17][7] = (sum_out[17][7] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[17][8] = (sum_out[17][8] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[17][9] = (sum_out[17][9] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[17][10] = (sum_out[17][10] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[17][11] = (sum_out[17][11] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[17][12] = (sum_out[17][12] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[17][13] = (sum_out[17][13] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[17][14] = (sum_out[17][14] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[17][15] = (sum_out[17][15] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[17][16] = (sum_out[17][16] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[17][17] = (sum_out[17][17] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[17][18] = (sum_out[17][18] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[17][19] = (sum_out[17][19] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[17][20] = (sum_out[17][20] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[17][21] = (sum_out[17][21] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[17][22] = (sum_out[17][22] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[17][23] = (sum_out[17][23] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[18][0] = (sum_out[18][0] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[18][1] = (sum_out[18][1] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[18][2] = (sum_out[18][2] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[18][3] = (sum_out[18][3] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[18][4] = (sum_out[18][4] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[18][5] = (sum_out[18][5] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[18][6] = (sum_out[18][6] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[18][7] = (sum_out[18][7] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[18][8] = (sum_out[18][8] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[18][9] = (sum_out[18][9] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[18][10] = (sum_out[18][10] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[18][11] = (sum_out[18][11] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[18][12] = (sum_out[18][12] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[18][13] = (sum_out[18][13] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[18][14] = (sum_out[18][14] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[18][15] = (sum_out[18][15] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[18][16] = (sum_out[18][16] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[18][17] = (sum_out[18][17] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[18][18] = (sum_out[18][18] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[18][19] = (sum_out[18][19] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[18][20] = (sum_out[18][20] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[18][21] = (sum_out[18][21] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[18][22] = (sum_out[18][22] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[18][23] = (sum_out[18][23] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[19][0] = (sum_out[19][0] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[19][1] = (sum_out[19][1] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[19][2] = (sum_out[19][2] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[19][3] = (sum_out[19][3] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[19][4] = (sum_out[19][4] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[19][5] = (sum_out[19][5] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[19][6] = (sum_out[19][6] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[19][7] = (sum_out[19][7] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[19][8] = (sum_out[19][8] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[19][9] = (sum_out[19][9] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[19][10] = (sum_out[19][10] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[19][11] = (sum_out[19][11] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[19][12] = (sum_out[19][12] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[19][13] = (sum_out[19][13] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[19][14] = (sum_out[19][14] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[19][15] = (sum_out[19][15] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[19][16] = (sum_out[19][16] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[19][17] = (sum_out[19][17] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[19][18] = (sum_out[19][18] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[19][19] = (sum_out[19][19] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[19][20] = (sum_out[19][20] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[19][21] = (sum_out[19][21] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[19][22] = (sum_out[19][22] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[19][23] = (sum_out[19][23] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[20][0] = (sum_out[20][0] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[20][1] = (sum_out[20][1] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[20][2] = (sum_out[20][2] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[20][3] = (sum_out[20][3] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[20][4] = (sum_out[20][4] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[20][5] = (sum_out[20][5] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[20][6] = (sum_out[20][6] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[20][7] = (sum_out[20][7] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[20][8] = (sum_out[20][8] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[20][9] = (sum_out[20][9] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[20][10] = (sum_out[20][10] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[20][11] = (sum_out[20][11] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[20][12] = (sum_out[20][12] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[20][13] = (sum_out[20][13] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[20][14] = (sum_out[20][14] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[20][15] = (sum_out[20][15] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[20][16] = (sum_out[20][16] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[20][17] = (sum_out[20][17] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[20][18] = (sum_out[20][18] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[20][19] = (sum_out[20][19] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[20][20] = (sum_out[20][20] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[20][21] = (sum_out[20][21] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[20][22] = (sum_out[20][22] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[20][23] = (sum_out[20][23] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[21][0] = (sum_out[21][0] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[21][1] = (sum_out[21][1] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[21][2] = (sum_out[21][2] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[21][3] = (sum_out[21][3] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[21][4] = (sum_out[21][4] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[21][5] = (sum_out[21][5] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[21][6] = (sum_out[21][6] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[21][7] = (sum_out[21][7] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[21][8] = (sum_out[21][8] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[21][9] = (sum_out[21][9] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[21][10] = (sum_out[21][10] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[21][11] = (sum_out[21][11] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[21][12] = (sum_out[21][12] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[21][13] = (sum_out[21][13] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[21][14] = (sum_out[21][14] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[21][15] = (sum_out[21][15] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[21][16] = (sum_out[21][16] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[21][17] = (sum_out[21][17] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[21][18] = (sum_out[21][18] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[21][19] = (sum_out[21][19] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[21][20] = (sum_out[21][20] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[21][21] = (sum_out[21][21] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[21][22] = (sum_out[21][22] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[21][23] = (sum_out[21][23] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[22][0] = (sum_out[22][0] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[22][1] = (sum_out[22][1] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[22][2] = (sum_out[22][2] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[22][3] = (sum_out[22][3] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[22][4] = (sum_out[22][4] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[22][5] = (sum_out[22][5] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[22][6] = (sum_out[22][6] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[22][7] = (sum_out[22][7] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[22][8] = (sum_out[22][8] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[22][9] = (sum_out[22][9] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[22][10] = (sum_out[22][10] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[22][11] = (sum_out[22][11] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[22][12] = (sum_out[22][12] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[22][13] = (sum_out[22][13] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[22][14] = (sum_out[22][14] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[22][15] = (sum_out[22][15] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[22][16] = (sum_out[22][16] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[22][17] = (sum_out[22][17] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[22][18] = (sum_out[22][18] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[22][19] = (sum_out[22][19] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[22][20] = (sum_out[22][20] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[22][21] = (sum_out[22][21] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[22][22] = (sum_out[22][22] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[22][23] = (sum_out[22][23] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[23][0] = (sum_out[23][0] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[23][1] = (sum_out[23][1] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[23][2] = (sum_out[23][2] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[23][3] = (sum_out[23][3] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[23][4] = (sum_out[23][4] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[23][5] = (sum_out[23][5] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[23][6] = (sum_out[23][6] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[23][7] = (sum_out[23][7] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[23][8] = (sum_out[23][8] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[23][9] = (sum_out[23][9] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[23][10] = (sum_out[23][10] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[23][11] = (sum_out[23][11] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[23][12] = (sum_out[23][12] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[23][13] = (sum_out[23][13] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[23][14] = (sum_out[23][14] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[23][15] = (sum_out[23][15] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[23][16] = (sum_out[23][16] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[23][17] = (sum_out[23][17] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[23][18] = (sum_out[23][18] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[23][19] = (sum_out[23][19] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[23][20] = (sum_out[23][20] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[23][21] = (sum_out[23][21] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[23][22] = (sum_out[23][22] > kernel_offset) ? 1'b1 : 1'b0;
assign accbin_out[23][23] = (sum_out[23][23] > kernel_offset) ? 1'b1 : 1'b0;

endmodule