module convchan1( 
    input  logic signed image     [0:27][0:27],
    input  logic        kernel    [0:4] [0:4],
    output logic        out_fmap  [0:23][0:23]
    );

logic signed [bW-1:0] xor_sum       [0:23][0:23];
logic signed [1   :0] signed_kernel [0: 4][0: 4];


// Make kernel signed 

always_ff @(posedge clk) begin
    if(~rst_n) begin
        for(i=0; i<5; i=i+1) begin
            for(j=0; j<5; j=j+1) begin
                signed_kernel[i][j] <= 2'b00;
            end
        end
    end else begin
        for(i=0; i<5; i=i+1) begin
            for(j=0; j<5; j=j+1) begin
                signed_kernel[i][j] <= (kernel[i][j] == 1'b1) ? 2'b01 : 2'b11;
            end
        end
    end
end

assign xor_sum[0][0] = signed_kernel[0][0] ~^ image[0][0] + signed_kernel[0][1] ~^ image[0][1] + signed_kernel[0][2] ~^ image[0][2] + signed_kernel[0][3] ~^ image[0][3] + signed_kernel[0][4] ~^ image[0][4] + signed_kernel[1][0] ~^ image[1][0] + signed_kernel[1][1] ~^ image[1][1] + signed_kernel[1][2] ~^ image[1][2] + signed_kernel[1][3] ~^ image[1][3] + signed_kernel[1][4] ~^ image[1][4] + signed_kernel[2][0] ~^ image[2][0] + signed_kernel[2][1] ~^ image[2][1] + signed_kernel[2][2] ~^ image[2][2] + signed_kernel[2][3] ~^ image[2][3] + signed_kernel[2][4] ~^ image[2][4] + signed_kernel[3][0] ~^ image[3][0] + signed_kernel[3][1] ~^ image[3][1] + signed_kernel[3][2] ~^ image[3][2] + signed_kernel[3][3] ~^ image[3][3] + signed_kernel[3][4] ~^ image[3][4] + signed_kernel[4][0] ~^ image[4][0] + signed_kernel[4][1] ~^ image[4][1] + signed_kernel[4][2] ~^ image[4][2] + signed_kernel[4][3] ~^ image[4][3] + signed_kernel[4][4] ~^ image[4][4];
assign xor_sum[0][1] = signed_kernel[0][0] ~^ image[0][1] + signed_kernel[0][1] ~^ image[0][2] + signed_kernel[0][2] ~^ image[0][3] + signed_kernel[0][3] ~^ image[0][4] + signed_kernel[0][4] ~^ image[0][5] + signed_kernel[1][0] ~^ image[1][1] + signed_kernel[1][1] ~^ image[1][2] + signed_kernel[1][2] ~^ image[1][3] + signed_kernel[1][3] ~^ image[1][4] + signed_kernel[1][4] ~^ image[1][5] + signed_kernel[2][0] ~^ image[2][1] + signed_kernel[2][1] ~^ image[2][2] + signed_kernel[2][2] ~^ image[2][3] + signed_kernel[2][3] ~^ image[2][4] + signed_kernel[2][4] ~^ image[2][5] + signed_kernel[3][0] ~^ image[3][1] + signed_kernel[3][1] ~^ image[3][2] + signed_kernel[3][2] ~^ image[3][3] + signed_kernel[3][3] ~^ image[3][4] + signed_kernel[3][4] ~^ image[3][5] + signed_kernel[4][0] ~^ image[4][1] + signed_kernel[4][1] ~^ image[4][2] + signed_kernel[4][2] ~^ image[4][3] + signed_kernel[4][3] ~^ image[4][4] + signed_kernel[4][4] ~^ image[4][5];
assign xor_sum[0][2] = signed_kernel[0][0] ~^ image[0][2] + signed_kernel[0][1] ~^ image[0][3] + signed_kernel[0][2] ~^ image[0][4] + signed_kernel[0][3] ~^ image[0][5] + signed_kernel[0][4] ~^ image[0][6] + signed_kernel[1][0] ~^ image[1][2] + signed_kernel[1][1] ~^ image[1][3] + signed_kernel[1][2] ~^ image[1][4] + signed_kernel[1][3] ~^ image[1][5] + signed_kernel[1][4] ~^ image[1][6] + signed_kernel[2][0] ~^ image[2][2] + signed_kernel[2][1] ~^ image[2][3] + signed_kernel[2][2] ~^ image[2][4] + signed_kernel[2][3] ~^ image[2][5] + signed_kernel[2][4] ~^ image[2][6] + signed_kernel[3][0] ~^ image[3][2] + signed_kernel[3][1] ~^ image[3][3] + signed_kernel[3][2] ~^ image[3][4] + signed_kernel[3][3] ~^ image[3][5] + signed_kernel[3][4] ~^ image[3][6] + signed_kernel[4][0] ~^ image[4][2] + signed_kernel[4][1] ~^ image[4][3] + signed_kernel[4][2] ~^ image[4][4] + signed_kernel[4][3] ~^ image[4][5] + signed_kernel[4][4] ~^ image[4][6];
assign xor_sum[0][3] = signed_kernel[0][0] ~^ image[0][3] + signed_kernel[0][1] ~^ image[0][4] + signed_kernel[0][2] ~^ image[0][5] + signed_kernel[0][3] ~^ image[0][6] + signed_kernel[0][4] ~^ image[0][7] + signed_kernel[1][0] ~^ image[1][3] + signed_kernel[1][1] ~^ image[1][4] + signed_kernel[1][2] ~^ image[1][5] + signed_kernel[1][3] ~^ image[1][6] + signed_kernel[1][4] ~^ image[1][7] + signed_kernel[2][0] ~^ image[2][3] + signed_kernel[2][1] ~^ image[2][4] + signed_kernel[2][2] ~^ image[2][5] + signed_kernel[2][3] ~^ image[2][6] + signed_kernel[2][4] ~^ image[2][7] + signed_kernel[3][0] ~^ image[3][3] + signed_kernel[3][1] ~^ image[3][4] + signed_kernel[3][2] ~^ image[3][5] + signed_kernel[3][3] ~^ image[3][6] + signed_kernel[3][4] ~^ image[3][7] + signed_kernel[4][0] ~^ image[4][3] + signed_kernel[4][1] ~^ image[4][4] + signed_kernel[4][2] ~^ image[4][5] + signed_kernel[4][3] ~^ image[4][6] + signed_kernel[4][4] ~^ image[4][7];
assign xor_sum[0][4] = signed_kernel[0][0] ~^ image[0][4] + signed_kernel[0][1] ~^ image[0][5] + signed_kernel[0][2] ~^ image[0][6] + signed_kernel[0][3] ~^ image[0][7] + signed_kernel[0][4] ~^ image[0][8] + signed_kernel[1][0] ~^ image[1][4] + signed_kernel[1][1] ~^ image[1][5] + signed_kernel[1][2] ~^ image[1][6] + signed_kernel[1][3] ~^ image[1][7] + signed_kernel[1][4] ~^ image[1][8] + signed_kernel[2][0] ~^ image[2][4] + signed_kernel[2][1] ~^ image[2][5] + signed_kernel[2][2] ~^ image[2][6] + signed_kernel[2][3] ~^ image[2][7] + signed_kernel[2][4] ~^ image[2][8] + signed_kernel[3][0] ~^ image[3][4] + signed_kernel[3][1] ~^ image[3][5] + signed_kernel[3][2] ~^ image[3][6] + signed_kernel[3][3] ~^ image[3][7] + signed_kernel[3][4] ~^ image[3][8] + signed_kernel[4][0] ~^ image[4][4] + signed_kernel[4][1] ~^ image[4][5] + signed_kernel[4][2] ~^ image[4][6] + signed_kernel[4][3] ~^ image[4][7] + signed_kernel[4][4] ~^ image[4][8];
assign xor_sum[0][5] = signed_kernel[0][0] ~^ image[0][5] + signed_kernel[0][1] ~^ image[0][6] + signed_kernel[0][2] ~^ image[0][7] + signed_kernel[0][3] ~^ image[0][8] + signed_kernel[0][4] ~^ image[0][9] + signed_kernel[1][0] ~^ image[1][5] + signed_kernel[1][1] ~^ image[1][6] + signed_kernel[1][2] ~^ image[1][7] + signed_kernel[1][3] ~^ image[1][8] + signed_kernel[1][4] ~^ image[1][9] + signed_kernel[2][0] ~^ image[2][5] + signed_kernel[2][1] ~^ image[2][6] + signed_kernel[2][2] ~^ image[2][7] + signed_kernel[2][3] ~^ image[2][8] + signed_kernel[2][4] ~^ image[2][9] + signed_kernel[3][0] ~^ image[3][5] + signed_kernel[3][1] ~^ image[3][6] + signed_kernel[3][2] ~^ image[3][7] + signed_kernel[3][3] ~^ image[3][8] + signed_kernel[3][4] ~^ image[3][9] + signed_kernel[4][0] ~^ image[4][5] + signed_kernel[4][1] ~^ image[4][6] + signed_kernel[4][2] ~^ image[4][7] + signed_kernel[4][3] ~^ image[4][8] + signed_kernel[4][4] ~^ image[4][9];
assign xor_sum[0][6] = signed_kernel[0][0] ~^ image[0][6] + signed_kernel[0][1] ~^ image[0][7] + signed_kernel[0][2] ~^ image[0][8] + signed_kernel[0][3] ~^ image[0][9] + signed_kernel[0][4] ~^ image[0][10] + signed_kernel[1][0] ~^ image[1][6] + signed_kernel[1][1] ~^ image[1][7] + signed_kernel[1][2] ~^ image[1][8] + signed_kernel[1][3] ~^ image[1][9] + signed_kernel[1][4] ~^ image[1][10] + signed_kernel[2][0] ~^ image[2][6] + signed_kernel[2][1] ~^ image[2][7] + signed_kernel[2][2] ~^ image[2][8] + signed_kernel[2][3] ~^ image[2][9] + signed_kernel[2][4] ~^ image[2][10] + signed_kernel[3][0] ~^ image[3][6] + signed_kernel[3][1] ~^ image[3][7] + signed_kernel[3][2] ~^ image[3][8] + signed_kernel[3][3] ~^ image[3][9] + signed_kernel[3][4] ~^ image[3][10] + signed_kernel[4][0] ~^ image[4][6] + signed_kernel[4][1] ~^ image[4][7] + signed_kernel[4][2] ~^ image[4][8] + signed_kernel[4][3] ~^ image[4][9] + signed_kernel[4][4] ~^ image[4][10];
assign xor_sum[0][7] = signed_kernel[0][0] ~^ image[0][7] + signed_kernel[0][1] ~^ image[0][8] + signed_kernel[0][2] ~^ image[0][9] + signed_kernel[0][3] ~^ image[0][10] + signed_kernel[0][4] ~^ image[0][11] + signed_kernel[1][0] ~^ image[1][7] + signed_kernel[1][1] ~^ image[1][8] + signed_kernel[1][2] ~^ image[1][9] + signed_kernel[1][3] ~^ image[1][10] + signed_kernel[1][4] ~^ image[1][11] + signed_kernel[2][0] ~^ image[2][7] + signed_kernel[2][1] ~^ image[2][8] + signed_kernel[2][2] ~^ image[2][9] + signed_kernel[2][3] ~^ image[2][10] + signed_kernel[2][4] ~^ image[2][11] + signed_kernel[3][0] ~^ image[3][7] + signed_kernel[3][1] ~^ image[3][8] + signed_kernel[3][2] ~^ image[3][9] + signed_kernel[3][3] ~^ image[3][10] + signed_kernel[3][4] ~^ image[3][11] + signed_kernel[4][0] ~^ image[4][7] + signed_kernel[4][1] ~^ image[4][8] + signed_kernel[4][2] ~^ image[4][9] + signed_kernel[4][3] ~^ image[4][10] + signed_kernel[4][4] ~^ image[4][11];
assign xor_sum[0][8] = signed_kernel[0][0] ~^ image[0][8] + signed_kernel[0][1] ~^ image[0][9] + signed_kernel[0][2] ~^ image[0][10] + signed_kernel[0][3] ~^ image[0][11] + signed_kernel[0][4] ~^ image[0][12] + signed_kernel[1][0] ~^ image[1][8] + signed_kernel[1][1] ~^ image[1][9] + signed_kernel[1][2] ~^ image[1][10] + signed_kernel[1][3] ~^ image[1][11] + signed_kernel[1][4] ~^ image[1][12] + signed_kernel[2][0] ~^ image[2][8] + signed_kernel[2][1] ~^ image[2][9] + signed_kernel[2][2] ~^ image[2][10] + signed_kernel[2][3] ~^ image[2][11] + signed_kernel[2][4] ~^ image[2][12] + signed_kernel[3][0] ~^ image[3][8] + signed_kernel[3][1] ~^ image[3][9] + signed_kernel[3][2] ~^ image[3][10] + signed_kernel[3][3] ~^ image[3][11] + signed_kernel[3][4] ~^ image[3][12] + signed_kernel[4][0] ~^ image[4][8] + signed_kernel[4][1] ~^ image[4][9] + signed_kernel[4][2] ~^ image[4][10] + signed_kernel[4][3] ~^ image[4][11] + signed_kernel[4][4] ~^ image[4][12];
assign xor_sum[0][9] = signed_kernel[0][0] ~^ image[0][9] + signed_kernel[0][1] ~^ image[0][10] + signed_kernel[0][2] ~^ image[0][11] + signed_kernel[0][3] ~^ image[0][12] + signed_kernel[0][4] ~^ image[0][13] + signed_kernel[1][0] ~^ image[1][9] + signed_kernel[1][1] ~^ image[1][10] + signed_kernel[1][2] ~^ image[1][11] + signed_kernel[1][3] ~^ image[1][12] + signed_kernel[1][4] ~^ image[1][13] + signed_kernel[2][0] ~^ image[2][9] + signed_kernel[2][1] ~^ image[2][10] + signed_kernel[2][2] ~^ image[2][11] + signed_kernel[2][3] ~^ image[2][12] + signed_kernel[2][4] ~^ image[2][13] + signed_kernel[3][0] ~^ image[3][9] + signed_kernel[3][1] ~^ image[3][10] + signed_kernel[3][2] ~^ image[3][11] + signed_kernel[3][3] ~^ image[3][12] + signed_kernel[3][4] ~^ image[3][13] + signed_kernel[4][0] ~^ image[4][9] + signed_kernel[4][1] ~^ image[4][10] + signed_kernel[4][2] ~^ image[4][11] + signed_kernel[4][3] ~^ image[4][12] + signed_kernel[4][4] ~^ image[4][13];
assign xor_sum[0][10] = signed_kernel[0][0] ~^ image[0][10] + signed_kernel[0][1] ~^ image[0][11] + signed_kernel[0][2] ~^ image[0][12] + signed_kernel[0][3] ~^ image[0][13] + signed_kernel[0][4] ~^ image[0][14] + signed_kernel[1][0] ~^ image[1][10] + signed_kernel[1][1] ~^ image[1][11] + signed_kernel[1][2] ~^ image[1][12] + signed_kernel[1][3] ~^ image[1][13] + signed_kernel[1][4] ~^ image[1][14] + signed_kernel[2][0] ~^ image[2][10] + signed_kernel[2][1] ~^ image[2][11] + signed_kernel[2][2] ~^ image[2][12] + signed_kernel[2][3] ~^ image[2][13] + signed_kernel[2][4] ~^ image[2][14] + signed_kernel[3][0] ~^ image[3][10] + signed_kernel[3][1] ~^ image[3][11] + signed_kernel[3][2] ~^ image[3][12] + signed_kernel[3][3] ~^ image[3][13] + signed_kernel[3][4] ~^ image[3][14] + signed_kernel[4][0] ~^ image[4][10] + signed_kernel[4][1] ~^ image[4][11] + signed_kernel[4][2] ~^ image[4][12] + signed_kernel[4][3] ~^ image[4][13] + signed_kernel[4][4] ~^ image[4][14];
assign xor_sum[0][11] = signed_kernel[0][0] ~^ image[0][11] + signed_kernel[0][1] ~^ image[0][12] + signed_kernel[0][2] ~^ image[0][13] + signed_kernel[0][3] ~^ image[0][14] + signed_kernel[0][4] ~^ image[0][15] + signed_kernel[1][0] ~^ image[1][11] + signed_kernel[1][1] ~^ image[1][12] + signed_kernel[1][2] ~^ image[1][13] + signed_kernel[1][3] ~^ image[1][14] + signed_kernel[1][4] ~^ image[1][15] + signed_kernel[2][0] ~^ image[2][11] + signed_kernel[2][1] ~^ image[2][12] + signed_kernel[2][2] ~^ image[2][13] + signed_kernel[2][3] ~^ image[2][14] + signed_kernel[2][4] ~^ image[2][15] + signed_kernel[3][0] ~^ image[3][11] + signed_kernel[3][1] ~^ image[3][12] + signed_kernel[3][2] ~^ image[3][13] + signed_kernel[3][3] ~^ image[3][14] + signed_kernel[3][4] ~^ image[3][15] + signed_kernel[4][0] ~^ image[4][11] + signed_kernel[4][1] ~^ image[4][12] + signed_kernel[4][2] ~^ image[4][13] + signed_kernel[4][3] ~^ image[4][14] + signed_kernel[4][4] ~^ image[4][15];
assign xor_sum[0][12] = signed_kernel[0][0] ~^ image[0][12] + signed_kernel[0][1] ~^ image[0][13] + signed_kernel[0][2] ~^ image[0][14] + signed_kernel[0][3] ~^ image[0][15] + signed_kernel[0][4] ~^ image[0][16] + signed_kernel[1][0] ~^ image[1][12] + signed_kernel[1][1] ~^ image[1][13] + signed_kernel[1][2] ~^ image[1][14] + signed_kernel[1][3] ~^ image[1][15] + signed_kernel[1][4] ~^ image[1][16] + signed_kernel[2][0] ~^ image[2][12] + signed_kernel[2][1] ~^ image[2][13] + signed_kernel[2][2] ~^ image[2][14] + signed_kernel[2][3] ~^ image[2][15] + signed_kernel[2][4] ~^ image[2][16] + signed_kernel[3][0] ~^ image[3][12] + signed_kernel[3][1] ~^ image[3][13] + signed_kernel[3][2] ~^ image[3][14] + signed_kernel[3][3] ~^ image[3][15] + signed_kernel[3][4] ~^ image[3][16] + signed_kernel[4][0] ~^ image[4][12] + signed_kernel[4][1] ~^ image[4][13] + signed_kernel[4][2] ~^ image[4][14] + signed_kernel[4][3] ~^ image[4][15] + signed_kernel[4][4] ~^ image[4][16];
assign xor_sum[0][13] = signed_kernel[0][0] ~^ image[0][13] + signed_kernel[0][1] ~^ image[0][14] + signed_kernel[0][2] ~^ image[0][15] + signed_kernel[0][3] ~^ image[0][16] + signed_kernel[0][4] ~^ image[0][17] + signed_kernel[1][0] ~^ image[1][13] + signed_kernel[1][1] ~^ image[1][14] + signed_kernel[1][2] ~^ image[1][15] + signed_kernel[1][3] ~^ image[1][16] + signed_kernel[1][4] ~^ image[1][17] + signed_kernel[2][0] ~^ image[2][13] + signed_kernel[2][1] ~^ image[2][14] + signed_kernel[2][2] ~^ image[2][15] + signed_kernel[2][3] ~^ image[2][16] + signed_kernel[2][4] ~^ image[2][17] + signed_kernel[3][0] ~^ image[3][13] + signed_kernel[3][1] ~^ image[3][14] + signed_kernel[3][2] ~^ image[3][15] + signed_kernel[3][3] ~^ image[3][16] + signed_kernel[3][4] ~^ image[3][17] + signed_kernel[4][0] ~^ image[4][13] + signed_kernel[4][1] ~^ image[4][14] + signed_kernel[4][2] ~^ image[4][15] + signed_kernel[4][3] ~^ image[4][16] + signed_kernel[4][4] ~^ image[4][17];
assign xor_sum[0][14] = signed_kernel[0][0] ~^ image[0][14] + signed_kernel[0][1] ~^ image[0][15] + signed_kernel[0][2] ~^ image[0][16] + signed_kernel[0][3] ~^ image[0][17] + signed_kernel[0][4] ~^ image[0][18] + signed_kernel[1][0] ~^ image[1][14] + signed_kernel[1][1] ~^ image[1][15] + signed_kernel[1][2] ~^ image[1][16] + signed_kernel[1][3] ~^ image[1][17] + signed_kernel[1][4] ~^ image[1][18] + signed_kernel[2][0] ~^ image[2][14] + signed_kernel[2][1] ~^ image[2][15] + signed_kernel[2][2] ~^ image[2][16] + signed_kernel[2][3] ~^ image[2][17] + signed_kernel[2][4] ~^ image[2][18] + signed_kernel[3][0] ~^ image[3][14] + signed_kernel[3][1] ~^ image[3][15] + signed_kernel[3][2] ~^ image[3][16] + signed_kernel[3][3] ~^ image[3][17] + signed_kernel[3][4] ~^ image[3][18] + signed_kernel[4][0] ~^ image[4][14] + signed_kernel[4][1] ~^ image[4][15] + signed_kernel[4][2] ~^ image[4][16] + signed_kernel[4][3] ~^ image[4][17] + signed_kernel[4][4] ~^ image[4][18];
assign xor_sum[0][15] = signed_kernel[0][0] ~^ image[0][15] + signed_kernel[0][1] ~^ image[0][16] + signed_kernel[0][2] ~^ image[0][17] + signed_kernel[0][3] ~^ image[0][18] + signed_kernel[0][4] ~^ image[0][19] + signed_kernel[1][0] ~^ image[1][15] + signed_kernel[1][1] ~^ image[1][16] + signed_kernel[1][2] ~^ image[1][17] + signed_kernel[1][3] ~^ image[1][18] + signed_kernel[1][4] ~^ image[1][19] + signed_kernel[2][0] ~^ image[2][15] + signed_kernel[2][1] ~^ image[2][16] + signed_kernel[2][2] ~^ image[2][17] + signed_kernel[2][3] ~^ image[2][18] + signed_kernel[2][4] ~^ image[2][19] + signed_kernel[3][0] ~^ image[3][15] + signed_kernel[3][1] ~^ image[3][16] + signed_kernel[3][2] ~^ image[3][17] + signed_kernel[3][3] ~^ image[3][18] + signed_kernel[3][4] ~^ image[3][19] + signed_kernel[4][0] ~^ image[4][15] + signed_kernel[4][1] ~^ image[4][16] + signed_kernel[4][2] ~^ image[4][17] + signed_kernel[4][3] ~^ image[4][18] + signed_kernel[4][4] ~^ image[4][19];
assign xor_sum[0][16] = signed_kernel[0][0] ~^ image[0][16] + signed_kernel[0][1] ~^ image[0][17] + signed_kernel[0][2] ~^ image[0][18] + signed_kernel[0][3] ~^ image[0][19] + signed_kernel[0][4] ~^ image[0][20] + signed_kernel[1][0] ~^ image[1][16] + signed_kernel[1][1] ~^ image[1][17] + signed_kernel[1][2] ~^ image[1][18] + signed_kernel[1][3] ~^ image[1][19] + signed_kernel[1][4] ~^ image[1][20] + signed_kernel[2][0] ~^ image[2][16] + signed_kernel[2][1] ~^ image[2][17] + signed_kernel[2][2] ~^ image[2][18] + signed_kernel[2][3] ~^ image[2][19] + signed_kernel[2][4] ~^ image[2][20] + signed_kernel[3][0] ~^ image[3][16] + signed_kernel[3][1] ~^ image[3][17] + signed_kernel[3][2] ~^ image[3][18] + signed_kernel[3][3] ~^ image[3][19] + signed_kernel[3][4] ~^ image[3][20] + signed_kernel[4][0] ~^ image[4][16] + signed_kernel[4][1] ~^ image[4][17] + signed_kernel[4][2] ~^ image[4][18] + signed_kernel[4][3] ~^ image[4][19] + signed_kernel[4][4] ~^ image[4][20];
assign xor_sum[0][17] = signed_kernel[0][0] ~^ image[0][17] + signed_kernel[0][1] ~^ image[0][18] + signed_kernel[0][2] ~^ image[0][19] + signed_kernel[0][3] ~^ image[0][20] + signed_kernel[0][4] ~^ image[0][21] + signed_kernel[1][0] ~^ image[1][17] + signed_kernel[1][1] ~^ image[1][18] + signed_kernel[1][2] ~^ image[1][19] + signed_kernel[1][3] ~^ image[1][20] + signed_kernel[1][4] ~^ image[1][21] + signed_kernel[2][0] ~^ image[2][17] + signed_kernel[2][1] ~^ image[2][18] + signed_kernel[2][2] ~^ image[2][19] + signed_kernel[2][3] ~^ image[2][20] + signed_kernel[2][4] ~^ image[2][21] + signed_kernel[3][0] ~^ image[3][17] + signed_kernel[3][1] ~^ image[3][18] + signed_kernel[3][2] ~^ image[3][19] + signed_kernel[3][3] ~^ image[3][20] + signed_kernel[3][4] ~^ image[3][21] + signed_kernel[4][0] ~^ image[4][17] + signed_kernel[4][1] ~^ image[4][18] + signed_kernel[4][2] ~^ image[4][19] + signed_kernel[4][3] ~^ image[4][20] + signed_kernel[4][4] ~^ image[4][21];
assign xor_sum[0][18] = signed_kernel[0][0] ~^ image[0][18] + signed_kernel[0][1] ~^ image[0][19] + signed_kernel[0][2] ~^ image[0][20] + signed_kernel[0][3] ~^ image[0][21] + signed_kernel[0][4] ~^ image[0][22] + signed_kernel[1][0] ~^ image[1][18] + signed_kernel[1][1] ~^ image[1][19] + signed_kernel[1][2] ~^ image[1][20] + signed_kernel[1][3] ~^ image[1][21] + signed_kernel[1][4] ~^ image[1][22] + signed_kernel[2][0] ~^ image[2][18] + signed_kernel[2][1] ~^ image[2][19] + signed_kernel[2][2] ~^ image[2][20] + signed_kernel[2][3] ~^ image[2][21] + signed_kernel[2][4] ~^ image[2][22] + signed_kernel[3][0] ~^ image[3][18] + signed_kernel[3][1] ~^ image[3][19] + signed_kernel[3][2] ~^ image[3][20] + signed_kernel[3][3] ~^ image[3][21] + signed_kernel[3][4] ~^ image[3][22] + signed_kernel[4][0] ~^ image[4][18] + signed_kernel[4][1] ~^ image[4][19] + signed_kernel[4][2] ~^ image[4][20] + signed_kernel[4][3] ~^ image[4][21] + signed_kernel[4][4] ~^ image[4][22];
assign xor_sum[0][19] = signed_kernel[0][0] ~^ image[0][19] + signed_kernel[0][1] ~^ image[0][20] + signed_kernel[0][2] ~^ image[0][21] + signed_kernel[0][3] ~^ image[0][22] + signed_kernel[0][4] ~^ image[0][23] + signed_kernel[1][0] ~^ image[1][19] + signed_kernel[1][1] ~^ image[1][20] + signed_kernel[1][2] ~^ image[1][21] + signed_kernel[1][3] ~^ image[1][22] + signed_kernel[1][4] ~^ image[1][23] + signed_kernel[2][0] ~^ image[2][19] + signed_kernel[2][1] ~^ image[2][20] + signed_kernel[2][2] ~^ image[2][21] + signed_kernel[2][3] ~^ image[2][22] + signed_kernel[2][4] ~^ image[2][23] + signed_kernel[3][0] ~^ image[3][19] + signed_kernel[3][1] ~^ image[3][20] + signed_kernel[3][2] ~^ image[3][21] + signed_kernel[3][3] ~^ image[3][22] + signed_kernel[3][4] ~^ image[3][23] + signed_kernel[4][0] ~^ image[4][19] + signed_kernel[4][1] ~^ image[4][20] + signed_kernel[4][2] ~^ image[4][21] + signed_kernel[4][3] ~^ image[4][22] + signed_kernel[4][4] ~^ image[4][23];
assign xor_sum[0][20] = signed_kernel[0][0] ~^ image[0][20] + signed_kernel[0][1] ~^ image[0][21] + signed_kernel[0][2] ~^ image[0][22] + signed_kernel[0][3] ~^ image[0][23] + signed_kernel[0][4] ~^ image[0][24] + signed_kernel[1][0] ~^ image[1][20] + signed_kernel[1][1] ~^ image[1][21] + signed_kernel[1][2] ~^ image[1][22] + signed_kernel[1][3] ~^ image[1][23] + signed_kernel[1][4] ~^ image[1][24] + signed_kernel[2][0] ~^ image[2][20] + signed_kernel[2][1] ~^ image[2][21] + signed_kernel[2][2] ~^ image[2][22] + signed_kernel[2][3] ~^ image[2][23] + signed_kernel[2][4] ~^ image[2][24] + signed_kernel[3][0] ~^ image[3][20] + signed_kernel[3][1] ~^ image[3][21] + signed_kernel[3][2] ~^ image[3][22] + signed_kernel[3][3] ~^ image[3][23] + signed_kernel[3][4] ~^ image[3][24] + signed_kernel[4][0] ~^ image[4][20] + signed_kernel[4][1] ~^ image[4][21] + signed_kernel[4][2] ~^ image[4][22] + signed_kernel[4][3] ~^ image[4][23] + signed_kernel[4][4] ~^ image[4][24];
assign xor_sum[0][21] = signed_kernel[0][0] ~^ image[0][21] + signed_kernel[0][1] ~^ image[0][22] + signed_kernel[0][2] ~^ image[0][23] + signed_kernel[0][3] ~^ image[0][24] + signed_kernel[0][4] ~^ image[0][25] + signed_kernel[1][0] ~^ image[1][21] + signed_kernel[1][1] ~^ image[1][22] + signed_kernel[1][2] ~^ image[1][23] + signed_kernel[1][3] ~^ image[1][24] + signed_kernel[1][4] ~^ image[1][25] + signed_kernel[2][0] ~^ image[2][21] + signed_kernel[2][1] ~^ image[2][22] + signed_kernel[2][2] ~^ image[2][23] + signed_kernel[2][3] ~^ image[2][24] + signed_kernel[2][4] ~^ image[2][25] + signed_kernel[3][0] ~^ image[3][21] + signed_kernel[3][1] ~^ image[3][22] + signed_kernel[3][2] ~^ image[3][23] + signed_kernel[3][3] ~^ image[3][24] + signed_kernel[3][4] ~^ image[3][25] + signed_kernel[4][0] ~^ image[4][21] + signed_kernel[4][1] ~^ image[4][22] + signed_kernel[4][2] ~^ image[4][23] + signed_kernel[4][3] ~^ image[4][24] + signed_kernel[4][4] ~^ image[4][25];
assign xor_sum[0][22] = signed_kernel[0][0] ~^ image[0][22] + signed_kernel[0][1] ~^ image[0][23] + signed_kernel[0][2] ~^ image[0][24] + signed_kernel[0][3] ~^ image[0][25] + signed_kernel[0][4] ~^ image[0][26] + signed_kernel[1][0] ~^ image[1][22] + signed_kernel[1][1] ~^ image[1][23] + signed_kernel[1][2] ~^ image[1][24] + signed_kernel[1][3] ~^ image[1][25] + signed_kernel[1][4] ~^ image[1][26] + signed_kernel[2][0] ~^ image[2][22] + signed_kernel[2][1] ~^ image[2][23] + signed_kernel[2][2] ~^ image[2][24] + signed_kernel[2][3] ~^ image[2][25] + signed_kernel[2][4] ~^ image[2][26] + signed_kernel[3][0] ~^ image[3][22] + signed_kernel[3][1] ~^ image[3][23] + signed_kernel[3][2] ~^ image[3][24] + signed_kernel[3][3] ~^ image[3][25] + signed_kernel[3][4] ~^ image[3][26] + signed_kernel[4][0] ~^ image[4][22] + signed_kernel[4][1] ~^ image[4][23] + signed_kernel[4][2] ~^ image[4][24] + signed_kernel[4][3] ~^ image[4][25] + signed_kernel[4][4] ~^ image[4][26];
assign xor_sum[0][23] = signed_kernel[0][0] ~^ image[0][23] + signed_kernel[0][1] ~^ image[0][24] + signed_kernel[0][2] ~^ image[0][25] + signed_kernel[0][3] ~^ image[0][26] + signed_kernel[0][4] ~^ image[0][27] + signed_kernel[1][0] ~^ image[1][23] + signed_kernel[1][1] ~^ image[1][24] + signed_kernel[1][2] ~^ image[1][25] + signed_kernel[1][3] ~^ image[1][26] + signed_kernel[1][4] ~^ image[1][27] + signed_kernel[2][0] ~^ image[2][23] + signed_kernel[2][1] ~^ image[2][24] + signed_kernel[2][2] ~^ image[2][25] + signed_kernel[2][3] ~^ image[2][26] + signed_kernel[2][4] ~^ image[2][27] + signed_kernel[3][0] ~^ image[3][23] + signed_kernel[3][1] ~^ image[3][24] + signed_kernel[3][2] ~^ image[3][25] + signed_kernel[3][3] ~^ image[3][26] + signed_kernel[3][4] ~^ image[3][27] + signed_kernel[4][0] ~^ image[4][23] + signed_kernel[4][1] ~^ image[4][24] + signed_kernel[4][2] ~^ image[4][25] + signed_kernel[4][3] ~^ image[4][26] + signed_kernel[4][4] ~^ image[4][27];
assign xor_sum[1][0] = signed_kernel[0][0] ~^ image[1][0] + signed_kernel[0][1] ~^ image[1][1] + signed_kernel[0][2] ~^ image[1][2] + signed_kernel[0][3] ~^ image[1][3] + signed_kernel[0][4] ~^ image[1][4] + signed_kernel[1][0] ~^ image[2][0] + signed_kernel[1][1] ~^ image[2][1] + signed_kernel[1][2] ~^ image[2][2] + signed_kernel[1][3] ~^ image[2][3] + signed_kernel[1][4] ~^ image[2][4] + signed_kernel[2][0] ~^ image[3][0] + signed_kernel[2][1] ~^ image[3][1] + signed_kernel[2][2] ~^ image[3][2] + signed_kernel[2][3] ~^ image[3][3] + signed_kernel[2][4] ~^ image[3][4] + signed_kernel[3][0] ~^ image[4][0] + signed_kernel[3][1] ~^ image[4][1] + signed_kernel[3][2] ~^ image[4][2] + signed_kernel[3][3] ~^ image[4][3] + signed_kernel[3][4] ~^ image[4][4] + signed_kernel[4][0] ~^ image[5][0] + signed_kernel[4][1] ~^ image[5][1] + signed_kernel[4][2] ~^ image[5][2] + signed_kernel[4][3] ~^ image[5][3] + signed_kernel[4][4] ~^ image[5][4];
assign xor_sum[1][1] = signed_kernel[0][0] ~^ image[1][1] + signed_kernel[0][1] ~^ image[1][2] + signed_kernel[0][2] ~^ image[1][3] + signed_kernel[0][3] ~^ image[1][4] + signed_kernel[0][4] ~^ image[1][5] + signed_kernel[1][0] ~^ image[2][1] + signed_kernel[1][1] ~^ image[2][2] + signed_kernel[1][2] ~^ image[2][3] + signed_kernel[1][3] ~^ image[2][4] + signed_kernel[1][4] ~^ image[2][5] + signed_kernel[2][0] ~^ image[3][1] + signed_kernel[2][1] ~^ image[3][2] + signed_kernel[2][2] ~^ image[3][3] + signed_kernel[2][3] ~^ image[3][4] + signed_kernel[2][4] ~^ image[3][5] + signed_kernel[3][0] ~^ image[4][1] + signed_kernel[3][1] ~^ image[4][2] + signed_kernel[3][2] ~^ image[4][3] + signed_kernel[3][3] ~^ image[4][4] + signed_kernel[3][4] ~^ image[4][5] + signed_kernel[4][0] ~^ image[5][1] + signed_kernel[4][1] ~^ image[5][2] + signed_kernel[4][2] ~^ image[5][3] + signed_kernel[4][3] ~^ image[5][4] + signed_kernel[4][4] ~^ image[5][5];
assign xor_sum[1][2] = signed_kernel[0][0] ~^ image[1][2] + signed_kernel[0][1] ~^ image[1][3] + signed_kernel[0][2] ~^ image[1][4] + signed_kernel[0][3] ~^ image[1][5] + signed_kernel[0][4] ~^ image[1][6] + signed_kernel[1][0] ~^ image[2][2] + signed_kernel[1][1] ~^ image[2][3] + signed_kernel[1][2] ~^ image[2][4] + signed_kernel[1][3] ~^ image[2][5] + signed_kernel[1][4] ~^ image[2][6] + signed_kernel[2][0] ~^ image[3][2] + signed_kernel[2][1] ~^ image[3][3] + signed_kernel[2][2] ~^ image[3][4] + signed_kernel[2][3] ~^ image[3][5] + signed_kernel[2][4] ~^ image[3][6] + signed_kernel[3][0] ~^ image[4][2] + signed_kernel[3][1] ~^ image[4][3] + signed_kernel[3][2] ~^ image[4][4] + signed_kernel[3][3] ~^ image[4][5] + signed_kernel[3][4] ~^ image[4][6] + signed_kernel[4][0] ~^ image[5][2] + signed_kernel[4][1] ~^ image[5][3] + signed_kernel[4][2] ~^ image[5][4] + signed_kernel[4][3] ~^ image[5][5] + signed_kernel[4][4] ~^ image[5][6];
assign xor_sum[1][3] = signed_kernel[0][0] ~^ image[1][3] + signed_kernel[0][1] ~^ image[1][4] + signed_kernel[0][2] ~^ image[1][5] + signed_kernel[0][3] ~^ image[1][6] + signed_kernel[0][4] ~^ image[1][7] + signed_kernel[1][0] ~^ image[2][3] + signed_kernel[1][1] ~^ image[2][4] + signed_kernel[1][2] ~^ image[2][5] + signed_kernel[1][3] ~^ image[2][6] + signed_kernel[1][4] ~^ image[2][7] + signed_kernel[2][0] ~^ image[3][3] + signed_kernel[2][1] ~^ image[3][4] + signed_kernel[2][2] ~^ image[3][5] + signed_kernel[2][3] ~^ image[3][6] + signed_kernel[2][4] ~^ image[3][7] + signed_kernel[3][0] ~^ image[4][3] + signed_kernel[3][1] ~^ image[4][4] + signed_kernel[3][2] ~^ image[4][5] + signed_kernel[3][3] ~^ image[4][6] + signed_kernel[3][4] ~^ image[4][7] + signed_kernel[4][0] ~^ image[5][3] + signed_kernel[4][1] ~^ image[5][4] + signed_kernel[4][2] ~^ image[5][5] + signed_kernel[4][3] ~^ image[5][6] + signed_kernel[4][4] ~^ image[5][7];
assign xor_sum[1][4] = signed_kernel[0][0] ~^ image[1][4] + signed_kernel[0][1] ~^ image[1][5] + signed_kernel[0][2] ~^ image[1][6] + signed_kernel[0][3] ~^ image[1][7] + signed_kernel[0][4] ~^ image[1][8] + signed_kernel[1][0] ~^ image[2][4] + signed_kernel[1][1] ~^ image[2][5] + signed_kernel[1][2] ~^ image[2][6] + signed_kernel[1][3] ~^ image[2][7] + signed_kernel[1][4] ~^ image[2][8] + signed_kernel[2][0] ~^ image[3][4] + signed_kernel[2][1] ~^ image[3][5] + signed_kernel[2][2] ~^ image[3][6] + signed_kernel[2][3] ~^ image[3][7] + signed_kernel[2][4] ~^ image[3][8] + signed_kernel[3][0] ~^ image[4][4] + signed_kernel[3][1] ~^ image[4][5] + signed_kernel[3][2] ~^ image[4][6] + signed_kernel[3][3] ~^ image[4][7] + signed_kernel[3][4] ~^ image[4][8] + signed_kernel[4][0] ~^ image[5][4] + signed_kernel[4][1] ~^ image[5][5] + signed_kernel[4][2] ~^ image[5][6] + signed_kernel[4][3] ~^ image[5][7] + signed_kernel[4][4] ~^ image[5][8];
assign xor_sum[1][5] = signed_kernel[0][0] ~^ image[1][5] + signed_kernel[0][1] ~^ image[1][6] + signed_kernel[0][2] ~^ image[1][7] + signed_kernel[0][3] ~^ image[1][8] + signed_kernel[0][4] ~^ image[1][9] + signed_kernel[1][0] ~^ image[2][5] + signed_kernel[1][1] ~^ image[2][6] + signed_kernel[1][2] ~^ image[2][7] + signed_kernel[1][3] ~^ image[2][8] + signed_kernel[1][4] ~^ image[2][9] + signed_kernel[2][0] ~^ image[3][5] + signed_kernel[2][1] ~^ image[3][6] + signed_kernel[2][2] ~^ image[3][7] + signed_kernel[2][3] ~^ image[3][8] + signed_kernel[2][4] ~^ image[3][9] + signed_kernel[3][0] ~^ image[4][5] + signed_kernel[3][1] ~^ image[4][6] + signed_kernel[3][2] ~^ image[4][7] + signed_kernel[3][3] ~^ image[4][8] + signed_kernel[3][4] ~^ image[4][9] + signed_kernel[4][0] ~^ image[5][5] + signed_kernel[4][1] ~^ image[5][6] + signed_kernel[4][2] ~^ image[5][7] + signed_kernel[4][3] ~^ image[5][8] + signed_kernel[4][4] ~^ image[5][9];
assign xor_sum[1][6] = signed_kernel[0][0] ~^ image[1][6] + signed_kernel[0][1] ~^ image[1][7] + signed_kernel[0][2] ~^ image[1][8] + signed_kernel[0][3] ~^ image[1][9] + signed_kernel[0][4] ~^ image[1][10] + signed_kernel[1][0] ~^ image[2][6] + signed_kernel[1][1] ~^ image[2][7] + signed_kernel[1][2] ~^ image[2][8] + signed_kernel[1][3] ~^ image[2][9] + signed_kernel[1][4] ~^ image[2][10] + signed_kernel[2][0] ~^ image[3][6] + signed_kernel[2][1] ~^ image[3][7] + signed_kernel[2][2] ~^ image[3][8] + signed_kernel[2][3] ~^ image[3][9] + signed_kernel[2][4] ~^ image[3][10] + signed_kernel[3][0] ~^ image[4][6] + signed_kernel[3][1] ~^ image[4][7] + signed_kernel[3][2] ~^ image[4][8] + signed_kernel[3][3] ~^ image[4][9] + signed_kernel[3][4] ~^ image[4][10] + signed_kernel[4][0] ~^ image[5][6] + signed_kernel[4][1] ~^ image[5][7] + signed_kernel[4][2] ~^ image[5][8] + signed_kernel[4][3] ~^ image[5][9] + signed_kernel[4][4] ~^ image[5][10];
assign xor_sum[1][7] = signed_kernel[0][0] ~^ image[1][7] + signed_kernel[0][1] ~^ image[1][8] + signed_kernel[0][2] ~^ image[1][9] + signed_kernel[0][3] ~^ image[1][10] + signed_kernel[0][4] ~^ image[1][11] + signed_kernel[1][0] ~^ image[2][7] + signed_kernel[1][1] ~^ image[2][8] + signed_kernel[1][2] ~^ image[2][9] + signed_kernel[1][3] ~^ image[2][10] + signed_kernel[1][4] ~^ image[2][11] + signed_kernel[2][0] ~^ image[3][7] + signed_kernel[2][1] ~^ image[3][8] + signed_kernel[2][2] ~^ image[3][9] + signed_kernel[2][3] ~^ image[3][10] + signed_kernel[2][4] ~^ image[3][11] + signed_kernel[3][0] ~^ image[4][7] + signed_kernel[3][1] ~^ image[4][8] + signed_kernel[3][2] ~^ image[4][9] + signed_kernel[3][3] ~^ image[4][10] + signed_kernel[3][4] ~^ image[4][11] + signed_kernel[4][0] ~^ image[5][7] + signed_kernel[4][1] ~^ image[5][8] + signed_kernel[4][2] ~^ image[5][9] + signed_kernel[4][3] ~^ image[5][10] + signed_kernel[4][4] ~^ image[5][11];
assign xor_sum[1][8] = signed_kernel[0][0] ~^ image[1][8] + signed_kernel[0][1] ~^ image[1][9] + signed_kernel[0][2] ~^ image[1][10] + signed_kernel[0][3] ~^ image[1][11] + signed_kernel[0][4] ~^ image[1][12] + signed_kernel[1][0] ~^ image[2][8] + signed_kernel[1][1] ~^ image[2][9] + signed_kernel[1][2] ~^ image[2][10] + signed_kernel[1][3] ~^ image[2][11] + signed_kernel[1][4] ~^ image[2][12] + signed_kernel[2][0] ~^ image[3][8] + signed_kernel[2][1] ~^ image[3][9] + signed_kernel[2][2] ~^ image[3][10] + signed_kernel[2][3] ~^ image[3][11] + signed_kernel[2][4] ~^ image[3][12] + signed_kernel[3][0] ~^ image[4][8] + signed_kernel[3][1] ~^ image[4][9] + signed_kernel[3][2] ~^ image[4][10] + signed_kernel[3][3] ~^ image[4][11] + signed_kernel[3][4] ~^ image[4][12] + signed_kernel[4][0] ~^ image[5][8] + signed_kernel[4][1] ~^ image[5][9] + signed_kernel[4][2] ~^ image[5][10] + signed_kernel[4][3] ~^ image[5][11] + signed_kernel[4][4] ~^ image[5][12];
assign xor_sum[1][9] = signed_kernel[0][0] ~^ image[1][9] + signed_kernel[0][1] ~^ image[1][10] + signed_kernel[0][2] ~^ image[1][11] + signed_kernel[0][3] ~^ image[1][12] + signed_kernel[0][4] ~^ image[1][13] + signed_kernel[1][0] ~^ image[2][9] + signed_kernel[1][1] ~^ image[2][10] + signed_kernel[1][2] ~^ image[2][11] + signed_kernel[1][3] ~^ image[2][12] + signed_kernel[1][4] ~^ image[2][13] + signed_kernel[2][0] ~^ image[3][9] + signed_kernel[2][1] ~^ image[3][10] + signed_kernel[2][2] ~^ image[3][11] + signed_kernel[2][3] ~^ image[3][12] + signed_kernel[2][4] ~^ image[3][13] + signed_kernel[3][0] ~^ image[4][9] + signed_kernel[3][1] ~^ image[4][10] + signed_kernel[3][2] ~^ image[4][11] + signed_kernel[3][3] ~^ image[4][12] + signed_kernel[3][4] ~^ image[4][13] + signed_kernel[4][0] ~^ image[5][9] + signed_kernel[4][1] ~^ image[5][10] + signed_kernel[4][2] ~^ image[5][11] + signed_kernel[4][3] ~^ image[5][12] + signed_kernel[4][4] ~^ image[5][13];
assign xor_sum[1][10] = signed_kernel[0][0] ~^ image[1][10] + signed_kernel[0][1] ~^ image[1][11] + signed_kernel[0][2] ~^ image[1][12] + signed_kernel[0][3] ~^ image[1][13] + signed_kernel[0][4] ~^ image[1][14] + signed_kernel[1][0] ~^ image[2][10] + signed_kernel[1][1] ~^ image[2][11] + signed_kernel[1][2] ~^ image[2][12] + signed_kernel[1][3] ~^ image[2][13] + signed_kernel[1][4] ~^ image[2][14] + signed_kernel[2][0] ~^ image[3][10] + signed_kernel[2][1] ~^ image[3][11] + signed_kernel[2][2] ~^ image[3][12] + signed_kernel[2][3] ~^ image[3][13] + signed_kernel[2][4] ~^ image[3][14] + signed_kernel[3][0] ~^ image[4][10] + signed_kernel[3][1] ~^ image[4][11] + signed_kernel[3][2] ~^ image[4][12] + signed_kernel[3][3] ~^ image[4][13] + signed_kernel[3][4] ~^ image[4][14] + signed_kernel[4][0] ~^ image[5][10] + signed_kernel[4][1] ~^ image[5][11] + signed_kernel[4][2] ~^ image[5][12] + signed_kernel[4][3] ~^ image[5][13] + signed_kernel[4][4] ~^ image[5][14];
assign xor_sum[1][11] = signed_kernel[0][0] ~^ image[1][11] + signed_kernel[0][1] ~^ image[1][12] + signed_kernel[0][2] ~^ image[1][13] + signed_kernel[0][3] ~^ image[1][14] + signed_kernel[0][4] ~^ image[1][15] + signed_kernel[1][0] ~^ image[2][11] + signed_kernel[1][1] ~^ image[2][12] + signed_kernel[1][2] ~^ image[2][13] + signed_kernel[1][3] ~^ image[2][14] + signed_kernel[1][4] ~^ image[2][15] + signed_kernel[2][0] ~^ image[3][11] + signed_kernel[2][1] ~^ image[3][12] + signed_kernel[2][2] ~^ image[3][13] + signed_kernel[2][3] ~^ image[3][14] + signed_kernel[2][4] ~^ image[3][15] + signed_kernel[3][0] ~^ image[4][11] + signed_kernel[3][1] ~^ image[4][12] + signed_kernel[3][2] ~^ image[4][13] + signed_kernel[3][3] ~^ image[4][14] + signed_kernel[3][4] ~^ image[4][15] + signed_kernel[4][0] ~^ image[5][11] + signed_kernel[4][1] ~^ image[5][12] + signed_kernel[4][2] ~^ image[5][13] + signed_kernel[4][3] ~^ image[5][14] + signed_kernel[4][4] ~^ image[5][15];
assign xor_sum[1][12] = signed_kernel[0][0] ~^ image[1][12] + signed_kernel[0][1] ~^ image[1][13] + signed_kernel[0][2] ~^ image[1][14] + signed_kernel[0][3] ~^ image[1][15] + signed_kernel[0][4] ~^ image[1][16] + signed_kernel[1][0] ~^ image[2][12] + signed_kernel[1][1] ~^ image[2][13] + signed_kernel[1][2] ~^ image[2][14] + signed_kernel[1][3] ~^ image[2][15] + signed_kernel[1][4] ~^ image[2][16] + signed_kernel[2][0] ~^ image[3][12] + signed_kernel[2][1] ~^ image[3][13] + signed_kernel[2][2] ~^ image[3][14] + signed_kernel[2][3] ~^ image[3][15] + signed_kernel[2][4] ~^ image[3][16] + signed_kernel[3][0] ~^ image[4][12] + signed_kernel[3][1] ~^ image[4][13] + signed_kernel[3][2] ~^ image[4][14] + signed_kernel[3][3] ~^ image[4][15] + signed_kernel[3][4] ~^ image[4][16] + signed_kernel[4][0] ~^ image[5][12] + signed_kernel[4][1] ~^ image[5][13] + signed_kernel[4][2] ~^ image[5][14] + signed_kernel[4][3] ~^ image[5][15] + signed_kernel[4][4] ~^ image[5][16];
assign xor_sum[1][13] = signed_kernel[0][0] ~^ image[1][13] + signed_kernel[0][1] ~^ image[1][14] + signed_kernel[0][2] ~^ image[1][15] + signed_kernel[0][3] ~^ image[1][16] + signed_kernel[0][4] ~^ image[1][17] + signed_kernel[1][0] ~^ image[2][13] + signed_kernel[1][1] ~^ image[2][14] + signed_kernel[1][2] ~^ image[2][15] + signed_kernel[1][3] ~^ image[2][16] + signed_kernel[1][4] ~^ image[2][17] + signed_kernel[2][0] ~^ image[3][13] + signed_kernel[2][1] ~^ image[3][14] + signed_kernel[2][2] ~^ image[3][15] + signed_kernel[2][3] ~^ image[3][16] + signed_kernel[2][4] ~^ image[3][17] + signed_kernel[3][0] ~^ image[4][13] + signed_kernel[3][1] ~^ image[4][14] + signed_kernel[3][2] ~^ image[4][15] + signed_kernel[3][3] ~^ image[4][16] + signed_kernel[3][4] ~^ image[4][17] + signed_kernel[4][0] ~^ image[5][13] + signed_kernel[4][1] ~^ image[5][14] + signed_kernel[4][2] ~^ image[5][15] + signed_kernel[4][3] ~^ image[5][16] + signed_kernel[4][4] ~^ image[5][17];
assign xor_sum[1][14] = signed_kernel[0][0] ~^ image[1][14] + signed_kernel[0][1] ~^ image[1][15] + signed_kernel[0][2] ~^ image[1][16] + signed_kernel[0][3] ~^ image[1][17] + signed_kernel[0][4] ~^ image[1][18] + signed_kernel[1][0] ~^ image[2][14] + signed_kernel[1][1] ~^ image[2][15] + signed_kernel[1][2] ~^ image[2][16] + signed_kernel[1][3] ~^ image[2][17] + signed_kernel[1][4] ~^ image[2][18] + signed_kernel[2][0] ~^ image[3][14] + signed_kernel[2][1] ~^ image[3][15] + signed_kernel[2][2] ~^ image[3][16] + signed_kernel[2][3] ~^ image[3][17] + signed_kernel[2][4] ~^ image[3][18] + signed_kernel[3][0] ~^ image[4][14] + signed_kernel[3][1] ~^ image[4][15] + signed_kernel[3][2] ~^ image[4][16] + signed_kernel[3][3] ~^ image[4][17] + signed_kernel[3][4] ~^ image[4][18] + signed_kernel[4][0] ~^ image[5][14] + signed_kernel[4][1] ~^ image[5][15] + signed_kernel[4][2] ~^ image[5][16] + signed_kernel[4][3] ~^ image[5][17] + signed_kernel[4][4] ~^ image[5][18];
assign xor_sum[1][15] = signed_kernel[0][0] ~^ image[1][15] + signed_kernel[0][1] ~^ image[1][16] + signed_kernel[0][2] ~^ image[1][17] + signed_kernel[0][3] ~^ image[1][18] + signed_kernel[0][4] ~^ image[1][19] + signed_kernel[1][0] ~^ image[2][15] + signed_kernel[1][1] ~^ image[2][16] + signed_kernel[1][2] ~^ image[2][17] + signed_kernel[1][3] ~^ image[2][18] + signed_kernel[1][4] ~^ image[2][19] + signed_kernel[2][0] ~^ image[3][15] + signed_kernel[2][1] ~^ image[3][16] + signed_kernel[2][2] ~^ image[3][17] + signed_kernel[2][3] ~^ image[3][18] + signed_kernel[2][4] ~^ image[3][19] + signed_kernel[3][0] ~^ image[4][15] + signed_kernel[3][1] ~^ image[4][16] + signed_kernel[3][2] ~^ image[4][17] + signed_kernel[3][3] ~^ image[4][18] + signed_kernel[3][4] ~^ image[4][19] + signed_kernel[4][0] ~^ image[5][15] + signed_kernel[4][1] ~^ image[5][16] + signed_kernel[4][2] ~^ image[5][17] + signed_kernel[4][3] ~^ image[5][18] + signed_kernel[4][4] ~^ image[5][19];
assign xor_sum[1][16] = signed_kernel[0][0] ~^ image[1][16] + signed_kernel[0][1] ~^ image[1][17] + signed_kernel[0][2] ~^ image[1][18] + signed_kernel[0][3] ~^ image[1][19] + signed_kernel[0][4] ~^ image[1][20] + signed_kernel[1][0] ~^ image[2][16] + signed_kernel[1][1] ~^ image[2][17] + signed_kernel[1][2] ~^ image[2][18] + signed_kernel[1][3] ~^ image[2][19] + signed_kernel[1][4] ~^ image[2][20] + signed_kernel[2][0] ~^ image[3][16] + signed_kernel[2][1] ~^ image[3][17] + signed_kernel[2][2] ~^ image[3][18] + signed_kernel[2][3] ~^ image[3][19] + signed_kernel[2][4] ~^ image[3][20] + signed_kernel[3][0] ~^ image[4][16] + signed_kernel[3][1] ~^ image[4][17] + signed_kernel[3][2] ~^ image[4][18] + signed_kernel[3][3] ~^ image[4][19] + signed_kernel[3][4] ~^ image[4][20] + signed_kernel[4][0] ~^ image[5][16] + signed_kernel[4][1] ~^ image[5][17] + signed_kernel[4][2] ~^ image[5][18] + signed_kernel[4][3] ~^ image[5][19] + signed_kernel[4][4] ~^ image[5][20];
assign xor_sum[1][17] = signed_kernel[0][0] ~^ image[1][17] + signed_kernel[0][1] ~^ image[1][18] + signed_kernel[0][2] ~^ image[1][19] + signed_kernel[0][3] ~^ image[1][20] + signed_kernel[0][4] ~^ image[1][21] + signed_kernel[1][0] ~^ image[2][17] + signed_kernel[1][1] ~^ image[2][18] + signed_kernel[1][2] ~^ image[2][19] + signed_kernel[1][3] ~^ image[2][20] + signed_kernel[1][4] ~^ image[2][21] + signed_kernel[2][0] ~^ image[3][17] + signed_kernel[2][1] ~^ image[3][18] + signed_kernel[2][2] ~^ image[3][19] + signed_kernel[2][3] ~^ image[3][20] + signed_kernel[2][4] ~^ image[3][21] + signed_kernel[3][0] ~^ image[4][17] + signed_kernel[3][1] ~^ image[4][18] + signed_kernel[3][2] ~^ image[4][19] + signed_kernel[3][3] ~^ image[4][20] + signed_kernel[3][4] ~^ image[4][21] + signed_kernel[4][0] ~^ image[5][17] + signed_kernel[4][1] ~^ image[5][18] + signed_kernel[4][2] ~^ image[5][19] + signed_kernel[4][3] ~^ image[5][20] + signed_kernel[4][4] ~^ image[5][21];
assign xor_sum[1][18] = signed_kernel[0][0] ~^ image[1][18] + signed_kernel[0][1] ~^ image[1][19] + signed_kernel[0][2] ~^ image[1][20] + signed_kernel[0][3] ~^ image[1][21] + signed_kernel[0][4] ~^ image[1][22] + signed_kernel[1][0] ~^ image[2][18] + signed_kernel[1][1] ~^ image[2][19] + signed_kernel[1][2] ~^ image[2][20] + signed_kernel[1][3] ~^ image[2][21] + signed_kernel[1][4] ~^ image[2][22] + signed_kernel[2][0] ~^ image[3][18] + signed_kernel[2][1] ~^ image[3][19] + signed_kernel[2][2] ~^ image[3][20] + signed_kernel[2][3] ~^ image[3][21] + signed_kernel[2][4] ~^ image[3][22] + signed_kernel[3][0] ~^ image[4][18] + signed_kernel[3][1] ~^ image[4][19] + signed_kernel[3][2] ~^ image[4][20] + signed_kernel[3][3] ~^ image[4][21] + signed_kernel[3][4] ~^ image[4][22] + signed_kernel[4][0] ~^ image[5][18] + signed_kernel[4][1] ~^ image[5][19] + signed_kernel[4][2] ~^ image[5][20] + signed_kernel[4][3] ~^ image[5][21] + signed_kernel[4][4] ~^ image[5][22];
assign xor_sum[1][19] = signed_kernel[0][0] ~^ image[1][19] + signed_kernel[0][1] ~^ image[1][20] + signed_kernel[0][2] ~^ image[1][21] + signed_kernel[0][3] ~^ image[1][22] + signed_kernel[0][4] ~^ image[1][23] + signed_kernel[1][0] ~^ image[2][19] + signed_kernel[1][1] ~^ image[2][20] + signed_kernel[1][2] ~^ image[2][21] + signed_kernel[1][3] ~^ image[2][22] + signed_kernel[1][4] ~^ image[2][23] + signed_kernel[2][0] ~^ image[3][19] + signed_kernel[2][1] ~^ image[3][20] + signed_kernel[2][2] ~^ image[3][21] + signed_kernel[2][3] ~^ image[3][22] + signed_kernel[2][4] ~^ image[3][23] + signed_kernel[3][0] ~^ image[4][19] + signed_kernel[3][1] ~^ image[4][20] + signed_kernel[3][2] ~^ image[4][21] + signed_kernel[3][3] ~^ image[4][22] + signed_kernel[3][4] ~^ image[4][23] + signed_kernel[4][0] ~^ image[5][19] + signed_kernel[4][1] ~^ image[5][20] + signed_kernel[4][2] ~^ image[5][21] + signed_kernel[4][3] ~^ image[5][22] + signed_kernel[4][4] ~^ image[5][23];
assign xor_sum[1][20] = signed_kernel[0][0] ~^ image[1][20] + signed_kernel[0][1] ~^ image[1][21] + signed_kernel[0][2] ~^ image[1][22] + signed_kernel[0][3] ~^ image[1][23] + signed_kernel[0][4] ~^ image[1][24] + signed_kernel[1][0] ~^ image[2][20] + signed_kernel[1][1] ~^ image[2][21] + signed_kernel[1][2] ~^ image[2][22] + signed_kernel[1][3] ~^ image[2][23] + signed_kernel[1][4] ~^ image[2][24] + signed_kernel[2][0] ~^ image[3][20] + signed_kernel[2][1] ~^ image[3][21] + signed_kernel[2][2] ~^ image[3][22] + signed_kernel[2][3] ~^ image[3][23] + signed_kernel[2][4] ~^ image[3][24] + signed_kernel[3][0] ~^ image[4][20] + signed_kernel[3][1] ~^ image[4][21] + signed_kernel[3][2] ~^ image[4][22] + signed_kernel[3][3] ~^ image[4][23] + signed_kernel[3][4] ~^ image[4][24] + signed_kernel[4][0] ~^ image[5][20] + signed_kernel[4][1] ~^ image[5][21] + signed_kernel[4][2] ~^ image[5][22] + signed_kernel[4][3] ~^ image[5][23] + signed_kernel[4][4] ~^ image[5][24];
assign xor_sum[1][21] = signed_kernel[0][0] ~^ image[1][21] + signed_kernel[0][1] ~^ image[1][22] + signed_kernel[0][2] ~^ image[1][23] + signed_kernel[0][3] ~^ image[1][24] + signed_kernel[0][4] ~^ image[1][25] + signed_kernel[1][0] ~^ image[2][21] + signed_kernel[1][1] ~^ image[2][22] + signed_kernel[1][2] ~^ image[2][23] + signed_kernel[1][3] ~^ image[2][24] + signed_kernel[1][4] ~^ image[2][25] + signed_kernel[2][0] ~^ image[3][21] + signed_kernel[2][1] ~^ image[3][22] + signed_kernel[2][2] ~^ image[3][23] + signed_kernel[2][3] ~^ image[3][24] + signed_kernel[2][4] ~^ image[3][25] + signed_kernel[3][0] ~^ image[4][21] + signed_kernel[3][1] ~^ image[4][22] + signed_kernel[3][2] ~^ image[4][23] + signed_kernel[3][3] ~^ image[4][24] + signed_kernel[3][4] ~^ image[4][25] + signed_kernel[4][0] ~^ image[5][21] + signed_kernel[4][1] ~^ image[5][22] + signed_kernel[4][2] ~^ image[5][23] + signed_kernel[4][3] ~^ image[5][24] + signed_kernel[4][4] ~^ image[5][25];
assign xor_sum[1][22] = signed_kernel[0][0] ~^ image[1][22] + signed_kernel[0][1] ~^ image[1][23] + signed_kernel[0][2] ~^ image[1][24] + signed_kernel[0][3] ~^ image[1][25] + signed_kernel[0][4] ~^ image[1][26] + signed_kernel[1][0] ~^ image[2][22] + signed_kernel[1][1] ~^ image[2][23] + signed_kernel[1][2] ~^ image[2][24] + signed_kernel[1][3] ~^ image[2][25] + signed_kernel[1][4] ~^ image[2][26] + signed_kernel[2][0] ~^ image[3][22] + signed_kernel[2][1] ~^ image[3][23] + signed_kernel[2][2] ~^ image[3][24] + signed_kernel[2][3] ~^ image[3][25] + signed_kernel[2][4] ~^ image[3][26] + signed_kernel[3][0] ~^ image[4][22] + signed_kernel[3][1] ~^ image[4][23] + signed_kernel[3][2] ~^ image[4][24] + signed_kernel[3][3] ~^ image[4][25] + signed_kernel[3][4] ~^ image[4][26] + signed_kernel[4][0] ~^ image[5][22] + signed_kernel[4][1] ~^ image[5][23] + signed_kernel[4][2] ~^ image[5][24] + signed_kernel[4][3] ~^ image[5][25] + signed_kernel[4][4] ~^ image[5][26];
assign xor_sum[1][23] = signed_kernel[0][0] ~^ image[1][23] + signed_kernel[0][1] ~^ image[1][24] + signed_kernel[0][2] ~^ image[1][25] + signed_kernel[0][3] ~^ image[1][26] + signed_kernel[0][4] ~^ image[1][27] + signed_kernel[1][0] ~^ image[2][23] + signed_kernel[1][1] ~^ image[2][24] + signed_kernel[1][2] ~^ image[2][25] + signed_kernel[1][3] ~^ image[2][26] + signed_kernel[1][4] ~^ image[2][27] + signed_kernel[2][0] ~^ image[3][23] + signed_kernel[2][1] ~^ image[3][24] + signed_kernel[2][2] ~^ image[3][25] + signed_kernel[2][3] ~^ image[3][26] + signed_kernel[2][4] ~^ image[3][27] + signed_kernel[3][0] ~^ image[4][23] + signed_kernel[3][1] ~^ image[4][24] + signed_kernel[3][2] ~^ image[4][25] + signed_kernel[3][3] ~^ image[4][26] + signed_kernel[3][4] ~^ image[4][27] + signed_kernel[4][0] ~^ image[5][23] + signed_kernel[4][1] ~^ image[5][24] + signed_kernel[4][2] ~^ image[5][25] + signed_kernel[4][3] ~^ image[5][26] + signed_kernel[4][4] ~^ image[5][27];
assign xor_sum[2][0] = signed_kernel[0][0] ~^ image[2][0] + signed_kernel[0][1] ~^ image[2][1] + signed_kernel[0][2] ~^ image[2][2] + signed_kernel[0][3] ~^ image[2][3] + signed_kernel[0][4] ~^ image[2][4] + signed_kernel[1][0] ~^ image[3][0] + signed_kernel[1][1] ~^ image[3][1] + signed_kernel[1][2] ~^ image[3][2] + signed_kernel[1][3] ~^ image[3][3] + signed_kernel[1][4] ~^ image[3][4] + signed_kernel[2][0] ~^ image[4][0] + signed_kernel[2][1] ~^ image[4][1] + signed_kernel[2][2] ~^ image[4][2] + signed_kernel[2][3] ~^ image[4][3] + signed_kernel[2][4] ~^ image[4][4] + signed_kernel[3][0] ~^ image[5][0] + signed_kernel[3][1] ~^ image[5][1] + signed_kernel[3][2] ~^ image[5][2] + signed_kernel[3][3] ~^ image[5][3] + signed_kernel[3][4] ~^ image[5][4] + signed_kernel[4][0] ~^ image[6][0] + signed_kernel[4][1] ~^ image[6][1] + signed_kernel[4][2] ~^ image[6][2] + signed_kernel[4][3] ~^ image[6][3] + signed_kernel[4][4] ~^ image[6][4];
assign xor_sum[2][1] = signed_kernel[0][0] ~^ image[2][1] + signed_kernel[0][1] ~^ image[2][2] + signed_kernel[0][2] ~^ image[2][3] + signed_kernel[0][3] ~^ image[2][4] + signed_kernel[0][4] ~^ image[2][5] + signed_kernel[1][0] ~^ image[3][1] + signed_kernel[1][1] ~^ image[3][2] + signed_kernel[1][2] ~^ image[3][3] + signed_kernel[1][3] ~^ image[3][4] + signed_kernel[1][4] ~^ image[3][5] + signed_kernel[2][0] ~^ image[4][1] + signed_kernel[2][1] ~^ image[4][2] + signed_kernel[2][2] ~^ image[4][3] + signed_kernel[2][3] ~^ image[4][4] + signed_kernel[2][4] ~^ image[4][5] + signed_kernel[3][0] ~^ image[5][1] + signed_kernel[3][1] ~^ image[5][2] + signed_kernel[3][2] ~^ image[5][3] + signed_kernel[3][3] ~^ image[5][4] + signed_kernel[3][4] ~^ image[5][5] + signed_kernel[4][0] ~^ image[6][1] + signed_kernel[4][1] ~^ image[6][2] + signed_kernel[4][2] ~^ image[6][3] + signed_kernel[4][3] ~^ image[6][4] + signed_kernel[4][4] ~^ image[6][5];
assign xor_sum[2][2] = signed_kernel[0][0] ~^ image[2][2] + signed_kernel[0][1] ~^ image[2][3] + signed_kernel[0][2] ~^ image[2][4] + signed_kernel[0][3] ~^ image[2][5] + signed_kernel[0][4] ~^ image[2][6] + signed_kernel[1][0] ~^ image[3][2] + signed_kernel[1][1] ~^ image[3][3] + signed_kernel[1][2] ~^ image[3][4] + signed_kernel[1][3] ~^ image[3][5] + signed_kernel[1][4] ~^ image[3][6] + signed_kernel[2][0] ~^ image[4][2] + signed_kernel[2][1] ~^ image[4][3] + signed_kernel[2][2] ~^ image[4][4] + signed_kernel[2][3] ~^ image[4][5] + signed_kernel[2][4] ~^ image[4][6] + signed_kernel[3][0] ~^ image[5][2] + signed_kernel[3][1] ~^ image[5][3] + signed_kernel[3][2] ~^ image[5][4] + signed_kernel[3][3] ~^ image[5][5] + signed_kernel[3][4] ~^ image[5][6] + signed_kernel[4][0] ~^ image[6][2] + signed_kernel[4][1] ~^ image[6][3] + signed_kernel[4][2] ~^ image[6][4] + signed_kernel[4][3] ~^ image[6][5] + signed_kernel[4][4] ~^ image[6][6];
assign xor_sum[2][3] = signed_kernel[0][0] ~^ image[2][3] + signed_kernel[0][1] ~^ image[2][4] + signed_kernel[0][2] ~^ image[2][5] + signed_kernel[0][3] ~^ image[2][6] + signed_kernel[0][4] ~^ image[2][7] + signed_kernel[1][0] ~^ image[3][3] + signed_kernel[1][1] ~^ image[3][4] + signed_kernel[1][2] ~^ image[3][5] + signed_kernel[1][3] ~^ image[3][6] + signed_kernel[1][4] ~^ image[3][7] + signed_kernel[2][0] ~^ image[4][3] + signed_kernel[2][1] ~^ image[4][4] + signed_kernel[2][2] ~^ image[4][5] + signed_kernel[2][3] ~^ image[4][6] + signed_kernel[2][4] ~^ image[4][7] + signed_kernel[3][0] ~^ image[5][3] + signed_kernel[3][1] ~^ image[5][4] + signed_kernel[3][2] ~^ image[5][5] + signed_kernel[3][3] ~^ image[5][6] + signed_kernel[3][4] ~^ image[5][7] + signed_kernel[4][0] ~^ image[6][3] + signed_kernel[4][1] ~^ image[6][4] + signed_kernel[4][2] ~^ image[6][5] + signed_kernel[4][3] ~^ image[6][6] + signed_kernel[4][4] ~^ image[6][7];
assign xor_sum[2][4] = signed_kernel[0][0] ~^ image[2][4] + signed_kernel[0][1] ~^ image[2][5] + signed_kernel[0][2] ~^ image[2][6] + signed_kernel[0][3] ~^ image[2][7] + signed_kernel[0][4] ~^ image[2][8] + signed_kernel[1][0] ~^ image[3][4] + signed_kernel[1][1] ~^ image[3][5] + signed_kernel[1][2] ~^ image[3][6] + signed_kernel[1][3] ~^ image[3][7] + signed_kernel[1][4] ~^ image[3][8] + signed_kernel[2][0] ~^ image[4][4] + signed_kernel[2][1] ~^ image[4][5] + signed_kernel[2][2] ~^ image[4][6] + signed_kernel[2][3] ~^ image[4][7] + signed_kernel[2][4] ~^ image[4][8] + signed_kernel[3][0] ~^ image[5][4] + signed_kernel[3][1] ~^ image[5][5] + signed_kernel[3][2] ~^ image[5][6] + signed_kernel[3][3] ~^ image[5][7] + signed_kernel[3][4] ~^ image[5][8] + signed_kernel[4][0] ~^ image[6][4] + signed_kernel[4][1] ~^ image[6][5] + signed_kernel[4][2] ~^ image[6][6] + signed_kernel[4][3] ~^ image[6][7] + signed_kernel[4][4] ~^ image[6][8];
assign xor_sum[2][5] = signed_kernel[0][0] ~^ image[2][5] + signed_kernel[0][1] ~^ image[2][6] + signed_kernel[0][2] ~^ image[2][7] + signed_kernel[0][3] ~^ image[2][8] + signed_kernel[0][4] ~^ image[2][9] + signed_kernel[1][0] ~^ image[3][5] + signed_kernel[1][1] ~^ image[3][6] + signed_kernel[1][2] ~^ image[3][7] + signed_kernel[1][3] ~^ image[3][8] + signed_kernel[1][4] ~^ image[3][9] + signed_kernel[2][0] ~^ image[4][5] + signed_kernel[2][1] ~^ image[4][6] + signed_kernel[2][2] ~^ image[4][7] + signed_kernel[2][3] ~^ image[4][8] + signed_kernel[2][4] ~^ image[4][9] + signed_kernel[3][0] ~^ image[5][5] + signed_kernel[3][1] ~^ image[5][6] + signed_kernel[3][2] ~^ image[5][7] + signed_kernel[3][3] ~^ image[5][8] + signed_kernel[3][4] ~^ image[5][9] + signed_kernel[4][0] ~^ image[6][5] + signed_kernel[4][1] ~^ image[6][6] + signed_kernel[4][2] ~^ image[6][7] + signed_kernel[4][3] ~^ image[6][8] + signed_kernel[4][4] ~^ image[6][9];
assign xor_sum[2][6] = signed_kernel[0][0] ~^ image[2][6] + signed_kernel[0][1] ~^ image[2][7] + signed_kernel[0][2] ~^ image[2][8] + signed_kernel[0][3] ~^ image[2][9] + signed_kernel[0][4] ~^ image[2][10] + signed_kernel[1][0] ~^ image[3][6] + signed_kernel[1][1] ~^ image[3][7] + signed_kernel[1][2] ~^ image[3][8] + signed_kernel[1][3] ~^ image[3][9] + signed_kernel[1][4] ~^ image[3][10] + signed_kernel[2][0] ~^ image[4][6] + signed_kernel[2][1] ~^ image[4][7] + signed_kernel[2][2] ~^ image[4][8] + signed_kernel[2][3] ~^ image[4][9] + signed_kernel[2][4] ~^ image[4][10] + signed_kernel[3][0] ~^ image[5][6] + signed_kernel[3][1] ~^ image[5][7] + signed_kernel[3][2] ~^ image[5][8] + signed_kernel[3][3] ~^ image[5][9] + signed_kernel[3][4] ~^ image[5][10] + signed_kernel[4][0] ~^ image[6][6] + signed_kernel[4][1] ~^ image[6][7] + signed_kernel[4][2] ~^ image[6][8] + signed_kernel[4][3] ~^ image[6][9] + signed_kernel[4][4] ~^ image[6][10];
assign xor_sum[2][7] = signed_kernel[0][0] ~^ image[2][7] + signed_kernel[0][1] ~^ image[2][8] + signed_kernel[0][2] ~^ image[2][9] + signed_kernel[0][3] ~^ image[2][10] + signed_kernel[0][4] ~^ image[2][11] + signed_kernel[1][0] ~^ image[3][7] + signed_kernel[1][1] ~^ image[3][8] + signed_kernel[1][2] ~^ image[3][9] + signed_kernel[1][3] ~^ image[3][10] + signed_kernel[1][4] ~^ image[3][11] + signed_kernel[2][0] ~^ image[4][7] + signed_kernel[2][1] ~^ image[4][8] + signed_kernel[2][2] ~^ image[4][9] + signed_kernel[2][3] ~^ image[4][10] + signed_kernel[2][4] ~^ image[4][11] + signed_kernel[3][0] ~^ image[5][7] + signed_kernel[3][1] ~^ image[5][8] + signed_kernel[3][2] ~^ image[5][9] + signed_kernel[3][3] ~^ image[5][10] + signed_kernel[3][4] ~^ image[5][11] + signed_kernel[4][0] ~^ image[6][7] + signed_kernel[4][1] ~^ image[6][8] + signed_kernel[4][2] ~^ image[6][9] + signed_kernel[4][3] ~^ image[6][10] + signed_kernel[4][4] ~^ image[6][11];
assign xor_sum[2][8] = signed_kernel[0][0] ~^ image[2][8] + signed_kernel[0][1] ~^ image[2][9] + signed_kernel[0][2] ~^ image[2][10] + signed_kernel[0][3] ~^ image[2][11] + signed_kernel[0][4] ~^ image[2][12] + signed_kernel[1][0] ~^ image[3][8] + signed_kernel[1][1] ~^ image[3][9] + signed_kernel[1][2] ~^ image[3][10] + signed_kernel[1][3] ~^ image[3][11] + signed_kernel[1][4] ~^ image[3][12] + signed_kernel[2][0] ~^ image[4][8] + signed_kernel[2][1] ~^ image[4][9] + signed_kernel[2][2] ~^ image[4][10] + signed_kernel[2][3] ~^ image[4][11] + signed_kernel[2][4] ~^ image[4][12] + signed_kernel[3][0] ~^ image[5][8] + signed_kernel[3][1] ~^ image[5][9] + signed_kernel[3][2] ~^ image[5][10] + signed_kernel[3][3] ~^ image[5][11] + signed_kernel[3][4] ~^ image[5][12] + signed_kernel[4][0] ~^ image[6][8] + signed_kernel[4][1] ~^ image[6][9] + signed_kernel[4][2] ~^ image[6][10] + signed_kernel[4][3] ~^ image[6][11] + signed_kernel[4][4] ~^ image[6][12];
assign xor_sum[2][9] = signed_kernel[0][0] ~^ image[2][9] + signed_kernel[0][1] ~^ image[2][10] + signed_kernel[0][2] ~^ image[2][11] + signed_kernel[0][3] ~^ image[2][12] + signed_kernel[0][4] ~^ image[2][13] + signed_kernel[1][0] ~^ image[3][9] + signed_kernel[1][1] ~^ image[3][10] + signed_kernel[1][2] ~^ image[3][11] + signed_kernel[1][3] ~^ image[3][12] + signed_kernel[1][4] ~^ image[3][13] + signed_kernel[2][0] ~^ image[4][9] + signed_kernel[2][1] ~^ image[4][10] + signed_kernel[2][2] ~^ image[4][11] + signed_kernel[2][3] ~^ image[4][12] + signed_kernel[2][4] ~^ image[4][13] + signed_kernel[3][0] ~^ image[5][9] + signed_kernel[3][1] ~^ image[5][10] + signed_kernel[3][2] ~^ image[5][11] + signed_kernel[3][3] ~^ image[5][12] + signed_kernel[3][4] ~^ image[5][13] + signed_kernel[4][0] ~^ image[6][9] + signed_kernel[4][1] ~^ image[6][10] + signed_kernel[4][2] ~^ image[6][11] + signed_kernel[4][3] ~^ image[6][12] + signed_kernel[4][4] ~^ image[6][13];
assign xor_sum[2][10] = signed_kernel[0][0] ~^ image[2][10] + signed_kernel[0][1] ~^ image[2][11] + signed_kernel[0][2] ~^ image[2][12] + signed_kernel[0][3] ~^ image[2][13] + signed_kernel[0][4] ~^ image[2][14] + signed_kernel[1][0] ~^ image[3][10] + signed_kernel[1][1] ~^ image[3][11] + signed_kernel[1][2] ~^ image[3][12] + signed_kernel[1][3] ~^ image[3][13] + signed_kernel[1][4] ~^ image[3][14] + signed_kernel[2][0] ~^ image[4][10] + signed_kernel[2][1] ~^ image[4][11] + signed_kernel[2][2] ~^ image[4][12] + signed_kernel[2][3] ~^ image[4][13] + signed_kernel[2][4] ~^ image[4][14] + signed_kernel[3][0] ~^ image[5][10] + signed_kernel[3][1] ~^ image[5][11] + signed_kernel[3][2] ~^ image[5][12] + signed_kernel[3][3] ~^ image[5][13] + signed_kernel[3][4] ~^ image[5][14] + signed_kernel[4][0] ~^ image[6][10] + signed_kernel[4][1] ~^ image[6][11] + signed_kernel[4][2] ~^ image[6][12] + signed_kernel[4][3] ~^ image[6][13] + signed_kernel[4][4] ~^ image[6][14];
assign xor_sum[2][11] = signed_kernel[0][0] ~^ image[2][11] + signed_kernel[0][1] ~^ image[2][12] + signed_kernel[0][2] ~^ image[2][13] + signed_kernel[0][3] ~^ image[2][14] + signed_kernel[0][4] ~^ image[2][15] + signed_kernel[1][0] ~^ image[3][11] + signed_kernel[1][1] ~^ image[3][12] + signed_kernel[1][2] ~^ image[3][13] + signed_kernel[1][3] ~^ image[3][14] + signed_kernel[1][4] ~^ image[3][15] + signed_kernel[2][0] ~^ image[4][11] + signed_kernel[2][1] ~^ image[4][12] + signed_kernel[2][2] ~^ image[4][13] + signed_kernel[2][3] ~^ image[4][14] + signed_kernel[2][4] ~^ image[4][15] + signed_kernel[3][0] ~^ image[5][11] + signed_kernel[3][1] ~^ image[5][12] + signed_kernel[3][2] ~^ image[5][13] + signed_kernel[3][3] ~^ image[5][14] + signed_kernel[3][4] ~^ image[5][15] + signed_kernel[4][0] ~^ image[6][11] + signed_kernel[4][1] ~^ image[6][12] + signed_kernel[4][2] ~^ image[6][13] + signed_kernel[4][3] ~^ image[6][14] + signed_kernel[4][4] ~^ image[6][15];
assign xor_sum[2][12] = signed_kernel[0][0] ~^ image[2][12] + signed_kernel[0][1] ~^ image[2][13] + signed_kernel[0][2] ~^ image[2][14] + signed_kernel[0][3] ~^ image[2][15] + signed_kernel[0][4] ~^ image[2][16] + signed_kernel[1][0] ~^ image[3][12] + signed_kernel[1][1] ~^ image[3][13] + signed_kernel[1][2] ~^ image[3][14] + signed_kernel[1][3] ~^ image[3][15] + signed_kernel[1][4] ~^ image[3][16] + signed_kernel[2][0] ~^ image[4][12] + signed_kernel[2][1] ~^ image[4][13] + signed_kernel[2][2] ~^ image[4][14] + signed_kernel[2][3] ~^ image[4][15] + signed_kernel[2][4] ~^ image[4][16] + signed_kernel[3][0] ~^ image[5][12] + signed_kernel[3][1] ~^ image[5][13] + signed_kernel[3][2] ~^ image[5][14] + signed_kernel[3][3] ~^ image[5][15] + signed_kernel[3][4] ~^ image[5][16] + signed_kernel[4][0] ~^ image[6][12] + signed_kernel[4][1] ~^ image[6][13] + signed_kernel[4][2] ~^ image[6][14] + signed_kernel[4][3] ~^ image[6][15] + signed_kernel[4][4] ~^ image[6][16];
assign xor_sum[2][13] = signed_kernel[0][0] ~^ image[2][13] + signed_kernel[0][1] ~^ image[2][14] + signed_kernel[0][2] ~^ image[2][15] + signed_kernel[0][3] ~^ image[2][16] + signed_kernel[0][4] ~^ image[2][17] + signed_kernel[1][0] ~^ image[3][13] + signed_kernel[1][1] ~^ image[3][14] + signed_kernel[1][2] ~^ image[3][15] + signed_kernel[1][3] ~^ image[3][16] + signed_kernel[1][4] ~^ image[3][17] + signed_kernel[2][0] ~^ image[4][13] + signed_kernel[2][1] ~^ image[4][14] + signed_kernel[2][2] ~^ image[4][15] + signed_kernel[2][3] ~^ image[4][16] + signed_kernel[2][4] ~^ image[4][17] + signed_kernel[3][0] ~^ image[5][13] + signed_kernel[3][1] ~^ image[5][14] + signed_kernel[3][2] ~^ image[5][15] + signed_kernel[3][3] ~^ image[5][16] + signed_kernel[3][4] ~^ image[5][17] + signed_kernel[4][0] ~^ image[6][13] + signed_kernel[4][1] ~^ image[6][14] + signed_kernel[4][2] ~^ image[6][15] + signed_kernel[4][3] ~^ image[6][16] + signed_kernel[4][4] ~^ image[6][17];
assign xor_sum[2][14] = signed_kernel[0][0] ~^ image[2][14] + signed_kernel[0][1] ~^ image[2][15] + signed_kernel[0][2] ~^ image[2][16] + signed_kernel[0][3] ~^ image[2][17] + signed_kernel[0][4] ~^ image[2][18] + signed_kernel[1][0] ~^ image[3][14] + signed_kernel[1][1] ~^ image[3][15] + signed_kernel[1][2] ~^ image[3][16] + signed_kernel[1][3] ~^ image[3][17] + signed_kernel[1][4] ~^ image[3][18] + signed_kernel[2][0] ~^ image[4][14] + signed_kernel[2][1] ~^ image[4][15] + signed_kernel[2][2] ~^ image[4][16] + signed_kernel[2][3] ~^ image[4][17] + signed_kernel[2][4] ~^ image[4][18] + signed_kernel[3][0] ~^ image[5][14] + signed_kernel[3][1] ~^ image[5][15] + signed_kernel[3][2] ~^ image[5][16] + signed_kernel[3][3] ~^ image[5][17] + signed_kernel[3][4] ~^ image[5][18] + signed_kernel[4][0] ~^ image[6][14] + signed_kernel[4][1] ~^ image[6][15] + signed_kernel[4][2] ~^ image[6][16] + signed_kernel[4][3] ~^ image[6][17] + signed_kernel[4][4] ~^ image[6][18];
assign xor_sum[2][15] = signed_kernel[0][0] ~^ image[2][15] + signed_kernel[0][1] ~^ image[2][16] + signed_kernel[0][2] ~^ image[2][17] + signed_kernel[0][3] ~^ image[2][18] + signed_kernel[0][4] ~^ image[2][19] + signed_kernel[1][0] ~^ image[3][15] + signed_kernel[1][1] ~^ image[3][16] + signed_kernel[1][2] ~^ image[3][17] + signed_kernel[1][3] ~^ image[3][18] + signed_kernel[1][4] ~^ image[3][19] + signed_kernel[2][0] ~^ image[4][15] + signed_kernel[2][1] ~^ image[4][16] + signed_kernel[2][2] ~^ image[4][17] + signed_kernel[2][3] ~^ image[4][18] + signed_kernel[2][4] ~^ image[4][19] + signed_kernel[3][0] ~^ image[5][15] + signed_kernel[3][1] ~^ image[5][16] + signed_kernel[3][2] ~^ image[5][17] + signed_kernel[3][3] ~^ image[5][18] + signed_kernel[3][4] ~^ image[5][19] + signed_kernel[4][0] ~^ image[6][15] + signed_kernel[4][1] ~^ image[6][16] + signed_kernel[4][2] ~^ image[6][17] + signed_kernel[4][3] ~^ image[6][18] + signed_kernel[4][4] ~^ image[6][19];
assign xor_sum[2][16] = signed_kernel[0][0] ~^ image[2][16] + signed_kernel[0][1] ~^ image[2][17] + signed_kernel[0][2] ~^ image[2][18] + signed_kernel[0][3] ~^ image[2][19] + signed_kernel[0][4] ~^ image[2][20] + signed_kernel[1][0] ~^ image[3][16] + signed_kernel[1][1] ~^ image[3][17] + signed_kernel[1][2] ~^ image[3][18] + signed_kernel[1][3] ~^ image[3][19] + signed_kernel[1][4] ~^ image[3][20] + signed_kernel[2][0] ~^ image[4][16] + signed_kernel[2][1] ~^ image[4][17] + signed_kernel[2][2] ~^ image[4][18] + signed_kernel[2][3] ~^ image[4][19] + signed_kernel[2][4] ~^ image[4][20] + signed_kernel[3][0] ~^ image[5][16] + signed_kernel[3][1] ~^ image[5][17] + signed_kernel[3][2] ~^ image[5][18] + signed_kernel[3][3] ~^ image[5][19] + signed_kernel[3][4] ~^ image[5][20] + signed_kernel[4][0] ~^ image[6][16] + signed_kernel[4][1] ~^ image[6][17] + signed_kernel[4][2] ~^ image[6][18] + signed_kernel[4][3] ~^ image[6][19] + signed_kernel[4][4] ~^ image[6][20];
assign xor_sum[2][17] = signed_kernel[0][0] ~^ image[2][17] + signed_kernel[0][1] ~^ image[2][18] + signed_kernel[0][2] ~^ image[2][19] + signed_kernel[0][3] ~^ image[2][20] + signed_kernel[0][4] ~^ image[2][21] + signed_kernel[1][0] ~^ image[3][17] + signed_kernel[1][1] ~^ image[3][18] + signed_kernel[1][2] ~^ image[3][19] + signed_kernel[1][3] ~^ image[3][20] + signed_kernel[1][4] ~^ image[3][21] + signed_kernel[2][0] ~^ image[4][17] + signed_kernel[2][1] ~^ image[4][18] + signed_kernel[2][2] ~^ image[4][19] + signed_kernel[2][3] ~^ image[4][20] + signed_kernel[2][4] ~^ image[4][21] + signed_kernel[3][0] ~^ image[5][17] + signed_kernel[3][1] ~^ image[5][18] + signed_kernel[3][2] ~^ image[5][19] + signed_kernel[3][3] ~^ image[5][20] + signed_kernel[3][4] ~^ image[5][21] + signed_kernel[4][0] ~^ image[6][17] + signed_kernel[4][1] ~^ image[6][18] + signed_kernel[4][2] ~^ image[6][19] + signed_kernel[4][3] ~^ image[6][20] + signed_kernel[4][4] ~^ image[6][21];
assign xor_sum[2][18] = signed_kernel[0][0] ~^ image[2][18] + signed_kernel[0][1] ~^ image[2][19] + signed_kernel[0][2] ~^ image[2][20] + signed_kernel[0][3] ~^ image[2][21] + signed_kernel[0][4] ~^ image[2][22] + signed_kernel[1][0] ~^ image[3][18] + signed_kernel[1][1] ~^ image[3][19] + signed_kernel[1][2] ~^ image[3][20] + signed_kernel[1][3] ~^ image[3][21] + signed_kernel[1][4] ~^ image[3][22] + signed_kernel[2][0] ~^ image[4][18] + signed_kernel[2][1] ~^ image[4][19] + signed_kernel[2][2] ~^ image[4][20] + signed_kernel[2][3] ~^ image[4][21] + signed_kernel[2][4] ~^ image[4][22] + signed_kernel[3][0] ~^ image[5][18] + signed_kernel[3][1] ~^ image[5][19] + signed_kernel[3][2] ~^ image[5][20] + signed_kernel[3][3] ~^ image[5][21] + signed_kernel[3][4] ~^ image[5][22] + signed_kernel[4][0] ~^ image[6][18] + signed_kernel[4][1] ~^ image[6][19] + signed_kernel[4][2] ~^ image[6][20] + signed_kernel[4][3] ~^ image[6][21] + signed_kernel[4][4] ~^ image[6][22];
assign xor_sum[2][19] = signed_kernel[0][0] ~^ image[2][19] + signed_kernel[0][1] ~^ image[2][20] + signed_kernel[0][2] ~^ image[2][21] + signed_kernel[0][3] ~^ image[2][22] + signed_kernel[0][4] ~^ image[2][23] + signed_kernel[1][0] ~^ image[3][19] + signed_kernel[1][1] ~^ image[3][20] + signed_kernel[1][2] ~^ image[3][21] + signed_kernel[1][3] ~^ image[3][22] + signed_kernel[1][4] ~^ image[3][23] + signed_kernel[2][0] ~^ image[4][19] + signed_kernel[2][1] ~^ image[4][20] + signed_kernel[2][2] ~^ image[4][21] + signed_kernel[2][3] ~^ image[4][22] + signed_kernel[2][4] ~^ image[4][23] + signed_kernel[3][0] ~^ image[5][19] + signed_kernel[3][1] ~^ image[5][20] + signed_kernel[3][2] ~^ image[5][21] + signed_kernel[3][3] ~^ image[5][22] + signed_kernel[3][4] ~^ image[5][23] + signed_kernel[4][0] ~^ image[6][19] + signed_kernel[4][1] ~^ image[6][20] + signed_kernel[4][2] ~^ image[6][21] + signed_kernel[4][3] ~^ image[6][22] + signed_kernel[4][4] ~^ image[6][23];
assign xor_sum[2][20] = signed_kernel[0][0] ~^ image[2][20] + signed_kernel[0][1] ~^ image[2][21] + signed_kernel[0][2] ~^ image[2][22] + signed_kernel[0][3] ~^ image[2][23] + signed_kernel[0][4] ~^ image[2][24] + signed_kernel[1][0] ~^ image[3][20] + signed_kernel[1][1] ~^ image[3][21] + signed_kernel[1][2] ~^ image[3][22] + signed_kernel[1][3] ~^ image[3][23] + signed_kernel[1][4] ~^ image[3][24] + signed_kernel[2][0] ~^ image[4][20] + signed_kernel[2][1] ~^ image[4][21] + signed_kernel[2][2] ~^ image[4][22] + signed_kernel[2][3] ~^ image[4][23] + signed_kernel[2][4] ~^ image[4][24] + signed_kernel[3][0] ~^ image[5][20] + signed_kernel[3][1] ~^ image[5][21] + signed_kernel[3][2] ~^ image[5][22] + signed_kernel[3][3] ~^ image[5][23] + signed_kernel[3][4] ~^ image[5][24] + signed_kernel[4][0] ~^ image[6][20] + signed_kernel[4][1] ~^ image[6][21] + signed_kernel[4][2] ~^ image[6][22] + signed_kernel[4][3] ~^ image[6][23] + signed_kernel[4][4] ~^ image[6][24];
assign xor_sum[2][21] = signed_kernel[0][0] ~^ image[2][21] + signed_kernel[0][1] ~^ image[2][22] + signed_kernel[0][2] ~^ image[2][23] + signed_kernel[0][3] ~^ image[2][24] + signed_kernel[0][4] ~^ image[2][25] + signed_kernel[1][0] ~^ image[3][21] + signed_kernel[1][1] ~^ image[3][22] + signed_kernel[1][2] ~^ image[3][23] + signed_kernel[1][3] ~^ image[3][24] + signed_kernel[1][4] ~^ image[3][25] + signed_kernel[2][0] ~^ image[4][21] + signed_kernel[2][1] ~^ image[4][22] + signed_kernel[2][2] ~^ image[4][23] + signed_kernel[2][3] ~^ image[4][24] + signed_kernel[2][4] ~^ image[4][25] + signed_kernel[3][0] ~^ image[5][21] + signed_kernel[3][1] ~^ image[5][22] + signed_kernel[3][2] ~^ image[5][23] + signed_kernel[3][3] ~^ image[5][24] + signed_kernel[3][4] ~^ image[5][25] + signed_kernel[4][0] ~^ image[6][21] + signed_kernel[4][1] ~^ image[6][22] + signed_kernel[4][2] ~^ image[6][23] + signed_kernel[4][3] ~^ image[6][24] + signed_kernel[4][4] ~^ image[6][25];
assign xor_sum[2][22] = signed_kernel[0][0] ~^ image[2][22] + signed_kernel[0][1] ~^ image[2][23] + signed_kernel[0][2] ~^ image[2][24] + signed_kernel[0][3] ~^ image[2][25] + signed_kernel[0][4] ~^ image[2][26] + signed_kernel[1][0] ~^ image[3][22] + signed_kernel[1][1] ~^ image[3][23] + signed_kernel[1][2] ~^ image[3][24] + signed_kernel[1][3] ~^ image[3][25] + signed_kernel[1][4] ~^ image[3][26] + signed_kernel[2][0] ~^ image[4][22] + signed_kernel[2][1] ~^ image[4][23] + signed_kernel[2][2] ~^ image[4][24] + signed_kernel[2][3] ~^ image[4][25] + signed_kernel[2][4] ~^ image[4][26] + signed_kernel[3][0] ~^ image[5][22] + signed_kernel[3][1] ~^ image[5][23] + signed_kernel[3][2] ~^ image[5][24] + signed_kernel[3][3] ~^ image[5][25] + signed_kernel[3][4] ~^ image[5][26] + signed_kernel[4][0] ~^ image[6][22] + signed_kernel[4][1] ~^ image[6][23] + signed_kernel[4][2] ~^ image[6][24] + signed_kernel[4][3] ~^ image[6][25] + signed_kernel[4][4] ~^ image[6][26];
assign xor_sum[2][23] = signed_kernel[0][0] ~^ image[2][23] + signed_kernel[0][1] ~^ image[2][24] + signed_kernel[0][2] ~^ image[2][25] + signed_kernel[0][3] ~^ image[2][26] + signed_kernel[0][4] ~^ image[2][27] + signed_kernel[1][0] ~^ image[3][23] + signed_kernel[1][1] ~^ image[3][24] + signed_kernel[1][2] ~^ image[3][25] + signed_kernel[1][3] ~^ image[3][26] + signed_kernel[1][4] ~^ image[3][27] + signed_kernel[2][0] ~^ image[4][23] + signed_kernel[2][1] ~^ image[4][24] + signed_kernel[2][2] ~^ image[4][25] + signed_kernel[2][3] ~^ image[4][26] + signed_kernel[2][4] ~^ image[4][27] + signed_kernel[3][0] ~^ image[5][23] + signed_kernel[3][1] ~^ image[5][24] + signed_kernel[3][2] ~^ image[5][25] + signed_kernel[3][3] ~^ image[5][26] + signed_kernel[3][4] ~^ image[5][27] + signed_kernel[4][0] ~^ image[6][23] + signed_kernel[4][1] ~^ image[6][24] + signed_kernel[4][2] ~^ image[6][25] + signed_kernel[4][3] ~^ image[6][26] + signed_kernel[4][4] ~^ image[6][27];
assign xor_sum[3][0] = signed_kernel[0][0] ~^ image[3][0] + signed_kernel[0][1] ~^ image[3][1] + signed_kernel[0][2] ~^ image[3][2] + signed_kernel[0][3] ~^ image[3][3] + signed_kernel[0][4] ~^ image[3][4] + signed_kernel[1][0] ~^ image[4][0] + signed_kernel[1][1] ~^ image[4][1] + signed_kernel[1][2] ~^ image[4][2] + signed_kernel[1][3] ~^ image[4][3] + signed_kernel[1][4] ~^ image[4][4] + signed_kernel[2][0] ~^ image[5][0] + signed_kernel[2][1] ~^ image[5][1] + signed_kernel[2][2] ~^ image[5][2] + signed_kernel[2][3] ~^ image[5][3] + signed_kernel[2][4] ~^ image[5][4] + signed_kernel[3][0] ~^ image[6][0] + signed_kernel[3][1] ~^ image[6][1] + signed_kernel[3][2] ~^ image[6][2] + signed_kernel[3][3] ~^ image[6][3] + signed_kernel[3][4] ~^ image[6][4] + signed_kernel[4][0] ~^ image[7][0] + signed_kernel[4][1] ~^ image[7][1] + signed_kernel[4][2] ~^ image[7][2] + signed_kernel[4][3] ~^ image[7][3] + signed_kernel[4][4] ~^ image[7][4];
assign xor_sum[3][1] = signed_kernel[0][0] ~^ image[3][1] + signed_kernel[0][1] ~^ image[3][2] + signed_kernel[0][2] ~^ image[3][3] + signed_kernel[0][3] ~^ image[3][4] + signed_kernel[0][4] ~^ image[3][5] + signed_kernel[1][0] ~^ image[4][1] + signed_kernel[1][1] ~^ image[4][2] + signed_kernel[1][2] ~^ image[4][3] + signed_kernel[1][3] ~^ image[4][4] + signed_kernel[1][4] ~^ image[4][5] + signed_kernel[2][0] ~^ image[5][1] + signed_kernel[2][1] ~^ image[5][2] + signed_kernel[2][2] ~^ image[5][3] + signed_kernel[2][3] ~^ image[5][4] + signed_kernel[2][4] ~^ image[5][5] + signed_kernel[3][0] ~^ image[6][1] + signed_kernel[3][1] ~^ image[6][2] + signed_kernel[3][2] ~^ image[6][3] + signed_kernel[3][3] ~^ image[6][4] + signed_kernel[3][4] ~^ image[6][5] + signed_kernel[4][0] ~^ image[7][1] + signed_kernel[4][1] ~^ image[7][2] + signed_kernel[4][2] ~^ image[7][3] + signed_kernel[4][3] ~^ image[7][4] + signed_kernel[4][4] ~^ image[7][5];
assign xor_sum[3][2] = signed_kernel[0][0] ~^ image[3][2] + signed_kernel[0][1] ~^ image[3][3] + signed_kernel[0][2] ~^ image[3][4] + signed_kernel[0][3] ~^ image[3][5] + signed_kernel[0][4] ~^ image[3][6] + signed_kernel[1][0] ~^ image[4][2] + signed_kernel[1][1] ~^ image[4][3] + signed_kernel[1][2] ~^ image[4][4] + signed_kernel[1][3] ~^ image[4][5] + signed_kernel[1][4] ~^ image[4][6] + signed_kernel[2][0] ~^ image[5][2] + signed_kernel[2][1] ~^ image[5][3] + signed_kernel[2][2] ~^ image[5][4] + signed_kernel[2][3] ~^ image[5][5] + signed_kernel[2][4] ~^ image[5][6] + signed_kernel[3][0] ~^ image[6][2] + signed_kernel[3][1] ~^ image[6][3] + signed_kernel[3][2] ~^ image[6][4] + signed_kernel[3][3] ~^ image[6][5] + signed_kernel[3][4] ~^ image[6][6] + signed_kernel[4][0] ~^ image[7][2] + signed_kernel[4][1] ~^ image[7][3] + signed_kernel[4][2] ~^ image[7][4] + signed_kernel[4][3] ~^ image[7][5] + signed_kernel[4][4] ~^ image[7][6];
assign xor_sum[3][3] = signed_kernel[0][0] ~^ image[3][3] + signed_kernel[0][1] ~^ image[3][4] + signed_kernel[0][2] ~^ image[3][5] + signed_kernel[0][3] ~^ image[3][6] + signed_kernel[0][4] ~^ image[3][7] + signed_kernel[1][0] ~^ image[4][3] + signed_kernel[1][1] ~^ image[4][4] + signed_kernel[1][2] ~^ image[4][5] + signed_kernel[1][3] ~^ image[4][6] + signed_kernel[1][4] ~^ image[4][7] + signed_kernel[2][0] ~^ image[5][3] + signed_kernel[2][1] ~^ image[5][4] + signed_kernel[2][2] ~^ image[5][5] + signed_kernel[2][3] ~^ image[5][6] + signed_kernel[2][4] ~^ image[5][7] + signed_kernel[3][0] ~^ image[6][3] + signed_kernel[3][1] ~^ image[6][4] + signed_kernel[3][2] ~^ image[6][5] + signed_kernel[3][3] ~^ image[6][6] + signed_kernel[3][4] ~^ image[6][7] + signed_kernel[4][0] ~^ image[7][3] + signed_kernel[4][1] ~^ image[7][4] + signed_kernel[4][2] ~^ image[7][5] + signed_kernel[4][3] ~^ image[7][6] + signed_kernel[4][4] ~^ image[7][7];
assign xor_sum[3][4] = signed_kernel[0][0] ~^ image[3][4] + signed_kernel[0][1] ~^ image[3][5] + signed_kernel[0][2] ~^ image[3][6] + signed_kernel[0][3] ~^ image[3][7] + signed_kernel[0][4] ~^ image[3][8] + signed_kernel[1][0] ~^ image[4][4] + signed_kernel[1][1] ~^ image[4][5] + signed_kernel[1][2] ~^ image[4][6] + signed_kernel[1][3] ~^ image[4][7] + signed_kernel[1][4] ~^ image[4][8] + signed_kernel[2][0] ~^ image[5][4] + signed_kernel[2][1] ~^ image[5][5] + signed_kernel[2][2] ~^ image[5][6] + signed_kernel[2][3] ~^ image[5][7] + signed_kernel[2][4] ~^ image[5][8] + signed_kernel[3][0] ~^ image[6][4] + signed_kernel[3][1] ~^ image[6][5] + signed_kernel[3][2] ~^ image[6][6] + signed_kernel[3][3] ~^ image[6][7] + signed_kernel[3][4] ~^ image[6][8] + signed_kernel[4][0] ~^ image[7][4] + signed_kernel[4][1] ~^ image[7][5] + signed_kernel[4][2] ~^ image[7][6] + signed_kernel[4][3] ~^ image[7][7] + signed_kernel[4][4] ~^ image[7][8];
assign xor_sum[3][5] = signed_kernel[0][0] ~^ image[3][5] + signed_kernel[0][1] ~^ image[3][6] + signed_kernel[0][2] ~^ image[3][7] + signed_kernel[0][3] ~^ image[3][8] + signed_kernel[0][4] ~^ image[3][9] + signed_kernel[1][0] ~^ image[4][5] + signed_kernel[1][1] ~^ image[4][6] + signed_kernel[1][2] ~^ image[4][7] + signed_kernel[1][3] ~^ image[4][8] + signed_kernel[1][4] ~^ image[4][9] + signed_kernel[2][0] ~^ image[5][5] + signed_kernel[2][1] ~^ image[5][6] + signed_kernel[2][2] ~^ image[5][7] + signed_kernel[2][3] ~^ image[5][8] + signed_kernel[2][4] ~^ image[5][9] + signed_kernel[3][0] ~^ image[6][5] + signed_kernel[3][1] ~^ image[6][6] + signed_kernel[3][2] ~^ image[6][7] + signed_kernel[3][3] ~^ image[6][8] + signed_kernel[3][4] ~^ image[6][9] + signed_kernel[4][0] ~^ image[7][5] + signed_kernel[4][1] ~^ image[7][6] + signed_kernel[4][2] ~^ image[7][7] + signed_kernel[4][3] ~^ image[7][8] + signed_kernel[4][4] ~^ image[7][9];
assign xor_sum[3][6] = signed_kernel[0][0] ~^ image[3][6] + signed_kernel[0][1] ~^ image[3][7] + signed_kernel[0][2] ~^ image[3][8] + signed_kernel[0][3] ~^ image[3][9] + signed_kernel[0][4] ~^ image[3][10] + signed_kernel[1][0] ~^ image[4][6] + signed_kernel[1][1] ~^ image[4][7] + signed_kernel[1][2] ~^ image[4][8] + signed_kernel[1][3] ~^ image[4][9] + signed_kernel[1][4] ~^ image[4][10] + signed_kernel[2][0] ~^ image[5][6] + signed_kernel[2][1] ~^ image[5][7] + signed_kernel[2][2] ~^ image[5][8] + signed_kernel[2][3] ~^ image[5][9] + signed_kernel[2][4] ~^ image[5][10] + signed_kernel[3][0] ~^ image[6][6] + signed_kernel[3][1] ~^ image[6][7] + signed_kernel[3][2] ~^ image[6][8] + signed_kernel[3][3] ~^ image[6][9] + signed_kernel[3][4] ~^ image[6][10] + signed_kernel[4][0] ~^ image[7][6] + signed_kernel[4][1] ~^ image[7][7] + signed_kernel[4][2] ~^ image[7][8] + signed_kernel[4][3] ~^ image[7][9] + signed_kernel[4][4] ~^ image[7][10];
assign xor_sum[3][7] = signed_kernel[0][0] ~^ image[3][7] + signed_kernel[0][1] ~^ image[3][8] + signed_kernel[0][2] ~^ image[3][9] + signed_kernel[0][3] ~^ image[3][10] + signed_kernel[0][4] ~^ image[3][11] + signed_kernel[1][0] ~^ image[4][7] + signed_kernel[1][1] ~^ image[4][8] + signed_kernel[1][2] ~^ image[4][9] + signed_kernel[1][3] ~^ image[4][10] + signed_kernel[1][4] ~^ image[4][11] + signed_kernel[2][0] ~^ image[5][7] + signed_kernel[2][1] ~^ image[5][8] + signed_kernel[2][2] ~^ image[5][9] + signed_kernel[2][3] ~^ image[5][10] + signed_kernel[2][4] ~^ image[5][11] + signed_kernel[3][0] ~^ image[6][7] + signed_kernel[3][1] ~^ image[6][8] + signed_kernel[3][2] ~^ image[6][9] + signed_kernel[3][3] ~^ image[6][10] + signed_kernel[3][4] ~^ image[6][11] + signed_kernel[4][0] ~^ image[7][7] + signed_kernel[4][1] ~^ image[7][8] + signed_kernel[4][2] ~^ image[7][9] + signed_kernel[4][3] ~^ image[7][10] + signed_kernel[4][4] ~^ image[7][11];
assign xor_sum[3][8] = signed_kernel[0][0] ~^ image[3][8] + signed_kernel[0][1] ~^ image[3][9] + signed_kernel[0][2] ~^ image[3][10] + signed_kernel[0][3] ~^ image[3][11] + signed_kernel[0][4] ~^ image[3][12] + signed_kernel[1][0] ~^ image[4][8] + signed_kernel[1][1] ~^ image[4][9] + signed_kernel[1][2] ~^ image[4][10] + signed_kernel[1][3] ~^ image[4][11] + signed_kernel[1][4] ~^ image[4][12] + signed_kernel[2][0] ~^ image[5][8] + signed_kernel[2][1] ~^ image[5][9] + signed_kernel[2][2] ~^ image[5][10] + signed_kernel[2][3] ~^ image[5][11] + signed_kernel[2][4] ~^ image[5][12] + signed_kernel[3][0] ~^ image[6][8] + signed_kernel[3][1] ~^ image[6][9] + signed_kernel[3][2] ~^ image[6][10] + signed_kernel[3][3] ~^ image[6][11] + signed_kernel[3][4] ~^ image[6][12] + signed_kernel[4][0] ~^ image[7][8] + signed_kernel[4][1] ~^ image[7][9] + signed_kernel[4][2] ~^ image[7][10] + signed_kernel[4][3] ~^ image[7][11] + signed_kernel[4][4] ~^ image[7][12];
assign xor_sum[3][9] = signed_kernel[0][0] ~^ image[3][9] + signed_kernel[0][1] ~^ image[3][10] + signed_kernel[0][2] ~^ image[3][11] + signed_kernel[0][3] ~^ image[3][12] + signed_kernel[0][4] ~^ image[3][13] + signed_kernel[1][0] ~^ image[4][9] + signed_kernel[1][1] ~^ image[4][10] + signed_kernel[1][2] ~^ image[4][11] + signed_kernel[1][3] ~^ image[4][12] + signed_kernel[1][4] ~^ image[4][13] + signed_kernel[2][0] ~^ image[5][9] + signed_kernel[2][1] ~^ image[5][10] + signed_kernel[2][2] ~^ image[5][11] + signed_kernel[2][3] ~^ image[5][12] + signed_kernel[2][4] ~^ image[5][13] + signed_kernel[3][0] ~^ image[6][9] + signed_kernel[3][1] ~^ image[6][10] + signed_kernel[3][2] ~^ image[6][11] + signed_kernel[3][3] ~^ image[6][12] + signed_kernel[3][4] ~^ image[6][13] + signed_kernel[4][0] ~^ image[7][9] + signed_kernel[4][1] ~^ image[7][10] + signed_kernel[4][2] ~^ image[7][11] + signed_kernel[4][3] ~^ image[7][12] + signed_kernel[4][4] ~^ image[7][13];
assign xor_sum[3][10] = signed_kernel[0][0] ~^ image[3][10] + signed_kernel[0][1] ~^ image[3][11] + signed_kernel[0][2] ~^ image[3][12] + signed_kernel[0][3] ~^ image[3][13] + signed_kernel[0][4] ~^ image[3][14] + signed_kernel[1][0] ~^ image[4][10] + signed_kernel[1][1] ~^ image[4][11] + signed_kernel[1][2] ~^ image[4][12] + signed_kernel[1][3] ~^ image[4][13] + signed_kernel[1][4] ~^ image[4][14] + signed_kernel[2][0] ~^ image[5][10] + signed_kernel[2][1] ~^ image[5][11] + signed_kernel[2][2] ~^ image[5][12] + signed_kernel[2][3] ~^ image[5][13] + signed_kernel[2][4] ~^ image[5][14] + signed_kernel[3][0] ~^ image[6][10] + signed_kernel[3][1] ~^ image[6][11] + signed_kernel[3][2] ~^ image[6][12] + signed_kernel[3][3] ~^ image[6][13] + signed_kernel[3][4] ~^ image[6][14] + signed_kernel[4][0] ~^ image[7][10] + signed_kernel[4][1] ~^ image[7][11] + signed_kernel[4][2] ~^ image[7][12] + signed_kernel[4][3] ~^ image[7][13] + signed_kernel[4][4] ~^ image[7][14];
assign xor_sum[3][11] = signed_kernel[0][0] ~^ image[3][11] + signed_kernel[0][1] ~^ image[3][12] + signed_kernel[0][2] ~^ image[3][13] + signed_kernel[0][3] ~^ image[3][14] + signed_kernel[0][4] ~^ image[3][15] + signed_kernel[1][0] ~^ image[4][11] + signed_kernel[1][1] ~^ image[4][12] + signed_kernel[1][2] ~^ image[4][13] + signed_kernel[1][3] ~^ image[4][14] + signed_kernel[1][4] ~^ image[4][15] + signed_kernel[2][0] ~^ image[5][11] + signed_kernel[2][1] ~^ image[5][12] + signed_kernel[2][2] ~^ image[5][13] + signed_kernel[2][3] ~^ image[5][14] + signed_kernel[2][4] ~^ image[5][15] + signed_kernel[3][0] ~^ image[6][11] + signed_kernel[3][1] ~^ image[6][12] + signed_kernel[3][2] ~^ image[6][13] + signed_kernel[3][3] ~^ image[6][14] + signed_kernel[3][4] ~^ image[6][15] + signed_kernel[4][0] ~^ image[7][11] + signed_kernel[4][1] ~^ image[7][12] + signed_kernel[4][2] ~^ image[7][13] + signed_kernel[4][3] ~^ image[7][14] + signed_kernel[4][4] ~^ image[7][15];
assign xor_sum[3][12] = signed_kernel[0][0] ~^ image[3][12] + signed_kernel[0][1] ~^ image[3][13] + signed_kernel[0][2] ~^ image[3][14] + signed_kernel[0][3] ~^ image[3][15] + signed_kernel[0][4] ~^ image[3][16] + signed_kernel[1][0] ~^ image[4][12] + signed_kernel[1][1] ~^ image[4][13] + signed_kernel[1][2] ~^ image[4][14] + signed_kernel[1][3] ~^ image[4][15] + signed_kernel[1][4] ~^ image[4][16] + signed_kernel[2][0] ~^ image[5][12] + signed_kernel[2][1] ~^ image[5][13] + signed_kernel[2][2] ~^ image[5][14] + signed_kernel[2][3] ~^ image[5][15] + signed_kernel[2][4] ~^ image[5][16] + signed_kernel[3][0] ~^ image[6][12] + signed_kernel[3][1] ~^ image[6][13] + signed_kernel[3][2] ~^ image[6][14] + signed_kernel[3][3] ~^ image[6][15] + signed_kernel[3][4] ~^ image[6][16] + signed_kernel[4][0] ~^ image[7][12] + signed_kernel[4][1] ~^ image[7][13] + signed_kernel[4][2] ~^ image[7][14] + signed_kernel[4][3] ~^ image[7][15] + signed_kernel[4][4] ~^ image[7][16];
assign xor_sum[3][13] = signed_kernel[0][0] ~^ image[3][13] + signed_kernel[0][1] ~^ image[3][14] + signed_kernel[0][2] ~^ image[3][15] + signed_kernel[0][3] ~^ image[3][16] + signed_kernel[0][4] ~^ image[3][17] + signed_kernel[1][0] ~^ image[4][13] + signed_kernel[1][1] ~^ image[4][14] + signed_kernel[1][2] ~^ image[4][15] + signed_kernel[1][3] ~^ image[4][16] + signed_kernel[1][4] ~^ image[4][17] + signed_kernel[2][0] ~^ image[5][13] + signed_kernel[2][1] ~^ image[5][14] + signed_kernel[2][2] ~^ image[5][15] + signed_kernel[2][3] ~^ image[5][16] + signed_kernel[2][4] ~^ image[5][17] + signed_kernel[3][0] ~^ image[6][13] + signed_kernel[3][1] ~^ image[6][14] + signed_kernel[3][2] ~^ image[6][15] + signed_kernel[3][3] ~^ image[6][16] + signed_kernel[3][4] ~^ image[6][17] + signed_kernel[4][0] ~^ image[7][13] + signed_kernel[4][1] ~^ image[7][14] + signed_kernel[4][2] ~^ image[7][15] + signed_kernel[4][3] ~^ image[7][16] + signed_kernel[4][4] ~^ image[7][17];
assign xor_sum[3][14] = signed_kernel[0][0] ~^ image[3][14] + signed_kernel[0][1] ~^ image[3][15] + signed_kernel[0][2] ~^ image[3][16] + signed_kernel[0][3] ~^ image[3][17] + signed_kernel[0][4] ~^ image[3][18] + signed_kernel[1][0] ~^ image[4][14] + signed_kernel[1][1] ~^ image[4][15] + signed_kernel[1][2] ~^ image[4][16] + signed_kernel[1][3] ~^ image[4][17] + signed_kernel[1][4] ~^ image[4][18] + signed_kernel[2][0] ~^ image[5][14] + signed_kernel[2][1] ~^ image[5][15] + signed_kernel[2][2] ~^ image[5][16] + signed_kernel[2][3] ~^ image[5][17] + signed_kernel[2][4] ~^ image[5][18] + signed_kernel[3][0] ~^ image[6][14] + signed_kernel[3][1] ~^ image[6][15] + signed_kernel[3][2] ~^ image[6][16] + signed_kernel[3][3] ~^ image[6][17] + signed_kernel[3][4] ~^ image[6][18] + signed_kernel[4][0] ~^ image[7][14] + signed_kernel[4][1] ~^ image[7][15] + signed_kernel[4][2] ~^ image[7][16] + signed_kernel[4][3] ~^ image[7][17] + signed_kernel[4][4] ~^ image[7][18];
assign xor_sum[3][15] = signed_kernel[0][0] ~^ image[3][15] + signed_kernel[0][1] ~^ image[3][16] + signed_kernel[0][2] ~^ image[3][17] + signed_kernel[0][3] ~^ image[3][18] + signed_kernel[0][4] ~^ image[3][19] + signed_kernel[1][0] ~^ image[4][15] + signed_kernel[1][1] ~^ image[4][16] + signed_kernel[1][2] ~^ image[4][17] + signed_kernel[1][3] ~^ image[4][18] + signed_kernel[1][4] ~^ image[4][19] + signed_kernel[2][0] ~^ image[5][15] + signed_kernel[2][1] ~^ image[5][16] + signed_kernel[2][2] ~^ image[5][17] + signed_kernel[2][3] ~^ image[5][18] + signed_kernel[2][4] ~^ image[5][19] + signed_kernel[3][0] ~^ image[6][15] + signed_kernel[3][1] ~^ image[6][16] + signed_kernel[3][2] ~^ image[6][17] + signed_kernel[3][3] ~^ image[6][18] + signed_kernel[3][4] ~^ image[6][19] + signed_kernel[4][0] ~^ image[7][15] + signed_kernel[4][1] ~^ image[7][16] + signed_kernel[4][2] ~^ image[7][17] + signed_kernel[4][3] ~^ image[7][18] + signed_kernel[4][4] ~^ image[7][19];
assign xor_sum[3][16] = signed_kernel[0][0] ~^ image[3][16] + signed_kernel[0][1] ~^ image[3][17] + signed_kernel[0][2] ~^ image[3][18] + signed_kernel[0][3] ~^ image[3][19] + signed_kernel[0][4] ~^ image[3][20] + signed_kernel[1][0] ~^ image[4][16] + signed_kernel[1][1] ~^ image[4][17] + signed_kernel[1][2] ~^ image[4][18] + signed_kernel[1][3] ~^ image[4][19] + signed_kernel[1][4] ~^ image[4][20] + signed_kernel[2][0] ~^ image[5][16] + signed_kernel[2][1] ~^ image[5][17] + signed_kernel[2][2] ~^ image[5][18] + signed_kernel[2][3] ~^ image[5][19] + signed_kernel[2][4] ~^ image[5][20] + signed_kernel[3][0] ~^ image[6][16] + signed_kernel[3][1] ~^ image[6][17] + signed_kernel[3][2] ~^ image[6][18] + signed_kernel[3][3] ~^ image[6][19] + signed_kernel[3][4] ~^ image[6][20] + signed_kernel[4][0] ~^ image[7][16] + signed_kernel[4][1] ~^ image[7][17] + signed_kernel[4][2] ~^ image[7][18] + signed_kernel[4][3] ~^ image[7][19] + signed_kernel[4][4] ~^ image[7][20];
assign xor_sum[3][17] = signed_kernel[0][0] ~^ image[3][17] + signed_kernel[0][1] ~^ image[3][18] + signed_kernel[0][2] ~^ image[3][19] + signed_kernel[0][3] ~^ image[3][20] + signed_kernel[0][4] ~^ image[3][21] + signed_kernel[1][0] ~^ image[4][17] + signed_kernel[1][1] ~^ image[4][18] + signed_kernel[1][2] ~^ image[4][19] + signed_kernel[1][3] ~^ image[4][20] + signed_kernel[1][4] ~^ image[4][21] + signed_kernel[2][0] ~^ image[5][17] + signed_kernel[2][1] ~^ image[5][18] + signed_kernel[2][2] ~^ image[5][19] + signed_kernel[2][3] ~^ image[5][20] + signed_kernel[2][4] ~^ image[5][21] + signed_kernel[3][0] ~^ image[6][17] + signed_kernel[3][1] ~^ image[6][18] + signed_kernel[3][2] ~^ image[6][19] + signed_kernel[3][3] ~^ image[6][20] + signed_kernel[3][4] ~^ image[6][21] + signed_kernel[4][0] ~^ image[7][17] + signed_kernel[4][1] ~^ image[7][18] + signed_kernel[4][2] ~^ image[7][19] + signed_kernel[4][3] ~^ image[7][20] + signed_kernel[4][4] ~^ image[7][21];
assign xor_sum[3][18] = signed_kernel[0][0] ~^ image[3][18] + signed_kernel[0][1] ~^ image[3][19] + signed_kernel[0][2] ~^ image[3][20] + signed_kernel[0][3] ~^ image[3][21] + signed_kernel[0][4] ~^ image[3][22] + signed_kernel[1][0] ~^ image[4][18] + signed_kernel[1][1] ~^ image[4][19] + signed_kernel[1][2] ~^ image[4][20] + signed_kernel[1][3] ~^ image[4][21] + signed_kernel[1][4] ~^ image[4][22] + signed_kernel[2][0] ~^ image[5][18] + signed_kernel[2][1] ~^ image[5][19] + signed_kernel[2][2] ~^ image[5][20] + signed_kernel[2][3] ~^ image[5][21] + signed_kernel[2][4] ~^ image[5][22] + signed_kernel[3][0] ~^ image[6][18] + signed_kernel[3][1] ~^ image[6][19] + signed_kernel[3][2] ~^ image[6][20] + signed_kernel[3][3] ~^ image[6][21] + signed_kernel[3][4] ~^ image[6][22] + signed_kernel[4][0] ~^ image[7][18] + signed_kernel[4][1] ~^ image[7][19] + signed_kernel[4][2] ~^ image[7][20] + signed_kernel[4][3] ~^ image[7][21] + signed_kernel[4][4] ~^ image[7][22];
assign xor_sum[3][19] = signed_kernel[0][0] ~^ image[3][19] + signed_kernel[0][1] ~^ image[3][20] + signed_kernel[0][2] ~^ image[3][21] + signed_kernel[0][3] ~^ image[3][22] + signed_kernel[0][4] ~^ image[3][23] + signed_kernel[1][0] ~^ image[4][19] + signed_kernel[1][1] ~^ image[4][20] + signed_kernel[1][2] ~^ image[4][21] + signed_kernel[1][3] ~^ image[4][22] + signed_kernel[1][4] ~^ image[4][23] + signed_kernel[2][0] ~^ image[5][19] + signed_kernel[2][1] ~^ image[5][20] + signed_kernel[2][2] ~^ image[5][21] + signed_kernel[2][3] ~^ image[5][22] + signed_kernel[2][4] ~^ image[5][23] + signed_kernel[3][0] ~^ image[6][19] + signed_kernel[3][1] ~^ image[6][20] + signed_kernel[3][2] ~^ image[6][21] + signed_kernel[3][3] ~^ image[6][22] + signed_kernel[3][4] ~^ image[6][23] + signed_kernel[4][0] ~^ image[7][19] + signed_kernel[4][1] ~^ image[7][20] + signed_kernel[4][2] ~^ image[7][21] + signed_kernel[4][3] ~^ image[7][22] + signed_kernel[4][4] ~^ image[7][23];
assign xor_sum[3][20] = signed_kernel[0][0] ~^ image[3][20] + signed_kernel[0][1] ~^ image[3][21] + signed_kernel[0][2] ~^ image[3][22] + signed_kernel[0][3] ~^ image[3][23] + signed_kernel[0][4] ~^ image[3][24] + signed_kernel[1][0] ~^ image[4][20] + signed_kernel[1][1] ~^ image[4][21] + signed_kernel[1][2] ~^ image[4][22] + signed_kernel[1][3] ~^ image[4][23] + signed_kernel[1][4] ~^ image[4][24] + signed_kernel[2][0] ~^ image[5][20] + signed_kernel[2][1] ~^ image[5][21] + signed_kernel[2][2] ~^ image[5][22] + signed_kernel[2][3] ~^ image[5][23] + signed_kernel[2][4] ~^ image[5][24] + signed_kernel[3][0] ~^ image[6][20] + signed_kernel[3][1] ~^ image[6][21] + signed_kernel[3][2] ~^ image[6][22] + signed_kernel[3][3] ~^ image[6][23] + signed_kernel[3][4] ~^ image[6][24] + signed_kernel[4][0] ~^ image[7][20] + signed_kernel[4][1] ~^ image[7][21] + signed_kernel[4][2] ~^ image[7][22] + signed_kernel[4][3] ~^ image[7][23] + signed_kernel[4][4] ~^ image[7][24];
assign xor_sum[3][21] = signed_kernel[0][0] ~^ image[3][21] + signed_kernel[0][1] ~^ image[3][22] + signed_kernel[0][2] ~^ image[3][23] + signed_kernel[0][3] ~^ image[3][24] + signed_kernel[0][4] ~^ image[3][25] + signed_kernel[1][0] ~^ image[4][21] + signed_kernel[1][1] ~^ image[4][22] + signed_kernel[1][2] ~^ image[4][23] + signed_kernel[1][3] ~^ image[4][24] + signed_kernel[1][4] ~^ image[4][25] + signed_kernel[2][0] ~^ image[5][21] + signed_kernel[2][1] ~^ image[5][22] + signed_kernel[2][2] ~^ image[5][23] + signed_kernel[2][3] ~^ image[5][24] + signed_kernel[2][4] ~^ image[5][25] + signed_kernel[3][0] ~^ image[6][21] + signed_kernel[3][1] ~^ image[6][22] + signed_kernel[3][2] ~^ image[6][23] + signed_kernel[3][3] ~^ image[6][24] + signed_kernel[3][4] ~^ image[6][25] + signed_kernel[4][0] ~^ image[7][21] + signed_kernel[4][1] ~^ image[7][22] + signed_kernel[4][2] ~^ image[7][23] + signed_kernel[4][3] ~^ image[7][24] + signed_kernel[4][4] ~^ image[7][25];
assign xor_sum[3][22] = signed_kernel[0][0] ~^ image[3][22] + signed_kernel[0][1] ~^ image[3][23] + signed_kernel[0][2] ~^ image[3][24] + signed_kernel[0][3] ~^ image[3][25] + signed_kernel[0][4] ~^ image[3][26] + signed_kernel[1][0] ~^ image[4][22] + signed_kernel[1][1] ~^ image[4][23] + signed_kernel[1][2] ~^ image[4][24] + signed_kernel[1][3] ~^ image[4][25] + signed_kernel[1][4] ~^ image[4][26] + signed_kernel[2][0] ~^ image[5][22] + signed_kernel[2][1] ~^ image[5][23] + signed_kernel[2][2] ~^ image[5][24] + signed_kernel[2][3] ~^ image[5][25] + signed_kernel[2][4] ~^ image[5][26] + signed_kernel[3][0] ~^ image[6][22] + signed_kernel[3][1] ~^ image[6][23] + signed_kernel[3][2] ~^ image[6][24] + signed_kernel[3][3] ~^ image[6][25] + signed_kernel[3][4] ~^ image[6][26] + signed_kernel[4][0] ~^ image[7][22] + signed_kernel[4][1] ~^ image[7][23] + signed_kernel[4][2] ~^ image[7][24] + signed_kernel[4][3] ~^ image[7][25] + signed_kernel[4][4] ~^ image[7][26];
assign xor_sum[3][23] = signed_kernel[0][0] ~^ image[3][23] + signed_kernel[0][1] ~^ image[3][24] + signed_kernel[0][2] ~^ image[3][25] + signed_kernel[0][3] ~^ image[3][26] + signed_kernel[0][4] ~^ image[3][27] + signed_kernel[1][0] ~^ image[4][23] + signed_kernel[1][1] ~^ image[4][24] + signed_kernel[1][2] ~^ image[4][25] + signed_kernel[1][3] ~^ image[4][26] + signed_kernel[1][4] ~^ image[4][27] + signed_kernel[2][0] ~^ image[5][23] + signed_kernel[2][1] ~^ image[5][24] + signed_kernel[2][2] ~^ image[5][25] + signed_kernel[2][3] ~^ image[5][26] + signed_kernel[2][4] ~^ image[5][27] + signed_kernel[3][0] ~^ image[6][23] + signed_kernel[3][1] ~^ image[6][24] + signed_kernel[3][2] ~^ image[6][25] + signed_kernel[3][3] ~^ image[6][26] + signed_kernel[3][4] ~^ image[6][27] + signed_kernel[4][0] ~^ image[7][23] + signed_kernel[4][1] ~^ image[7][24] + signed_kernel[4][2] ~^ image[7][25] + signed_kernel[4][3] ~^ image[7][26] + signed_kernel[4][4] ~^ image[7][27];
assign xor_sum[4][0] = signed_kernel[0][0] ~^ image[4][0] + signed_kernel[0][1] ~^ image[4][1] + signed_kernel[0][2] ~^ image[4][2] + signed_kernel[0][3] ~^ image[4][3] + signed_kernel[0][4] ~^ image[4][4] + signed_kernel[1][0] ~^ image[5][0] + signed_kernel[1][1] ~^ image[5][1] + signed_kernel[1][2] ~^ image[5][2] + signed_kernel[1][3] ~^ image[5][3] + signed_kernel[1][4] ~^ image[5][4] + signed_kernel[2][0] ~^ image[6][0] + signed_kernel[2][1] ~^ image[6][1] + signed_kernel[2][2] ~^ image[6][2] + signed_kernel[2][3] ~^ image[6][3] + signed_kernel[2][4] ~^ image[6][4] + signed_kernel[3][0] ~^ image[7][0] + signed_kernel[3][1] ~^ image[7][1] + signed_kernel[3][2] ~^ image[7][2] + signed_kernel[3][3] ~^ image[7][3] + signed_kernel[3][4] ~^ image[7][4] + signed_kernel[4][0] ~^ image[8][0] + signed_kernel[4][1] ~^ image[8][1] + signed_kernel[4][2] ~^ image[8][2] + signed_kernel[4][3] ~^ image[8][3] + signed_kernel[4][4] ~^ image[8][4];
assign xor_sum[4][1] = signed_kernel[0][0] ~^ image[4][1] + signed_kernel[0][1] ~^ image[4][2] + signed_kernel[0][2] ~^ image[4][3] + signed_kernel[0][3] ~^ image[4][4] + signed_kernel[0][4] ~^ image[4][5] + signed_kernel[1][0] ~^ image[5][1] + signed_kernel[1][1] ~^ image[5][2] + signed_kernel[1][2] ~^ image[5][3] + signed_kernel[1][3] ~^ image[5][4] + signed_kernel[1][4] ~^ image[5][5] + signed_kernel[2][0] ~^ image[6][1] + signed_kernel[2][1] ~^ image[6][2] + signed_kernel[2][2] ~^ image[6][3] + signed_kernel[2][3] ~^ image[6][4] + signed_kernel[2][4] ~^ image[6][5] + signed_kernel[3][0] ~^ image[7][1] + signed_kernel[3][1] ~^ image[7][2] + signed_kernel[3][2] ~^ image[7][3] + signed_kernel[3][3] ~^ image[7][4] + signed_kernel[3][4] ~^ image[7][5] + signed_kernel[4][0] ~^ image[8][1] + signed_kernel[4][1] ~^ image[8][2] + signed_kernel[4][2] ~^ image[8][3] + signed_kernel[4][3] ~^ image[8][4] + signed_kernel[4][4] ~^ image[8][5];
assign xor_sum[4][2] = signed_kernel[0][0] ~^ image[4][2] + signed_kernel[0][1] ~^ image[4][3] + signed_kernel[0][2] ~^ image[4][4] + signed_kernel[0][3] ~^ image[4][5] + signed_kernel[0][4] ~^ image[4][6] + signed_kernel[1][0] ~^ image[5][2] + signed_kernel[1][1] ~^ image[5][3] + signed_kernel[1][2] ~^ image[5][4] + signed_kernel[1][3] ~^ image[5][5] + signed_kernel[1][4] ~^ image[5][6] + signed_kernel[2][0] ~^ image[6][2] + signed_kernel[2][1] ~^ image[6][3] + signed_kernel[2][2] ~^ image[6][4] + signed_kernel[2][3] ~^ image[6][5] + signed_kernel[2][4] ~^ image[6][6] + signed_kernel[3][0] ~^ image[7][2] + signed_kernel[3][1] ~^ image[7][3] + signed_kernel[3][2] ~^ image[7][4] + signed_kernel[3][3] ~^ image[7][5] + signed_kernel[3][4] ~^ image[7][6] + signed_kernel[4][0] ~^ image[8][2] + signed_kernel[4][1] ~^ image[8][3] + signed_kernel[4][2] ~^ image[8][4] + signed_kernel[4][3] ~^ image[8][5] + signed_kernel[4][4] ~^ image[8][6];
assign xor_sum[4][3] = signed_kernel[0][0] ~^ image[4][3] + signed_kernel[0][1] ~^ image[4][4] + signed_kernel[0][2] ~^ image[4][5] + signed_kernel[0][3] ~^ image[4][6] + signed_kernel[0][4] ~^ image[4][7] + signed_kernel[1][0] ~^ image[5][3] + signed_kernel[1][1] ~^ image[5][4] + signed_kernel[1][2] ~^ image[5][5] + signed_kernel[1][3] ~^ image[5][6] + signed_kernel[1][4] ~^ image[5][7] + signed_kernel[2][0] ~^ image[6][3] + signed_kernel[2][1] ~^ image[6][4] + signed_kernel[2][2] ~^ image[6][5] + signed_kernel[2][3] ~^ image[6][6] + signed_kernel[2][4] ~^ image[6][7] + signed_kernel[3][0] ~^ image[7][3] + signed_kernel[3][1] ~^ image[7][4] + signed_kernel[3][2] ~^ image[7][5] + signed_kernel[3][3] ~^ image[7][6] + signed_kernel[3][4] ~^ image[7][7] + signed_kernel[4][0] ~^ image[8][3] + signed_kernel[4][1] ~^ image[8][4] + signed_kernel[4][2] ~^ image[8][5] + signed_kernel[4][3] ~^ image[8][6] + signed_kernel[4][4] ~^ image[8][7];
assign xor_sum[4][4] = signed_kernel[0][0] ~^ image[4][4] + signed_kernel[0][1] ~^ image[4][5] + signed_kernel[0][2] ~^ image[4][6] + signed_kernel[0][3] ~^ image[4][7] + signed_kernel[0][4] ~^ image[4][8] + signed_kernel[1][0] ~^ image[5][4] + signed_kernel[1][1] ~^ image[5][5] + signed_kernel[1][2] ~^ image[5][6] + signed_kernel[1][3] ~^ image[5][7] + signed_kernel[1][4] ~^ image[5][8] + signed_kernel[2][0] ~^ image[6][4] + signed_kernel[2][1] ~^ image[6][5] + signed_kernel[2][2] ~^ image[6][6] + signed_kernel[2][3] ~^ image[6][7] + signed_kernel[2][4] ~^ image[6][8] + signed_kernel[3][0] ~^ image[7][4] + signed_kernel[3][1] ~^ image[7][5] + signed_kernel[3][2] ~^ image[7][6] + signed_kernel[3][3] ~^ image[7][7] + signed_kernel[3][4] ~^ image[7][8] + signed_kernel[4][0] ~^ image[8][4] + signed_kernel[4][1] ~^ image[8][5] + signed_kernel[4][2] ~^ image[8][6] + signed_kernel[4][3] ~^ image[8][7] + signed_kernel[4][4] ~^ image[8][8];
assign xor_sum[4][5] = signed_kernel[0][0] ~^ image[4][5] + signed_kernel[0][1] ~^ image[4][6] + signed_kernel[0][2] ~^ image[4][7] + signed_kernel[0][3] ~^ image[4][8] + signed_kernel[0][4] ~^ image[4][9] + signed_kernel[1][0] ~^ image[5][5] + signed_kernel[1][1] ~^ image[5][6] + signed_kernel[1][2] ~^ image[5][7] + signed_kernel[1][3] ~^ image[5][8] + signed_kernel[1][4] ~^ image[5][9] + signed_kernel[2][0] ~^ image[6][5] + signed_kernel[2][1] ~^ image[6][6] + signed_kernel[2][2] ~^ image[6][7] + signed_kernel[2][3] ~^ image[6][8] + signed_kernel[2][4] ~^ image[6][9] + signed_kernel[3][0] ~^ image[7][5] + signed_kernel[3][1] ~^ image[7][6] + signed_kernel[3][2] ~^ image[7][7] + signed_kernel[3][3] ~^ image[7][8] + signed_kernel[3][4] ~^ image[7][9] + signed_kernel[4][0] ~^ image[8][5] + signed_kernel[4][1] ~^ image[8][6] + signed_kernel[4][2] ~^ image[8][7] + signed_kernel[4][3] ~^ image[8][8] + signed_kernel[4][4] ~^ image[8][9];
assign xor_sum[4][6] = signed_kernel[0][0] ~^ image[4][6] + signed_kernel[0][1] ~^ image[4][7] + signed_kernel[0][2] ~^ image[4][8] + signed_kernel[0][3] ~^ image[4][9] + signed_kernel[0][4] ~^ image[4][10] + signed_kernel[1][0] ~^ image[5][6] + signed_kernel[1][1] ~^ image[5][7] + signed_kernel[1][2] ~^ image[5][8] + signed_kernel[1][3] ~^ image[5][9] + signed_kernel[1][4] ~^ image[5][10] + signed_kernel[2][0] ~^ image[6][6] + signed_kernel[2][1] ~^ image[6][7] + signed_kernel[2][2] ~^ image[6][8] + signed_kernel[2][3] ~^ image[6][9] + signed_kernel[2][4] ~^ image[6][10] + signed_kernel[3][0] ~^ image[7][6] + signed_kernel[3][1] ~^ image[7][7] + signed_kernel[3][2] ~^ image[7][8] + signed_kernel[3][3] ~^ image[7][9] + signed_kernel[3][4] ~^ image[7][10] + signed_kernel[4][0] ~^ image[8][6] + signed_kernel[4][1] ~^ image[8][7] + signed_kernel[4][2] ~^ image[8][8] + signed_kernel[4][3] ~^ image[8][9] + signed_kernel[4][4] ~^ image[8][10];
assign xor_sum[4][7] = signed_kernel[0][0] ~^ image[4][7] + signed_kernel[0][1] ~^ image[4][8] + signed_kernel[0][2] ~^ image[4][9] + signed_kernel[0][3] ~^ image[4][10] + signed_kernel[0][4] ~^ image[4][11] + signed_kernel[1][0] ~^ image[5][7] + signed_kernel[1][1] ~^ image[5][8] + signed_kernel[1][2] ~^ image[5][9] + signed_kernel[1][3] ~^ image[5][10] + signed_kernel[1][4] ~^ image[5][11] + signed_kernel[2][0] ~^ image[6][7] + signed_kernel[2][1] ~^ image[6][8] + signed_kernel[2][2] ~^ image[6][9] + signed_kernel[2][3] ~^ image[6][10] + signed_kernel[2][4] ~^ image[6][11] + signed_kernel[3][0] ~^ image[7][7] + signed_kernel[3][1] ~^ image[7][8] + signed_kernel[3][2] ~^ image[7][9] + signed_kernel[3][3] ~^ image[7][10] + signed_kernel[3][4] ~^ image[7][11] + signed_kernel[4][0] ~^ image[8][7] + signed_kernel[4][1] ~^ image[8][8] + signed_kernel[4][2] ~^ image[8][9] + signed_kernel[4][3] ~^ image[8][10] + signed_kernel[4][4] ~^ image[8][11];
assign xor_sum[4][8] = signed_kernel[0][0] ~^ image[4][8] + signed_kernel[0][1] ~^ image[4][9] + signed_kernel[0][2] ~^ image[4][10] + signed_kernel[0][3] ~^ image[4][11] + signed_kernel[0][4] ~^ image[4][12] + signed_kernel[1][0] ~^ image[5][8] + signed_kernel[1][1] ~^ image[5][9] + signed_kernel[1][2] ~^ image[5][10] + signed_kernel[1][3] ~^ image[5][11] + signed_kernel[1][4] ~^ image[5][12] + signed_kernel[2][0] ~^ image[6][8] + signed_kernel[2][1] ~^ image[6][9] + signed_kernel[2][2] ~^ image[6][10] + signed_kernel[2][3] ~^ image[6][11] + signed_kernel[2][4] ~^ image[6][12] + signed_kernel[3][0] ~^ image[7][8] + signed_kernel[3][1] ~^ image[7][9] + signed_kernel[3][2] ~^ image[7][10] + signed_kernel[3][3] ~^ image[7][11] + signed_kernel[3][4] ~^ image[7][12] + signed_kernel[4][0] ~^ image[8][8] + signed_kernel[4][1] ~^ image[8][9] + signed_kernel[4][2] ~^ image[8][10] + signed_kernel[4][3] ~^ image[8][11] + signed_kernel[4][4] ~^ image[8][12];
assign xor_sum[4][9] = signed_kernel[0][0] ~^ image[4][9] + signed_kernel[0][1] ~^ image[4][10] + signed_kernel[0][2] ~^ image[4][11] + signed_kernel[0][3] ~^ image[4][12] + signed_kernel[0][4] ~^ image[4][13] + signed_kernel[1][0] ~^ image[5][9] + signed_kernel[1][1] ~^ image[5][10] + signed_kernel[1][2] ~^ image[5][11] + signed_kernel[1][3] ~^ image[5][12] + signed_kernel[1][4] ~^ image[5][13] + signed_kernel[2][0] ~^ image[6][9] + signed_kernel[2][1] ~^ image[6][10] + signed_kernel[2][2] ~^ image[6][11] + signed_kernel[2][3] ~^ image[6][12] + signed_kernel[2][4] ~^ image[6][13] + signed_kernel[3][0] ~^ image[7][9] + signed_kernel[3][1] ~^ image[7][10] + signed_kernel[3][2] ~^ image[7][11] + signed_kernel[3][3] ~^ image[7][12] + signed_kernel[3][4] ~^ image[7][13] + signed_kernel[4][0] ~^ image[8][9] + signed_kernel[4][1] ~^ image[8][10] + signed_kernel[4][2] ~^ image[8][11] + signed_kernel[4][3] ~^ image[8][12] + signed_kernel[4][4] ~^ image[8][13];
assign xor_sum[4][10] = signed_kernel[0][0] ~^ image[4][10] + signed_kernel[0][1] ~^ image[4][11] + signed_kernel[0][2] ~^ image[4][12] + signed_kernel[0][3] ~^ image[4][13] + signed_kernel[0][4] ~^ image[4][14] + signed_kernel[1][0] ~^ image[5][10] + signed_kernel[1][1] ~^ image[5][11] + signed_kernel[1][2] ~^ image[5][12] + signed_kernel[1][3] ~^ image[5][13] + signed_kernel[1][4] ~^ image[5][14] + signed_kernel[2][0] ~^ image[6][10] + signed_kernel[2][1] ~^ image[6][11] + signed_kernel[2][2] ~^ image[6][12] + signed_kernel[2][3] ~^ image[6][13] + signed_kernel[2][4] ~^ image[6][14] + signed_kernel[3][0] ~^ image[7][10] + signed_kernel[3][1] ~^ image[7][11] + signed_kernel[3][2] ~^ image[7][12] + signed_kernel[3][3] ~^ image[7][13] + signed_kernel[3][4] ~^ image[7][14] + signed_kernel[4][0] ~^ image[8][10] + signed_kernel[4][1] ~^ image[8][11] + signed_kernel[4][2] ~^ image[8][12] + signed_kernel[4][3] ~^ image[8][13] + signed_kernel[4][4] ~^ image[8][14];
assign xor_sum[4][11] = signed_kernel[0][0] ~^ image[4][11] + signed_kernel[0][1] ~^ image[4][12] + signed_kernel[0][2] ~^ image[4][13] + signed_kernel[0][3] ~^ image[4][14] + signed_kernel[0][4] ~^ image[4][15] + signed_kernel[1][0] ~^ image[5][11] + signed_kernel[1][1] ~^ image[5][12] + signed_kernel[1][2] ~^ image[5][13] + signed_kernel[1][3] ~^ image[5][14] + signed_kernel[1][4] ~^ image[5][15] + signed_kernel[2][0] ~^ image[6][11] + signed_kernel[2][1] ~^ image[6][12] + signed_kernel[2][2] ~^ image[6][13] + signed_kernel[2][3] ~^ image[6][14] + signed_kernel[2][4] ~^ image[6][15] + signed_kernel[3][0] ~^ image[7][11] + signed_kernel[3][1] ~^ image[7][12] + signed_kernel[3][2] ~^ image[7][13] + signed_kernel[3][3] ~^ image[7][14] + signed_kernel[3][4] ~^ image[7][15] + signed_kernel[4][0] ~^ image[8][11] + signed_kernel[4][1] ~^ image[8][12] + signed_kernel[4][2] ~^ image[8][13] + signed_kernel[4][3] ~^ image[8][14] + signed_kernel[4][4] ~^ image[8][15];
assign xor_sum[4][12] = signed_kernel[0][0] ~^ image[4][12] + signed_kernel[0][1] ~^ image[4][13] + signed_kernel[0][2] ~^ image[4][14] + signed_kernel[0][3] ~^ image[4][15] + signed_kernel[0][4] ~^ image[4][16] + signed_kernel[1][0] ~^ image[5][12] + signed_kernel[1][1] ~^ image[5][13] + signed_kernel[1][2] ~^ image[5][14] + signed_kernel[1][3] ~^ image[5][15] + signed_kernel[1][4] ~^ image[5][16] + signed_kernel[2][0] ~^ image[6][12] + signed_kernel[2][1] ~^ image[6][13] + signed_kernel[2][2] ~^ image[6][14] + signed_kernel[2][3] ~^ image[6][15] + signed_kernel[2][4] ~^ image[6][16] + signed_kernel[3][0] ~^ image[7][12] + signed_kernel[3][1] ~^ image[7][13] + signed_kernel[3][2] ~^ image[7][14] + signed_kernel[3][3] ~^ image[7][15] + signed_kernel[3][4] ~^ image[7][16] + signed_kernel[4][0] ~^ image[8][12] + signed_kernel[4][1] ~^ image[8][13] + signed_kernel[4][2] ~^ image[8][14] + signed_kernel[4][3] ~^ image[8][15] + signed_kernel[4][4] ~^ image[8][16];
assign xor_sum[4][13] = signed_kernel[0][0] ~^ image[4][13] + signed_kernel[0][1] ~^ image[4][14] + signed_kernel[0][2] ~^ image[4][15] + signed_kernel[0][3] ~^ image[4][16] + signed_kernel[0][4] ~^ image[4][17] + signed_kernel[1][0] ~^ image[5][13] + signed_kernel[1][1] ~^ image[5][14] + signed_kernel[1][2] ~^ image[5][15] + signed_kernel[1][3] ~^ image[5][16] + signed_kernel[1][4] ~^ image[5][17] + signed_kernel[2][0] ~^ image[6][13] + signed_kernel[2][1] ~^ image[6][14] + signed_kernel[2][2] ~^ image[6][15] + signed_kernel[2][3] ~^ image[6][16] + signed_kernel[2][4] ~^ image[6][17] + signed_kernel[3][0] ~^ image[7][13] + signed_kernel[3][1] ~^ image[7][14] + signed_kernel[3][2] ~^ image[7][15] + signed_kernel[3][3] ~^ image[7][16] + signed_kernel[3][4] ~^ image[7][17] + signed_kernel[4][0] ~^ image[8][13] + signed_kernel[4][1] ~^ image[8][14] + signed_kernel[4][2] ~^ image[8][15] + signed_kernel[4][3] ~^ image[8][16] + signed_kernel[4][4] ~^ image[8][17];
assign xor_sum[4][14] = signed_kernel[0][0] ~^ image[4][14] + signed_kernel[0][1] ~^ image[4][15] + signed_kernel[0][2] ~^ image[4][16] + signed_kernel[0][3] ~^ image[4][17] + signed_kernel[0][4] ~^ image[4][18] + signed_kernel[1][0] ~^ image[5][14] + signed_kernel[1][1] ~^ image[5][15] + signed_kernel[1][2] ~^ image[5][16] + signed_kernel[1][3] ~^ image[5][17] + signed_kernel[1][4] ~^ image[5][18] + signed_kernel[2][0] ~^ image[6][14] + signed_kernel[2][1] ~^ image[6][15] + signed_kernel[2][2] ~^ image[6][16] + signed_kernel[2][3] ~^ image[6][17] + signed_kernel[2][4] ~^ image[6][18] + signed_kernel[3][0] ~^ image[7][14] + signed_kernel[3][1] ~^ image[7][15] + signed_kernel[3][2] ~^ image[7][16] + signed_kernel[3][3] ~^ image[7][17] + signed_kernel[3][4] ~^ image[7][18] + signed_kernel[4][0] ~^ image[8][14] + signed_kernel[4][1] ~^ image[8][15] + signed_kernel[4][2] ~^ image[8][16] + signed_kernel[4][3] ~^ image[8][17] + signed_kernel[4][4] ~^ image[8][18];
assign xor_sum[4][15] = signed_kernel[0][0] ~^ image[4][15] + signed_kernel[0][1] ~^ image[4][16] + signed_kernel[0][2] ~^ image[4][17] + signed_kernel[0][3] ~^ image[4][18] + signed_kernel[0][4] ~^ image[4][19] + signed_kernel[1][0] ~^ image[5][15] + signed_kernel[1][1] ~^ image[5][16] + signed_kernel[1][2] ~^ image[5][17] + signed_kernel[1][3] ~^ image[5][18] + signed_kernel[1][4] ~^ image[5][19] + signed_kernel[2][0] ~^ image[6][15] + signed_kernel[2][1] ~^ image[6][16] + signed_kernel[2][2] ~^ image[6][17] + signed_kernel[2][3] ~^ image[6][18] + signed_kernel[2][4] ~^ image[6][19] + signed_kernel[3][0] ~^ image[7][15] + signed_kernel[3][1] ~^ image[7][16] + signed_kernel[3][2] ~^ image[7][17] + signed_kernel[3][3] ~^ image[7][18] + signed_kernel[3][4] ~^ image[7][19] + signed_kernel[4][0] ~^ image[8][15] + signed_kernel[4][1] ~^ image[8][16] + signed_kernel[4][2] ~^ image[8][17] + signed_kernel[4][3] ~^ image[8][18] + signed_kernel[4][4] ~^ image[8][19];
assign xor_sum[4][16] = signed_kernel[0][0] ~^ image[4][16] + signed_kernel[0][1] ~^ image[4][17] + signed_kernel[0][2] ~^ image[4][18] + signed_kernel[0][3] ~^ image[4][19] + signed_kernel[0][4] ~^ image[4][20] + signed_kernel[1][0] ~^ image[5][16] + signed_kernel[1][1] ~^ image[5][17] + signed_kernel[1][2] ~^ image[5][18] + signed_kernel[1][3] ~^ image[5][19] + signed_kernel[1][4] ~^ image[5][20] + signed_kernel[2][0] ~^ image[6][16] + signed_kernel[2][1] ~^ image[6][17] + signed_kernel[2][2] ~^ image[6][18] + signed_kernel[2][3] ~^ image[6][19] + signed_kernel[2][4] ~^ image[6][20] + signed_kernel[3][0] ~^ image[7][16] + signed_kernel[3][1] ~^ image[7][17] + signed_kernel[3][2] ~^ image[7][18] + signed_kernel[3][3] ~^ image[7][19] + signed_kernel[3][4] ~^ image[7][20] + signed_kernel[4][0] ~^ image[8][16] + signed_kernel[4][1] ~^ image[8][17] + signed_kernel[4][2] ~^ image[8][18] + signed_kernel[4][3] ~^ image[8][19] + signed_kernel[4][4] ~^ image[8][20];
assign xor_sum[4][17] = signed_kernel[0][0] ~^ image[4][17] + signed_kernel[0][1] ~^ image[4][18] + signed_kernel[0][2] ~^ image[4][19] + signed_kernel[0][3] ~^ image[4][20] + signed_kernel[0][4] ~^ image[4][21] + signed_kernel[1][0] ~^ image[5][17] + signed_kernel[1][1] ~^ image[5][18] + signed_kernel[1][2] ~^ image[5][19] + signed_kernel[1][3] ~^ image[5][20] + signed_kernel[1][4] ~^ image[5][21] + signed_kernel[2][0] ~^ image[6][17] + signed_kernel[2][1] ~^ image[6][18] + signed_kernel[2][2] ~^ image[6][19] + signed_kernel[2][3] ~^ image[6][20] + signed_kernel[2][4] ~^ image[6][21] + signed_kernel[3][0] ~^ image[7][17] + signed_kernel[3][1] ~^ image[7][18] + signed_kernel[3][2] ~^ image[7][19] + signed_kernel[3][3] ~^ image[7][20] + signed_kernel[3][4] ~^ image[7][21] + signed_kernel[4][0] ~^ image[8][17] + signed_kernel[4][1] ~^ image[8][18] + signed_kernel[4][2] ~^ image[8][19] + signed_kernel[4][3] ~^ image[8][20] + signed_kernel[4][4] ~^ image[8][21];
assign xor_sum[4][18] = signed_kernel[0][0] ~^ image[4][18] + signed_kernel[0][1] ~^ image[4][19] + signed_kernel[0][2] ~^ image[4][20] + signed_kernel[0][3] ~^ image[4][21] + signed_kernel[0][4] ~^ image[4][22] + signed_kernel[1][0] ~^ image[5][18] + signed_kernel[1][1] ~^ image[5][19] + signed_kernel[1][2] ~^ image[5][20] + signed_kernel[1][3] ~^ image[5][21] + signed_kernel[1][4] ~^ image[5][22] + signed_kernel[2][0] ~^ image[6][18] + signed_kernel[2][1] ~^ image[6][19] + signed_kernel[2][2] ~^ image[6][20] + signed_kernel[2][3] ~^ image[6][21] + signed_kernel[2][4] ~^ image[6][22] + signed_kernel[3][0] ~^ image[7][18] + signed_kernel[3][1] ~^ image[7][19] + signed_kernel[3][2] ~^ image[7][20] + signed_kernel[3][3] ~^ image[7][21] + signed_kernel[3][4] ~^ image[7][22] + signed_kernel[4][0] ~^ image[8][18] + signed_kernel[4][1] ~^ image[8][19] + signed_kernel[4][2] ~^ image[8][20] + signed_kernel[4][3] ~^ image[8][21] + signed_kernel[4][4] ~^ image[8][22];
assign xor_sum[4][19] = signed_kernel[0][0] ~^ image[4][19] + signed_kernel[0][1] ~^ image[4][20] + signed_kernel[0][2] ~^ image[4][21] + signed_kernel[0][3] ~^ image[4][22] + signed_kernel[0][4] ~^ image[4][23] + signed_kernel[1][0] ~^ image[5][19] + signed_kernel[1][1] ~^ image[5][20] + signed_kernel[1][2] ~^ image[5][21] + signed_kernel[1][3] ~^ image[5][22] + signed_kernel[1][4] ~^ image[5][23] + signed_kernel[2][0] ~^ image[6][19] + signed_kernel[2][1] ~^ image[6][20] + signed_kernel[2][2] ~^ image[6][21] + signed_kernel[2][3] ~^ image[6][22] + signed_kernel[2][4] ~^ image[6][23] + signed_kernel[3][0] ~^ image[7][19] + signed_kernel[3][1] ~^ image[7][20] + signed_kernel[3][2] ~^ image[7][21] + signed_kernel[3][3] ~^ image[7][22] + signed_kernel[3][4] ~^ image[7][23] + signed_kernel[4][0] ~^ image[8][19] + signed_kernel[4][1] ~^ image[8][20] + signed_kernel[4][2] ~^ image[8][21] + signed_kernel[4][3] ~^ image[8][22] + signed_kernel[4][4] ~^ image[8][23];
assign xor_sum[4][20] = signed_kernel[0][0] ~^ image[4][20] + signed_kernel[0][1] ~^ image[4][21] + signed_kernel[0][2] ~^ image[4][22] + signed_kernel[0][3] ~^ image[4][23] + signed_kernel[0][4] ~^ image[4][24] + signed_kernel[1][0] ~^ image[5][20] + signed_kernel[1][1] ~^ image[5][21] + signed_kernel[1][2] ~^ image[5][22] + signed_kernel[1][3] ~^ image[5][23] + signed_kernel[1][4] ~^ image[5][24] + signed_kernel[2][0] ~^ image[6][20] + signed_kernel[2][1] ~^ image[6][21] + signed_kernel[2][2] ~^ image[6][22] + signed_kernel[2][3] ~^ image[6][23] + signed_kernel[2][4] ~^ image[6][24] + signed_kernel[3][0] ~^ image[7][20] + signed_kernel[3][1] ~^ image[7][21] + signed_kernel[3][2] ~^ image[7][22] + signed_kernel[3][3] ~^ image[7][23] + signed_kernel[3][4] ~^ image[7][24] + signed_kernel[4][0] ~^ image[8][20] + signed_kernel[4][1] ~^ image[8][21] + signed_kernel[4][2] ~^ image[8][22] + signed_kernel[4][3] ~^ image[8][23] + signed_kernel[4][4] ~^ image[8][24];
assign xor_sum[4][21] = signed_kernel[0][0] ~^ image[4][21] + signed_kernel[0][1] ~^ image[4][22] + signed_kernel[0][2] ~^ image[4][23] + signed_kernel[0][3] ~^ image[4][24] + signed_kernel[0][4] ~^ image[4][25] + signed_kernel[1][0] ~^ image[5][21] + signed_kernel[1][1] ~^ image[5][22] + signed_kernel[1][2] ~^ image[5][23] + signed_kernel[1][3] ~^ image[5][24] + signed_kernel[1][4] ~^ image[5][25] + signed_kernel[2][0] ~^ image[6][21] + signed_kernel[2][1] ~^ image[6][22] + signed_kernel[2][2] ~^ image[6][23] + signed_kernel[2][3] ~^ image[6][24] + signed_kernel[2][4] ~^ image[6][25] + signed_kernel[3][0] ~^ image[7][21] + signed_kernel[3][1] ~^ image[7][22] + signed_kernel[3][2] ~^ image[7][23] + signed_kernel[3][3] ~^ image[7][24] + signed_kernel[3][4] ~^ image[7][25] + signed_kernel[4][0] ~^ image[8][21] + signed_kernel[4][1] ~^ image[8][22] + signed_kernel[4][2] ~^ image[8][23] + signed_kernel[4][3] ~^ image[8][24] + signed_kernel[4][4] ~^ image[8][25];
assign xor_sum[4][22] = signed_kernel[0][0] ~^ image[4][22] + signed_kernel[0][1] ~^ image[4][23] + signed_kernel[0][2] ~^ image[4][24] + signed_kernel[0][3] ~^ image[4][25] + signed_kernel[0][4] ~^ image[4][26] + signed_kernel[1][0] ~^ image[5][22] + signed_kernel[1][1] ~^ image[5][23] + signed_kernel[1][2] ~^ image[5][24] + signed_kernel[1][3] ~^ image[5][25] + signed_kernel[1][4] ~^ image[5][26] + signed_kernel[2][0] ~^ image[6][22] + signed_kernel[2][1] ~^ image[6][23] + signed_kernel[2][2] ~^ image[6][24] + signed_kernel[2][3] ~^ image[6][25] + signed_kernel[2][4] ~^ image[6][26] + signed_kernel[3][0] ~^ image[7][22] + signed_kernel[3][1] ~^ image[7][23] + signed_kernel[3][2] ~^ image[7][24] + signed_kernel[3][3] ~^ image[7][25] + signed_kernel[3][4] ~^ image[7][26] + signed_kernel[4][0] ~^ image[8][22] + signed_kernel[4][1] ~^ image[8][23] + signed_kernel[4][2] ~^ image[8][24] + signed_kernel[4][3] ~^ image[8][25] + signed_kernel[4][4] ~^ image[8][26];
assign xor_sum[4][23] = signed_kernel[0][0] ~^ image[4][23] + signed_kernel[0][1] ~^ image[4][24] + signed_kernel[0][2] ~^ image[4][25] + signed_kernel[0][3] ~^ image[4][26] + signed_kernel[0][4] ~^ image[4][27] + signed_kernel[1][0] ~^ image[5][23] + signed_kernel[1][1] ~^ image[5][24] + signed_kernel[1][2] ~^ image[5][25] + signed_kernel[1][3] ~^ image[5][26] + signed_kernel[1][4] ~^ image[5][27] + signed_kernel[2][0] ~^ image[6][23] + signed_kernel[2][1] ~^ image[6][24] + signed_kernel[2][2] ~^ image[6][25] + signed_kernel[2][3] ~^ image[6][26] + signed_kernel[2][4] ~^ image[6][27] + signed_kernel[3][0] ~^ image[7][23] + signed_kernel[3][1] ~^ image[7][24] + signed_kernel[3][2] ~^ image[7][25] + signed_kernel[3][3] ~^ image[7][26] + signed_kernel[3][4] ~^ image[7][27] + signed_kernel[4][0] ~^ image[8][23] + signed_kernel[4][1] ~^ image[8][24] + signed_kernel[4][2] ~^ image[8][25] + signed_kernel[4][3] ~^ image[8][26] + signed_kernel[4][4] ~^ image[8][27];
assign xor_sum[5][0] = signed_kernel[0][0] ~^ image[5][0] + signed_kernel[0][1] ~^ image[5][1] + signed_kernel[0][2] ~^ image[5][2] + signed_kernel[0][3] ~^ image[5][3] + signed_kernel[0][4] ~^ image[5][4] + signed_kernel[1][0] ~^ image[6][0] + signed_kernel[1][1] ~^ image[6][1] + signed_kernel[1][2] ~^ image[6][2] + signed_kernel[1][3] ~^ image[6][3] + signed_kernel[1][4] ~^ image[6][4] + signed_kernel[2][0] ~^ image[7][0] + signed_kernel[2][1] ~^ image[7][1] + signed_kernel[2][2] ~^ image[7][2] + signed_kernel[2][3] ~^ image[7][3] + signed_kernel[2][4] ~^ image[7][4] + signed_kernel[3][0] ~^ image[8][0] + signed_kernel[3][1] ~^ image[8][1] + signed_kernel[3][2] ~^ image[8][2] + signed_kernel[3][3] ~^ image[8][3] + signed_kernel[3][4] ~^ image[8][4] + signed_kernel[4][0] ~^ image[9][0] + signed_kernel[4][1] ~^ image[9][1] + signed_kernel[4][2] ~^ image[9][2] + signed_kernel[4][3] ~^ image[9][3] + signed_kernel[4][4] ~^ image[9][4];
assign xor_sum[5][1] = signed_kernel[0][0] ~^ image[5][1] + signed_kernel[0][1] ~^ image[5][2] + signed_kernel[0][2] ~^ image[5][3] + signed_kernel[0][3] ~^ image[5][4] + signed_kernel[0][4] ~^ image[5][5] + signed_kernel[1][0] ~^ image[6][1] + signed_kernel[1][1] ~^ image[6][2] + signed_kernel[1][2] ~^ image[6][3] + signed_kernel[1][3] ~^ image[6][4] + signed_kernel[1][4] ~^ image[6][5] + signed_kernel[2][0] ~^ image[7][1] + signed_kernel[2][1] ~^ image[7][2] + signed_kernel[2][2] ~^ image[7][3] + signed_kernel[2][3] ~^ image[7][4] + signed_kernel[2][4] ~^ image[7][5] + signed_kernel[3][0] ~^ image[8][1] + signed_kernel[3][1] ~^ image[8][2] + signed_kernel[3][2] ~^ image[8][3] + signed_kernel[3][3] ~^ image[8][4] + signed_kernel[3][4] ~^ image[8][5] + signed_kernel[4][0] ~^ image[9][1] + signed_kernel[4][1] ~^ image[9][2] + signed_kernel[4][2] ~^ image[9][3] + signed_kernel[4][3] ~^ image[9][4] + signed_kernel[4][4] ~^ image[9][5];
assign xor_sum[5][2] = signed_kernel[0][0] ~^ image[5][2] + signed_kernel[0][1] ~^ image[5][3] + signed_kernel[0][2] ~^ image[5][4] + signed_kernel[0][3] ~^ image[5][5] + signed_kernel[0][4] ~^ image[5][6] + signed_kernel[1][0] ~^ image[6][2] + signed_kernel[1][1] ~^ image[6][3] + signed_kernel[1][2] ~^ image[6][4] + signed_kernel[1][3] ~^ image[6][5] + signed_kernel[1][4] ~^ image[6][6] + signed_kernel[2][0] ~^ image[7][2] + signed_kernel[2][1] ~^ image[7][3] + signed_kernel[2][2] ~^ image[7][4] + signed_kernel[2][3] ~^ image[7][5] + signed_kernel[2][4] ~^ image[7][6] + signed_kernel[3][0] ~^ image[8][2] + signed_kernel[3][1] ~^ image[8][3] + signed_kernel[3][2] ~^ image[8][4] + signed_kernel[3][3] ~^ image[8][5] + signed_kernel[3][4] ~^ image[8][6] + signed_kernel[4][0] ~^ image[9][2] + signed_kernel[4][1] ~^ image[9][3] + signed_kernel[4][2] ~^ image[9][4] + signed_kernel[4][3] ~^ image[9][5] + signed_kernel[4][4] ~^ image[9][6];
assign xor_sum[5][3] = signed_kernel[0][0] ~^ image[5][3] + signed_kernel[0][1] ~^ image[5][4] + signed_kernel[0][2] ~^ image[5][5] + signed_kernel[0][3] ~^ image[5][6] + signed_kernel[0][4] ~^ image[5][7] + signed_kernel[1][0] ~^ image[6][3] + signed_kernel[1][1] ~^ image[6][4] + signed_kernel[1][2] ~^ image[6][5] + signed_kernel[1][3] ~^ image[6][6] + signed_kernel[1][4] ~^ image[6][7] + signed_kernel[2][0] ~^ image[7][3] + signed_kernel[2][1] ~^ image[7][4] + signed_kernel[2][2] ~^ image[7][5] + signed_kernel[2][3] ~^ image[7][6] + signed_kernel[2][4] ~^ image[7][7] + signed_kernel[3][0] ~^ image[8][3] + signed_kernel[3][1] ~^ image[8][4] + signed_kernel[3][2] ~^ image[8][5] + signed_kernel[3][3] ~^ image[8][6] + signed_kernel[3][4] ~^ image[8][7] + signed_kernel[4][0] ~^ image[9][3] + signed_kernel[4][1] ~^ image[9][4] + signed_kernel[4][2] ~^ image[9][5] + signed_kernel[4][3] ~^ image[9][6] + signed_kernel[4][4] ~^ image[9][7];
assign xor_sum[5][4] = signed_kernel[0][0] ~^ image[5][4] + signed_kernel[0][1] ~^ image[5][5] + signed_kernel[0][2] ~^ image[5][6] + signed_kernel[0][3] ~^ image[5][7] + signed_kernel[0][4] ~^ image[5][8] + signed_kernel[1][0] ~^ image[6][4] + signed_kernel[1][1] ~^ image[6][5] + signed_kernel[1][2] ~^ image[6][6] + signed_kernel[1][3] ~^ image[6][7] + signed_kernel[1][4] ~^ image[6][8] + signed_kernel[2][0] ~^ image[7][4] + signed_kernel[2][1] ~^ image[7][5] + signed_kernel[2][2] ~^ image[7][6] + signed_kernel[2][3] ~^ image[7][7] + signed_kernel[2][4] ~^ image[7][8] + signed_kernel[3][0] ~^ image[8][4] + signed_kernel[3][1] ~^ image[8][5] + signed_kernel[3][2] ~^ image[8][6] + signed_kernel[3][3] ~^ image[8][7] + signed_kernel[3][4] ~^ image[8][8] + signed_kernel[4][0] ~^ image[9][4] + signed_kernel[4][1] ~^ image[9][5] + signed_kernel[4][2] ~^ image[9][6] + signed_kernel[4][3] ~^ image[9][7] + signed_kernel[4][4] ~^ image[9][8];
assign xor_sum[5][5] = signed_kernel[0][0] ~^ image[5][5] + signed_kernel[0][1] ~^ image[5][6] + signed_kernel[0][2] ~^ image[5][7] + signed_kernel[0][3] ~^ image[5][8] + signed_kernel[0][4] ~^ image[5][9] + signed_kernel[1][0] ~^ image[6][5] + signed_kernel[1][1] ~^ image[6][6] + signed_kernel[1][2] ~^ image[6][7] + signed_kernel[1][3] ~^ image[6][8] + signed_kernel[1][4] ~^ image[6][9] + signed_kernel[2][0] ~^ image[7][5] + signed_kernel[2][1] ~^ image[7][6] + signed_kernel[2][2] ~^ image[7][7] + signed_kernel[2][3] ~^ image[7][8] + signed_kernel[2][4] ~^ image[7][9] + signed_kernel[3][0] ~^ image[8][5] + signed_kernel[3][1] ~^ image[8][6] + signed_kernel[3][2] ~^ image[8][7] + signed_kernel[3][3] ~^ image[8][8] + signed_kernel[3][4] ~^ image[8][9] + signed_kernel[4][0] ~^ image[9][5] + signed_kernel[4][1] ~^ image[9][6] + signed_kernel[4][2] ~^ image[9][7] + signed_kernel[4][3] ~^ image[9][8] + signed_kernel[4][4] ~^ image[9][9];
assign xor_sum[5][6] = signed_kernel[0][0] ~^ image[5][6] + signed_kernel[0][1] ~^ image[5][7] + signed_kernel[0][2] ~^ image[5][8] + signed_kernel[0][3] ~^ image[5][9] + signed_kernel[0][4] ~^ image[5][10] + signed_kernel[1][0] ~^ image[6][6] + signed_kernel[1][1] ~^ image[6][7] + signed_kernel[1][2] ~^ image[6][8] + signed_kernel[1][3] ~^ image[6][9] + signed_kernel[1][4] ~^ image[6][10] + signed_kernel[2][0] ~^ image[7][6] + signed_kernel[2][1] ~^ image[7][7] + signed_kernel[2][2] ~^ image[7][8] + signed_kernel[2][3] ~^ image[7][9] + signed_kernel[2][4] ~^ image[7][10] + signed_kernel[3][0] ~^ image[8][6] + signed_kernel[3][1] ~^ image[8][7] + signed_kernel[3][2] ~^ image[8][8] + signed_kernel[3][3] ~^ image[8][9] + signed_kernel[3][4] ~^ image[8][10] + signed_kernel[4][0] ~^ image[9][6] + signed_kernel[4][1] ~^ image[9][7] + signed_kernel[4][2] ~^ image[9][8] + signed_kernel[4][3] ~^ image[9][9] + signed_kernel[4][4] ~^ image[9][10];
assign xor_sum[5][7] = signed_kernel[0][0] ~^ image[5][7] + signed_kernel[0][1] ~^ image[5][8] + signed_kernel[0][2] ~^ image[5][9] + signed_kernel[0][3] ~^ image[5][10] + signed_kernel[0][4] ~^ image[5][11] + signed_kernel[1][0] ~^ image[6][7] + signed_kernel[1][1] ~^ image[6][8] + signed_kernel[1][2] ~^ image[6][9] + signed_kernel[1][3] ~^ image[6][10] + signed_kernel[1][4] ~^ image[6][11] + signed_kernel[2][0] ~^ image[7][7] + signed_kernel[2][1] ~^ image[7][8] + signed_kernel[2][2] ~^ image[7][9] + signed_kernel[2][3] ~^ image[7][10] + signed_kernel[2][4] ~^ image[7][11] + signed_kernel[3][0] ~^ image[8][7] + signed_kernel[3][1] ~^ image[8][8] + signed_kernel[3][2] ~^ image[8][9] + signed_kernel[3][3] ~^ image[8][10] + signed_kernel[3][4] ~^ image[8][11] + signed_kernel[4][0] ~^ image[9][7] + signed_kernel[4][1] ~^ image[9][8] + signed_kernel[4][2] ~^ image[9][9] + signed_kernel[4][3] ~^ image[9][10] + signed_kernel[4][4] ~^ image[9][11];
assign xor_sum[5][8] = signed_kernel[0][0] ~^ image[5][8] + signed_kernel[0][1] ~^ image[5][9] + signed_kernel[0][2] ~^ image[5][10] + signed_kernel[0][3] ~^ image[5][11] + signed_kernel[0][4] ~^ image[5][12] + signed_kernel[1][0] ~^ image[6][8] + signed_kernel[1][1] ~^ image[6][9] + signed_kernel[1][2] ~^ image[6][10] + signed_kernel[1][3] ~^ image[6][11] + signed_kernel[1][4] ~^ image[6][12] + signed_kernel[2][0] ~^ image[7][8] + signed_kernel[2][1] ~^ image[7][9] + signed_kernel[2][2] ~^ image[7][10] + signed_kernel[2][3] ~^ image[7][11] + signed_kernel[2][4] ~^ image[7][12] + signed_kernel[3][0] ~^ image[8][8] + signed_kernel[3][1] ~^ image[8][9] + signed_kernel[3][2] ~^ image[8][10] + signed_kernel[3][3] ~^ image[8][11] + signed_kernel[3][4] ~^ image[8][12] + signed_kernel[4][0] ~^ image[9][8] + signed_kernel[4][1] ~^ image[9][9] + signed_kernel[4][2] ~^ image[9][10] + signed_kernel[4][3] ~^ image[9][11] + signed_kernel[4][4] ~^ image[9][12];
assign xor_sum[5][9] = signed_kernel[0][0] ~^ image[5][9] + signed_kernel[0][1] ~^ image[5][10] + signed_kernel[0][2] ~^ image[5][11] + signed_kernel[0][3] ~^ image[5][12] + signed_kernel[0][4] ~^ image[5][13] + signed_kernel[1][0] ~^ image[6][9] + signed_kernel[1][1] ~^ image[6][10] + signed_kernel[1][2] ~^ image[6][11] + signed_kernel[1][3] ~^ image[6][12] + signed_kernel[1][4] ~^ image[6][13] + signed_kernel[2][0] ~^ image[7][9] + signed_kernel[2][1] ~^ image[7][10] + signed_kernel[2][2] ~^ image[7][11] + signed_kernel[2][3] ~^ image[7][12] + signed_kernel[2][4] ~^ image[7][13] + signed_kernel[3][0] ~^ image[8][9] + signed_kernel[3][1] ~^ image[8][10] + signed_kernel[3][2] ~^ image[8][11] + signed_kernel[3][3] ~^ image[8][12] + signed_kernel[3][4] ~^ image[8][13] + signed_kernel[4][0] ~^ image[9][9] + signed_kernel[4][1] ~^ image[9][10] + signed_kernel[4][2] ~^ image[9][11] + signed_kernel[4][3] ~^ image[9][12] + signed_kernel[4][4] ~^ image[9][13];
assign xor_sum[5][10] = signed_kernel[0][0] ~^ image[5][10] + signed_kernel[0][1] ~^ image[5][11] + signed_kernel[0][2] ~^ image[5][12] + signed_kernel[0][3] ~^ image[5][13] + signed_kernel[0][4] ~^ image[5][14] + signed_kernel[1][0] ~^ image[6][10] + signed_kernel[1][1] ~^ image[6][11] + signed_kernel[1][2] ~^ image[6][12] + signed_kernel[1][3] ~^ image[6][13] + signed_kernel[1][4] ~^ image[6][14] + signed_kernel[2][0] ~^ image[7][10] + signed_kernel[2][1] ~^ image[7][11] + signed_kernel[2][2] ~^ image[7][12] + signed_kernel[2][3] ~^ image[7][13] + signed_kernel[2][4] ~^ image[7][14] + signed_kernel[3][0] ~^ image[8][10] + signed_kernel[3][1] ~^ image[8][11] + signed_kernel[3][2] ~^ image[8][12] + signed_kernel[3][3] ~^ image[8][13] + signed_kernel[3][4] ~^ image[8][14] + signed_kernel[4][0] ~^ image[9][10] + signed_kernel[4][1] ~^ image[9][11] + signed_kernel[4][2] ~^ image[9][12] + signed_kernel[4][3] ~^ image[9][13] + signed_kernel[4][4] ~^ image[9][14];
assign xor_sum[5][11] = signed_kernel[0][0] ~^ image[5][11] + signed_kernel[0][1] ~^ image[5][12] + signed_kernel[0][2] ~^ image[5][13] + signed_kernel[0][3] ~^ image[5][14] + signed_kernel[0][4] ~^ image[5][15] + signed_kernel[1][0] ~^ image[6][11] + signed_kernel[1][1] ~^ image[6][12] + signed_kernel[1][2] ~^ image[6][13] + signed_kernel[1][3] ~^ image[6][14] + signed_kernel[1][4] ~^ image[6][15] + signed_kernel[2][0] ~^ image[7][11] + signed_kernel[2][1] ~^ image[7][12] + signed_kernel[2][2] ~^ image[7][13] + signed_kernel[2][3] ~^ image[7][14] + signed_kernel[2][4] ~^ image[7][15] + signed_kernel[3][0] ~^ image[8][11] + signed_kernel[3][1] ~^ image[8][12] + signed_kernel[3][2] ~^ image[8][13] + signed_kernel[3][3] ~^ image[8][14] + signed_kernel[3][4] ~^ image[8][15] + signed_kernel[4][0] ~^ image[9][11] + signed_kernel[4][1] ~^ image[9][12] + signed_kernel[4][2] ~^ image[9][13] + signed_kernel[4][3] ~^ image[9][14] + signed_kernel[4][4] ~^ image[9][15];
assign xor_sum[5][12] = signed_kernel[0][0] ~^ image[5][12] + signed_kernel[0][1] ~^ image[5][13] + signed_kernel[0][2] ~^ image[5][14] + signed_kernel[0][3] ~^ image[5][15] + signed_kernel[0][4] ~^ image[5][16] + signed_kernel[1][0] ~^ image[6][12] + signed_kernel[1][1] ~^ image[6][13] + signed_kernel[1][2] ~^ image[6][14] + signed_kernel[1][3] ~^ image[6][15] + signed_kernel[1][4] ~^ image[6][16] + signed_kernel[2][0] ~^ image[7][12] + signed_kernel[2][1] ~^ image[7][13] + signed_kernel[2][2] ~^ image[7][14] + signed_kernel[2][3] ~^ image[7][15] + signed_kernel[2][4] ~^ image[7][16] + signed_kernel[3][0] ~^ image[8][12] + signed_kernel[3][1] ~^ image[8][13] + signed_kernel[3][2] ~^ image[8][14] + signed_kernel[3][3] ~^ image[8][15] + signed_kernel[3][4] ~^ image[8][16] + signed_kernel[4][0] ~^ image[9][12] + signed_kernel[4][1] ~^ image[9][13] + signed_kernel[4][2] ~^ image[9][14] + signed_kernel[4][3] ~^ image[9][15] + signed_kernel[4][4] ~^ image[9][16];
assign xor_sum[5][13] = signed_kernel[0][0] ~^ image[5][13] + signed_kernel[0][1] ~^ image[5][14] + signed_kernel[0][2] ~^ image[5][15] + signed_kernel[0][3] ~^ image[5][16] + signed_kernel[0][4] ~^ image[5][17] + signed_kernel[1][0] ~^ image[6][13] + signed_kernel[1][1] ~^ image[6][14] + signed_kernel[1][2] ~^ image[6][15] + signed_kernel[1][3] ~^ image[6][16] + signed_kernel[1][4] ~^ image[6][17] + signed_kernel[2][0] ~^ image[7][13] + signed_kernel[2][1] ~^ image[7][14] + signed_kernel[2][2] ~^ image[7][15] + signed_kernel[2][3] ~^ image[7][16] + signed_kernel[2][4] ~^ image[7][17] + signed_kernel[3][0] ~^ image[8][13] + signed_kernel[3][1] ~^ image[8][14] + signed_kernel[3][2] ~^ image[8][15] + signed_kernel[3][3] ~^ image[8][16] + signed_kernel[3][4] ~^ image[8][17] + signed_kernel[4][0] ~^ image[9][13] + signed_kernel[4][1] ~^ image[9][14] + signed_kernel[4][2] ~^ image[9][15] + signed_kernel[4][3] ~^ image[9][16] + signed_kernel[4][4] ~^ image[9][17];
assign xor_sum[5][14] = signed_kernel[0][0] ~^ image[5][14] + signed_kernel[0][1] ~^ image[5][15] + signed_kernel[0][2] ~^ image[5][16] + signed_kernel[0][3] ~^ image[5][17] + signed_kernel[0][4] ~^ image[5][18] + signed_kernel[1][0] ~^ image[6][14] + signed_kernel[1][1] ~^ image[6][15] + signed_kernel[1][2] ~^ image[6][16] + signed_kernel[1][3] ~^ image[6][17] + signed_kernel[1][4] ~^ image[6][18] + signed_kernel[2][0] ~^ image[7][14] + signed_kernel[2][1] ~^ image[7][15] + signed_kernel[2][2] ~^ image[7][16] + signed_kernel[2][3] ~^ image[7][17] + signed_kernel[2][4] ~^ image[7][18] + signed_kernel[3][0] ~^ image[8][14] + signed_kernel[3][1] ~^ image[8][15] + signed_kernel[3][2] ~^ image[8][16] + signed_kernel[3][3] ~^ image[8][17] + signed_kernel[3][4] ~^ image[8][18] + signed_kernel[4][0] ~^ image[9][14] + signed_kernel[4][1] ~^ image[9][15] + signed_kernel[4][2] ~^ image[9][16] + signed_kernel[4][3] ~^ image[9][17] + signed_kernel[4][4] ~^ image[9][18];
assign xor_sum[5][15] = signed_kernel[0][0] ~^ image[5][15] + signed_kernel[0][1] ~^ image[5][16] + signed_kernel[0][2] ~^ image[5][17] + signed_kernel[0][3] ~^ image[5][18] + signed_kernel[0][4] ~^ image[5][19] + signed_kernel[1][0] ~^ image[6][15] + signed_kernel[1][1] ~^ image[6][16] + signed_kernel[1][2] ~^ image[6][17] + signed_kernel[1][3] ~^ image[6][18] + signed_kernel[1][4] ~^ image[6][19] + signed_kernel[2][0] ~^ image[7][15] + signed_kernel[2][1] ~^ image[7][16] + signed_kernel[2][2] ~^ image[7][17] + signed_kernel[2][3] ~^ image[7][18] + signed_kernel[2][4] ~^ image[7][19] + signed_kernel[3][0] ~^ image[8][15] + signed_kernel[3][1] ~^ image[8][16] + signed_kernel[3][2] ~^ image[8][17] + signed_kernel[3][3] ~^ image[8][18] + signed_kernel[3][4] ~^ image[8][19] + signed_kernel[4][0] ~^ image[9][15] + signed_kernel[4][1] ~^ image[9][16] + signed_kernel[4][2] ~^ image[9][17] + signed_kernel[4][3] ~^ image[9][18] + signed_kernel[4][4] ~^ image[9][19];
assign xor_sum[5][16] = signed_kernel[0][0] ~^ image[5][16] + signed_kernel[0][1] ~^ image[5][17] + signed_kernel[0][2] ~^ image[5][18] + signed_kernel[0][3] ~^ image[5][19] + signed_kernel[0][4] ~^ image[5][20] + signed_kernel[1][0] ~^ image[6][16] + signed_kernel[1][1] ~^ image[6][17] + signed_kernel[1][2] ~^ image[6][18] + signed_kernel[1][3] ~^ image[6][19] + signed_kernel[1][4] ~^ image[6][20] + signed_kernel[2][0] ~^ image[7][16] + signed_kernel[2][1] ~^ image[7][17] + signed_kernel[2][2] ~^ image[7][18] + signed_kernel[2][3] ~^ image[7][19] + signed_kernel[2][4] ~^ image[7][20] + signed_kernel[3][0] ~^ image[8][16] + signed_kernel[3][1] ~^ image[8][17] + signed_kernel[3][2] ~^ image[8][18] + signed_kernel[3][3] ~^ image[8][19] + signed_kernel[3][4] ~^ image[8][20] + signed_kernel[4][0] ~^ image[9][16] + signed_kernel[4][1] ~^ image[9][17] + signed_kernel[4][2] ~^ image[9][18] + signed_kernel[4][3] ~^ image[9][19] + signed_kernel[4][4] ~^ image[9][20];
assign xor_sum[5][17] = signed_kernel[0][0] ~^ image[5][17] + signed_kernel[0][1] ~^ image[5][18] + signed_kernel[0][2] ~^ image[5][19] + signed_kernel[0][3] ~^ image[5][20] + signed_kernel[0][4] ~^ image[5][21] + signed_kernel[1][0] ~^ image[6][17] + signed_kernel[1][1] ~^ image[6][18] + signed_kernel[1][2] ~^ image[6][19] + signed_kernel[1][3] ~^ image[6][20] + signed_kernel[1][4] ~^ image[6][21] + signed_kernel[2][0] ~^ image[7][17] + signed_kernel[2][1] ~^ image[7][18] + signed_kernel[2][2] ~^ image[7][19] + signed_kernel[2][3] ~^ image[7][20] + signed_kernel[2][4] ~^ image[7][21] + signed_kernel[3][0] ~^ image[8][17] + signed_kernel[3][1] ~^ image[8][18] + signed_kernel[3][2] ~^ image[8][19] + signed_kernel[3][3] ~^ image[8][20] + signed_kernel[3][4] ~^ image[8][21] + signed_kernel[4][0] ~^ image[9][17] + signed_kernel[4][1] ~^ image[9][18] + signed_kernel[4][2] ~^ image[9][19] + signed_kernel[4][3] ~^ image[9][20] + signed_kernel[4][4] ~^ image[9][21];
assign xor_sum[5][18] = signed_kernel[0][0] ~^ image[5][18] + signed_kernel[0][1] ~^ image[5][19] + signed_kernel[0][2] ~^ image[5][20] + signed_kernel[0][3] ~^ image[5][21] + signed_kernel[0][4] ~^ image[5][22] + signed_kernel[1][0] ~^ image[6][18] + signed_kernel[1][1] ~^ image[6][19] + signed_kernel[1][2] ~^ image[6][20] + signed_kernel[1][3] ~^ image[6][21] + signed_kernel[1][4] ~^ image[6][22] + signed_kernel[2][0] ~^ image[7][18] + signed_kernel[2][1] ~^ image[7][19] + signed_kernel[2][2] ~^ image[7][20] + signed_kernel[2][3] ~^ image[7][21] + signed_kernel[2][4] ~^ image[7][22] + signed_kernel[3][0] ~^ image[8][18] + signed_kernel[3][1] ~^ image[8][19] + signed_kernel[3][2] ~^ image[8][20] + signed_kernel[3][3] ~^ image[8][21] + signed_kernel[3][4] ~^ image[8][22] + signed_kernel[4][0] ~^ image[9][18] + signed_kernel[4][1] ~^ image[9][19] + signed_kernel[4][2] ~^ image[9][20] + signed_kernel[4][3] ~^ image[9][21] + signed_kernel[4][4] ~^ image[9][22];
assign xor_sum[5][19] = signed_kernel[0][0] ~^ image[5][19] + signed_kernel[0][1] ~^ image[5][20] + signed_kernel[0][2] ~^ image[5][21] + signed_kernel[0][3] ~^ image[5][22] + signed_kernel[0][4] ~^ image[5][23] + signed_kernel[1][0] ~^ image[6][19] + signed_kernel[1][1] ~^ image[6][20] + signed_kernel[1][2] ~^ image[6][21] + signed_kernel[1][3] ~^ image[6][22] + signed_kernel[1][4] ~^ image[6][23] + signed_kernel[2][0] ~^ image[7][19] + signed_kernel[2][1] ~^ image[7][20] + signed_kernel[2][2] ~^ image[7][21] + signed_kernel[2][3] ~^ image[7][22] + signed_kernel[2][4] ~^ image[7][23] + signed_kernel[3][0] ~^ image[8][19] + signed_kernel[3][1] ~^ image[8][20] + signed_kernel[3][2] ~^ image[8][21] + signed_kernel[3][3] ~^ image[8][22] + signed_kernel[3][4] ~^ image[8][23] + signed_kernel[4][0] ~^ image[9][19] + signed_kernel[4][1] ~^ image[9][20] + signed_kernel[4][2] ~^ image[9][21] + signed_kernel[4][3] ~^ image[9][22] + signed_kernel[4][4] ~^ image[9][23];
assign xor_sum[5][20] = signed_kernel[0][0] ~^ image[5][20] + signed_kernel[0][1] ~^ image[5][21] + signed_kernel[0][2] ~^ image[5][22] + signed_kernel[0][3] ~^ image[5][23] + signed_kernel[0][4] ~^ image[5][24] + signed_kernel[1][0] ~^ image[6][20] + signed_kernel[1][1] ~^ image[6][21] + signed_kernel[1][2] ~^ image[6][22] + signed_kernel[1][3] ~^ image[6][23] + signed_kernel[1][4] ~^ image[6][24] + signed_kernel[2][0] ~^ image[7][20] + signed_kernel[2][1] ~^ image[7][21] + signed_kernel[2][2] ~^ image[7][22] + signed_kernel[2][3] ~^ image[7][23] + signed_kernel[2][4] ~^ image[7][24] + signed_kernel[3][0] ~^ image[8][20] + signed_kernel[3][1] ~^ image[8][21] + signed_kernel[3][2] ~^ image[8][22] + signed_kernel[3][3] ~^ image[8][23] + signed_kernel[3][4] ~^ image[8][24] + signed_kernel[4][0] ~^ image[9][20] + signed_kernel[4][1] ~^ image[9][21] + signed_kernel[4][2] ~^ image[9][22] + signed_kernel[4][3] ~^ image[9][23] + signed_kernel[4][4] ~^ image[9][24];
assign xor_sum[5][21] = signed_kernel[0][0] ~^ image[5][21] + signed_kernel[0][1] ~^ image[5][22] + signed_kernel[0][2] ~^ image[5][23] + signed_kernel[0][3] ~^ image[5][24] + signed_kernel[0][4] ~^ image[5][25] + signed_kernel[1][0] ~^ image[6][21] + signed_kernel[1][1] ~^ image[6][22] + signed_kernel[1][2] ~^ image[6][23] + signed_kernel[1][3] ~^ image[6][24] + signed_kernel[1][4] ~^ image[6][25] + signed_kernel[2][0] ~^ image[7][21] + signed_kernel[2][1] ~^ image[7][22] + signed_kernel[2][2] ~^ image[7][23] + signed_kernel[2][3] ~^ image[7][24] + signed_kernel[2][4] ~^ image[7][25] + signed_kernel[3][0] ~^ image[8][21] + signed_kernel[3][1] ~^ image[8][22] + signed_kernel[3][2] ~^ image[8][23] + signed_kernel[3][3] ~^ image[8][24] + signed_kernel[3][4] ~^ image[8][25] + signed_kernel[4][0] ~^ image[9][21] + signed_kernel[4][1] ~^ image[9][22] + signed_kernel[4][2] ~^ image[9][23] + signed_kernel[4][3] ~^ image[9][24] + signed_kernel[4][4] ~^ image[9][25];
assign xor_sum[5][22] = signed_kernel[0][0] ~^ image[5][22] + signed_kernel[0][1] ~^ image[5][23] + signed_kernel[0][2] ~^ image[5][24] + signed_kernel[0][3] ~^ image[5][25] + signed_kernel[0][4] ~^ image[5][26] + signed_kernel[1][0] ~^ image[6][22] + signed_kernel[1][1] ~^ image[6][23] + signed_kernel[1][2] ~^ image[6][24] + signed_kernel[1][3] ~^ image[6][25] + signed_kernel[1][4] ~^ image[6][26] + signed_kernel[2][0] ~^ image[7][22] + signed_kernel[2][1] ~^ image[7][23] + signed_kernel[2][2] ~^ image[7][24] + signed_kernel[2][3] ~^ image[7][25] + signed_kernel[2][4] ~^ image[7][26] + signed_kernel[3][0] ~^ image[8][22] + signed_kernel[3][1] ~^ image[8][23] + signed_kernel[3][2] ~^ image[8][24] + signed_kernel[3][3] ~^ image[8][25] + signed_kernel[3][4] ~^ image[8][26] + signed_kernel[4][0] ~^ image[9][22] + signed_kernel[4][1] ~^ image[9][23] + signed_kernel[4][2] ~^ image[9][24] + signed_kernel[4][3] ~^ image[9][25] + signed_kernel[4][4] ~^ image[9][26];
assign xor_sum[5][23] = signed_kernel[0][0] ~^ image[5][23] + signed_kernel[0][1] ~^ image[5][24] + signed_kernel[0][2] ~^ image[5][25] + signed_kernel[0][3] ~^ image[5][26] + signed_kernel[0][4] ~^ image[5][27] + signed_kernel[1][0] ~^ image[6][23] + signed_kernel[1][1] ~^ image[6][24] + signed_kernel[1][2] ~^ image[6][25] + signed_kernel[1][3] ~^ image[6][26] + signed_kernel[1][4] ~^ image[6][27] + signed_kernel[2][0] ~^ image[7][23] + signed_kernel[2][1] ~^ image[7][24] + signed_kernel[2][2] ~^ image[7][25] + signed_kernel[2][3] ~^ image[7][26] + signed_kernel[2][4] ~^ image[7][27] + signed_kernel[3][0] ~^ image[8][23] + signed_kernel[3][1] ~^ image[8][24] + signed_kernel[3][2] ~^ image[8][25] + signed_kernel[3][3] ~^ image[8][26] + signed_kernel[3][4] ~^ image[8][27] + signed_kernel[4][0] ~^ image[9][23] + signed_kernel[4][1] ~^ image[9][24] + signed_kernel[4][2] ~^ image[9][25] + signed_kernel[4][3] ~^ image[9][26] + signed_kernel[4][4] ~^ image[9][27];
assign xor_sum[6][0] = signed_kernel[0][0] ~^ image[6][0] + signed_kernel[0][1] ~^ image[6][1] + signed_kernel[0][2] ~^ image[6][2] + signed_kernel[0][3] ~^ image[6][3] + signed_kernel[0][4] ~^ image[6][4] + signed_kernel[1][0] ~^ image[7][0] + signed_kernel[1][1] ~^ image[7][1] + signed_kernel[1][2] ~^ image[7][2] + signed_kernel[1][3] ~^ image[7][3] + signed_kernel[1][4] ~^ image[7][4] + signed_kernel[2][0] ~^ image[8][0] + signed_kernel[2][1] ~^ image[8][1] + signed_kernel[2][2] ~^ image[8][2] + signed_kernel[2][3] ~^ image[8][3] + signed_kernel[2][4] ~^ image[8][4] + signed_kernel[3][0] ~^ image[9][0] + signed_kernel[3][1] ~^ image[9][1] + signed_kernel[3][2] ~^ image[9][2] + signed_kernel[3][3] ~^ image[9][3] + signed_kernel[3][4] ~^ image[9][4] + signed_kernel[4][0] ~^ image[10][0] + signed_kernel[4][1] ~^ image[10][1] + signed_kernel[4][2] ~^ image[10][2] + signed_kernel[4][3] ~^ image[10][3] + signed_kernel[4][4] ~^ image[10][4];
assign xor_sum[6][1] = signed_kernel[0][0] ~^ image[6][1] + signed_kernel[0][1] ~^ image[6][2] + signed_kernel[0][2] ~^ image[6][3] + signed_kernel[0][3] ~^ image[6][4] + signed_kernel[0][4] ~^ image[6][5] + signed_kernel[1][0] ~^ image[7][1] + signed_kernel[1][1] ~^ image[7][2] + signed_kernel[1][2] ~^ image[7][3] + signed_kernel[1][3] ~^ image[7][4] + signed_kernel[1][4] ~^ image[7][5] + signed_kernel[2][0] ~^ image[8][1] + signed_kernel[2][1] ~^ image[8][2] + signed_kernel[2][2] ~^ image[8][3] + signed_kernel[2][3] ~^ image[8][4] + signed_kernel[2][4] ~^ image[8][5] + signed_kernel[3][0] ~^ image[9][1] + signed_kernel[3][1] ~^ image[9][2] + signed_kernel[3][2] ~^ image[9][3] + signed_kernel[3][3] ~^ image[9][4] + signed_kernel[3][4] ~^ image[9][5] + signed_kernel[4][0] ~^ image[10][1] + signed_kernel[4][1] ~^ image[10][2] + signed_kernel[4][2] ~^ image[10][3] + signed_kernel[4][3] ~^ image[10][4] + signed_kernel[4][4] ~^ image[10][5];
assign xor_sum[6][2] = signed_kernel[0][0] ~^ image[6][2] + signed_kernel[0][1] ~^ image[6][3] + signed_kernel[0][2] ~^ image[6][4] + signed_kernel[0][3] ~^ image[6][5] + signed_kernel[0][4] ~^ image[6][6] + signed_kernel[1][0] ~^ image[7][2] + signed_kernel[1][1] ~^ image[7][3] + signed_kernel[1][2] ~^ image[7][4] + signed_kernel[1][3] ~^ image[7][5] + signed_kernel[1][4] ~^ image[7][6] + signed_kernel[2][0] ~^ image[8][2] + signed_kernel[2][1] ~^ image[8][3] + signed_kernel[2][2] ~^ image[8][4] + signed_kernel[2][3] ~^ image[8][5] + signed_kernel[2][4] ~^ image[8][6] + signed_kernel[3][0] ~^ image[9][2] + signed_kernel[3][1] ~^ image[9][3] + signed_kernel[3][2] ~^ image[9][4] + signed_kernel[3][3] ~^ image[9][5] + signed_kernel[3][4] ~^ image[9][6] + signed_kernel[4][0] ~^ image[10][2] + signed_kernel[4][1] ~^ image[10][3] + signed_kernel[4][2] ~^ image[10][4] + signed_kernel[4][3] ~^ image[10][5] + signed_kernel[4][4] ~^ image[10][6];
assign xor_sum[6][3] = signed_kernel[0][0] ~^ image[6][3] + signed_kernel[0][1] ~^ image[6][4] + signed_kernel[0][2] ~^ image[6][5] + signed_kernel[0][3] ~^ image[6][6] + signed_kernel[0][4] ~^ image[6][7] + signed_kernel[1][0] ~^ image[7][3] + signed_kernel[1][1] ~^ image[7][4] + signed_kernel[1][2] ~^ image[7][5] + signed_kernel[1][3] ~^ image[7][6] + signed_kernel[1][4] ~^ image[7][7] + signed_kernel[2][0] ~^ image[8][3] + signed_kernel[2][1] ~^ image[8][4] + signed_kernel[2][2] ~^ image[8][5] + signed_kernel[2][3] ~^ image[8][6] + signed_kernel[2][4] ~^ image[8][7] + signed_kernel[3][0] ~^ image[9][3] + signed_kernel[3][1] ~^ image[9][4] + signed_kernel[3][2] ~^ image[9][5] + signed_kernel[3][3] ~^ image[9][6] + signed_kernel[3][4] ~^ image[9][7] + signed_kernel[4][0] ~^ image[10][3] + signed_kernel[4][1] ~^ image[10][4] + signed_kernel[4][2] ~^ image[10][5] + signed_kernel[4][3] ~^ image[10][6] + signed_kernel[4][4] ~^ image[10][7];
assign xor_sum[6][4] = signed_kernel[0][0] ~^ image[6][4] + signed_kernel[0][1] ~^ image[6][5] + signed_kernel[0][2] ~^ image[6][6] + signed_kernel[0][3] ~^ image[6][7] + signed_kernel[0][4] ~^ image[6][8] + signed_kernel[1][0] ~^ image[7][4] + signed_kernel[1][1] ~^ image[7][5] + signed_kernel[1][2] ~^ image[7][6] + signed_kernel[1][3] ~^ image[7][7] + signed_kernel[1][4] ~^ image[7][8] + signed_kernel[2][0] ~^ image[8][4] + signed_kernel[2][1] ~^ image[8][5] + signed_kernel[2][2] ~^ image[8][6] + signed_kernel[2][3] ~^ image[8][7] + signed_kernel[2][4] ~^ image[8][8] + signed_kernel[3][0] ~^ image[9][4] + signed_kernel[3][1] ~^ image[9][5] + signed_kernel[3][2] ~^ image[9][6] + signed_kernel[3][3] ~^ image[9][7] + signed_kernel[3][4] ~^ image[9][8] + signed_kernel[4][0] ~^ image[10][4] + signed_kernel[4][1] ~^ image[10][5] + signed_kernel[4][2] ~^ image[10][6] + signed_kernel[4][3] ~^ image[10][7] + signed_kernel[4][4] ~^ image[10][8];
assign xor_sum[6][5] = signed_kernel[0][0] ~^ image[6][5] + signed_kernel[0][1] ~^ image[6][6] + signed_kernel[0][2] ~^ image[6][7] + signed_kernel[0][3] ~^ image[6][8] + signed_kernel[0][4] ~^ image[6][9] + signed_kernel[1][0] ~^ image[7][5] + signed_kernel[1][1] ~^ image[7][6] + signed_kernel[1][2] ~^ image[7][7] + signed_kernel[1][3] ~^ image[7][8] + signed_kernel[1][4] ~^ image[7][9] + signed_kernel[2][0] ~^ image[8][5] + signed_kernel[2][1] ~^ image[8][6] + signed_kernel[2][2] ~^ image[8][7] + signed_kernel[2][3] ~^ image[8][8] + signed_kernel[2][4] ~^ image[8][9] + signed_kernel[3][0] ~^ image[9][5] + signed_kernel[3][1] ~^ image[9][6] + signed_kernel[3][2] ~^ image[9][7] + signed_kernel[3][3] ~^ image[9][8] + signed_kernel[3][4] ~^ image[9][9] + signed_kernel[4][0] ~^ image[10][5] + signed_kernel[4][1] ~^ image[10][6] + signed_kernel[4][2] ~^ image[10][7] + signed_kernel[4][3] ~^ image[10][8] + signed_kernel[4][4] ~^ image[10][9];
assign xor_sum[6][6] = signed_kernel[0][0] ~^ image[6][6] + signed_kernel[0][1] ~^ image[6][7] + signed_kernel[0][2] ~^ image[6][8] + signed_kernel[0][3] ~^ image[6][9] + signed_kernel[0][4] ~^ image[6][10] + signed_kernel[1][0] ~^ image[7][6] + signed_kernel[1][1] ~^ image[7][7] + signed_kernel[1][2] ~^ image[7][8] + signed_kernel[1][3] ~^ image[7][9] + signed_kernel[1][4] ~^ image[7][10] + signed_kernel[2][0] ~^ image[8][6] + signed_kernel[2][1] ~^ image[8][7] + signed_kernel[2][2] ~^ image[8][8] + signed_kernel[2][3] ~^ image[8][9] + signed_kernel[2][4] ~^ image[8][10] + signed_kernel[3][0] ~^ image[9][6] + signed_kernel[3][1] ~^ image[9][7] + signed_kernel[3][2] ~^ image[9][8] + signed_kernel[3][3] ~^ image[9][9] + signed_kernel[3][4] ~^ image[9][10] + signed_kernel[4][0] ~^ image[10][6] + signed_kernel[4][1] ~^ image[10][7] + signed_kernel[4][2] ~^ image[10][8] + signed_kernel[4][3] ~^ image[10][9] + signed_kernel[4][4] ~^ image[10][10];
assign xor_sum[6][7] = signed_kernel[0][0] ~^ image[6][7] + signed_kernel[0][1] ~^ image[6][8] + signed_kernel[0][2] ~^ image[6][9] + signed_kernel[0][3] ~^ image[6][10] + signed_kernel[0][4] ~^ image[6][11] + signed_kernel[1][0] ~^ image[7][7] + signed_kernel[1][1] ~^ image[7][8] + signed_kernel[1][2] ~^ image[7][9] + signed_kernel[1][3] ~^ image[7][10] + signed_kernel[1][4] ~^ image[7][11] + signed_kernel[2][0] ~^ image[8][7] + signed_kernel[2][1] ~^ image[8][8] + signed_kernel[2][2] ~^ image[8][9] + signed_kernel[2][3] ~^ image[8][10] + signed_kernel[2][4] ~^ image[8][11] + signed_kernel[3][0] ~^ image[9][7] + signed_kernel[3][1] ~^ image[9][8] + signed_kernel[3][2] ~^ image[9][9] + signed_kernel[3][3] ~^ image[9][10] + signed_kernel[3][4] ~^ image[9][11] + signed_kernel[4][0] ~^ image[10][7] + signed_kernel[4][1] ~^ image[10][8] + signed_kernel[4][2] ~^ image[10][9] + signed_kernel[4][3] ~^ image[10][10] + signed_kernel[4][4] ~^ image[10][11];
assign xor_sum[6][8] = signed_kernel[0][0] ~^ image[6][8] + signed_kernel[0][1] ~^ image[6][9] + signed_kernel[0][2] ~^ image[6][10] + signed_kernel[0][3] ~^ image[6][11] + signed_kernel[0][4] ~^ image[6][12] + signed_kernel[1][0] ~^ image[7][8] + signed_kernel[1][1] ~^ image[7][9] + signed_kernel[1][2] ~^ image[7][10] + signed_kernel[1][3] ~^ image[7][11] + signed_kernel[1][4] ~^ image[7][12] + signed_kernel[2][0] ~^ image[8][8] + signed_kernel[2][1] ~^ image[8][9] + signed_kernel[2][2] ~^ image[8][10] + signed_kernel[2][3] ~^ image[8][11] + signed_kernel[2][4] ~^ image[8][12] + signed_kernel[3][0] ~^ image[9][8] + signed_kernel[3][1] ~^ image[9][9] + signed_kernel[3][2] ~^ image[9][10] + signed_kernel[3][3] ~^ image[9][11] + signed_kernel[3][4] ~^ image[9][12] + signed_kernel[4][0] ~^ image[10][8] + signed_kernel[4][1] ~^ image[10][9] + signed_kernel[4][2] ~^ image[10][10] + signed_kernel[4][3] ~^ image[10][11] + signed_kernel[4][4] ~^ image[10][12];
assign xor_sum[6][9] = signed_kernel[0][0] ~^ image[6][9] + signed_kernel[0][1] ~^ image[6][10] + signed_kernel[0][2] ~^ image[6][11] + signed_kernel[0][3] ~^ image[6][12] + signed_kernel[0][4] ~^ image[6][13] + signed_kernel[1][0] ~^ image[7][9] + signed_kernel[1][1] ~^ image[7][10] + signed_kernel[1][2] ~^ image[7][11] + signed_kernel[1][3] ~^ image[7][12] + signed_kernel[1][4] ~^ image[7][13] + signed_kernel[2][0] ~^ image[8][9] + signed_kernel[2][1] ~^ image[8][10] + signed_kernel[2][2] ~^ image[8][11] + signed_kernel[2][3] ~^ image[8][12] + signed_kernel[2][4] ~^ image[8][13] + signed_kernel[3][0] ~^ image[9][9] + signed_kernel[3][1] ~^ image[9][10] + signed_kernel[3][2] ~^ image[9][11] + signed_kernel[3][3] ~^ image[9][12] + signed_kernel[3][4] ~^ image[9][13] + signed_kernel[4][0] ~^ image[10][9] + signed_kernel[4][1] ~^ image[10][10] + signed_kernel[4][2] ~^ image[10][11] + signed_kernel[4][3] ~^ image[10][12] + signed_kernel[4][4] ~^ image[10][13];
assign xor_sum[6][10] = signed_kernel[0][0] ~^ image[6][10] + signed_kernel[0][1] ~^ image[6][11] + signed_kernel[0][2] ~^ image[6][12] + signed_kernel[0][3] ~^ image[6][13] + signed_kernel[0][4] ~^ image[6][14] + signed_kernel[1][0] ~^ image[7][10] + signed_kernel[1][1] ~^ image[7][11] + signed_kernel[1][2] ~^ image[7][12] + signed_kernel[1][3] ~^ image[7][13] + signed_kernel[1][4] ~^ image[7][14] + signed_kernel[2][0] ~^ image[8][10] + signed_kernel[2][1] ~^ image[8][11] + signed_kernel[2][2] ~^ image[8][12] + signed_kernel[2][3] ~^ image[8][13] + signed_kernel[2][4] ~^ image[8][14] + signed_kernel[3][0] ~^ image[9][10] + signed_kernel[3][1] ~^ image[9][11] + signed_kernel[3][2] ~^ image[9][12] + signed_kernel[3][3] ~^ image[9][13] + signed_kernel[3][4] ~^ image[9][14] + signed_kernel[4][0] ~^ image[10][10] + signed_kernel[4][1] ~^ image[10][11] + signed_kernel[4][2] ~^ image[10][12] + signed_kernel[4][3] ~^ image[10][13] + signed_kernel[4][4] ~^ image[10][14];
assign xor_sum[6][11] = signed_kernel[0][0] ~^ image[6][11] + signed_kernel[0][1] ~^ image[6][12] + signed_kernel[0][2] ~^ image[6][13] + signed_kernel[0][3] ~^ image[6][14] + signed_kernel[0][4] ~^ image[6][15] + signed_kernel[1][0] ~^ image[7][11] + signed_kernel[1][1] ~^ image[7][12] + signed_kernel[1][2] ~^ image[7][13] + signed_kernel[1][3] ~^ image[7][14] + signed_kernel[1][4] ~^ image[7][15] + signed_kernel[2][0] ~^ image[8][11] + signed_kernel[2][1] ~^ image[8][12] + signed_kernel[2][2] ~^ image[8][13] + signed_kernel[2][3] ~^ image[8][14] + signed_kernel[2][4] ~^ image[8][15] + signed_kernel[3][0] ~^ image[9][11] + signed_kernel[3][1] ~^ image[9][12] + signed_kernel[3][2] ~^ image[9][13] + signed_kernel[3][3] ~^ image[9][14] + signed_kernel[3][4] ~^ image[9][15] + signed_kernel[4][0] ~^ image[10][11] + signed_kernel[4][1] ~^ image[10][12] + signed_kernel[4][2] ~^ image[10][13] + signed_kernel[4][3] ~^ image[10][14] + signed_kernel[4][4] ~^ image[10][15];
assign xor_sum[6][12] = signed_kernel[0][0] ~^ image[6][12] + signed_kernel[0][1] ~^ image[6][13] + signed_kernel[0][2] ~^ image[6][14] + signed_kernel[0][3] ~^ image[6][15] + signed_kernel[0][4] ~^ image[6][16] + signed_kernel[1][0] ~^ image[7][12] + signed_kernel[1][1] ~^ image[7][13] + signed_kernel[1][2] ~^ image[7][14] + signed_kernel[1][3] ~^ image[7][15] + signed_kernel[1][4] ~^ image[7][16] + signed_kernel[2][0] ~^ image[8][12] + signed_kernel[2][1] ~^ image[8][13] + signed_kernel[2][2] ~^ image[8][14] + signed_kernel[2][3] ~^ image[8][15] + signed_kernel[2][4] ~^ image[8][16] + signed_kernel[3][0] ~^ image[9][12] + signed_kernel[3][1] ~^ image[9][13] + signed_kernel[3][2] ~^ image[9][14] + signed_kernel[3][3] ~^ image[9][15] + signed_kernel[3][4] ~^ image[9][16] + signed_kernel[4][0] ~^ image[10][12] + signed_kernel[4][1] ~^ image[10][13] + signed_kernel[4][2] ~^ image[10][14] + signed_kernel[4][3] ~^ image[10][15] + signed_kernel[4][4] ~^ image[10][16];
assign xor_sum[6][13] = signed_kernel[0][0] ~^ image[6][13] + signed_kernel[0][1] ~^ image[6][14] + signed_kernel[0][2] ~^ image[6][15] + signed_kernel[0][3] ~^ image[6][16] + signed_kernel[0][4] ~^ image[6][17] + signed_kernel[1][0] ~^ image[7][13] + signed_kernel[1][1] ~^ image[7][14] + signed_kernel[1][2] ~^ image[7][15] + signed_kernel[1][3] ~^ image[7][16] + signed_kernel[1][4] ~^ image[7][17] + signed_kernel[2][0] ~^ image[8][13] + signed_kernel[2][1] ~^ image[8][14] + signed_kernel[2][2] ~^ image[8][15] + signed_kernel[2][3] ~^ image[8][16] + signed_kernel[2][4] ~^ image[8][17] + signed_kernel[3][0] ~^ image[9][13] + signed_kernel[3][1] ~^ image[9][14] + signed_kernel[3][2] ~^ image[9][15] + signed_kernel[3][3] ~^ image[9][16] + signed_kernel[3][4] ~^ image[9][17] + signed_kernel[4][0] ~^ image[10][13] + signed_kernel[4][1] ~^ image[10][14] + signed_kernel[4][2] ~^ image[10][15] + signed_kernel[4][3] ~^ image[10][16] + signed_kernel[4][4] ~^ image[10][17];
assign xor_sum[6][14] = signed_kernel[0][0] ~^ image[6][14] + signed_kernel[0][1] ~^ image[6][15] + signed_kernel[0][2] ~^ image[6][16] + signed_kernel[0][3] ~^ image[6][17] + signed_kernel[0][4] ~^ image[6][18] + signed_kernel[1][0] ~^ image[7][14] + signed_kernel[1][1] ~^ image[7][15] + signed_kernel[1][2] ~^ image[7][16] + signed_kernel[1][3] ~^ image[7][17] + signed_kernel[1][4] ~^ image[7][18] + signed_kernel[2][0] ~^ image[8][14] + signed_kernel[2][1] ~^ image[8][15] + signed_kernel[2][2] ~^ image[8][16] + signed_kernel[2][3] ~^ image[8][17] + signed_kernel[2][4] ~^ image[8][18] + signed_kernel[3][0] ~^ image[9][14] + signed_kernel[3][1] ~^ image[9][15] + signed_kernel[3][2] ~^ image[9][16] + signed_kernel[3][3] ~^ image[9][17] + signed_kernel[3][4] ~^ image[9][18] + signed_kernel[4][0] ~^ image[10][14] + signed_kernel[4][1] ~^ image[10][15] + signed_kernel[4][2] ~^ image[10][16] + signed_kernel[4][3] ~^ image[10][17] + signed_kernel[4][4] ~^ image[10][18];
assign xor_sum[6][15] = signed_kernel[0][0] ~^ image[6][15] + signed_kernel[0][1] ~^ image[6][16] + signed_kernel[0][2] ~^ image[6][17] + signed_kernel[0][3] ~^ image[6][18] + signed_kernel[0][4] ~^ image[6][19] + signed_kernel[1][0] ~^ image[7][15] + signed_kernel[1][1] ~^ image[7][16] + signed_kernel[1][2] ~^ image[7][17] + signed_kernel[1][3] ~^ image[7][18] + signed_kernel[1][4] ~^ image[7][19] + signed_kernel[2][0] ~^ image[8][15] + signed_kernel[2][1] ~^ image[8][16] + signed_kernel[2][2] ~^ image[8][17] + signed_kernel[2][3] ~^ image[8][18] + signed_kernel[2][4] ~^ image[8][19] + signed_kernel[3][0] ~^ image[9][15] + signed_kernel[3][1] ~^ image[9][16] + signed_kernel[3][2] ~^ image[9][17] + signed_kernel[3][3] ~^ image[9][18] + signed_kernel[3][4] ~^ image[9][19] + signed_kernel[4][0] ~^ image[10][15] + signed_kernel[4][1] ~^ image[10][16] + signed_kernel[4][2] ~^ image[10][17] + signed_kernel[4][3] ~^ image[10][18] + signed_kernel[4][4] ~^ image[10][19];
assign xor_sum[6][16] = signed_kernel[0][0] ~^ image[6][16] + signed_kernel[0][1] ~^ image[6][17] + signed_kernel[0][2] ~^ image[6][18] + signed_kernel[0][3] ~^ image[6][19] + signed_kernel[0][4] ~^ image[6][20] + signed_kernel[1][0] ~^ image[7][16] + signed_kernel[1][1] ~^ image[7][17] + signed_kernel[1][2] ~^ image[7][18] + signed_kernel[1][3] ~^ image[7][19] + signed_kernel[1][4] ~^ image[7][20] + signed_kernel[2][0] ~^ image[8][16] + signed_kernel[2][1] ~^ image[8][17] + signed_kernel[2][2] ~^ image[8][18] + signed_kernel[2][3] ~^ image[8][19] + signed_kernel[2][4] ~^ image[8][20] + signed_kernel[3][0] ~^ image[9][16] + signed_kernel[3][1] ~^ image[9][17] + signed_kernel[3][2] ~^ image[9][18] + signed_kernel[3][3] ~^ image[9][19] + signed_kernel[3][4] ~^ image[9][20] + signed_kernel[4][0] ~^ image[10][16] + signed_kernel[4][1] ~^ image[10][17] + signed_kernel[4][2] ~^ image[10][18] + signed_kernel[4][3] ~^ image[10][19] + signed_kernel[4][4] ~^ image[10][20];
assign xor_sum[6][17] = signed_kernel[0][0] ~^ image[6][17] + signed_kernel[0][1] ~^ image[6][18] + signed_kernel[0][2] ~^ image[6][19] + signed_kernel[0][3] ~^ image[6][20] + signed_kernel[0][4] ~^ image[6][21] + signed_kernel[1][0] ~^ image[7][17] + signed_kernel[1][1] ~^ image[7][18] + signed_kernel[1][2] ~^ image[7][19] + signed_kernel[1][3] ~^ image[7][20] + signed_kernel[1][4] ~^ image[7][21] + signed_kernel[2][0] ~^ image[8][17] + signed_kernel[2][1] ~^ image[8][18] + signed_kernel[2][2] ~^ image[8][19] + signed_kernel[2][3] ~^ image[8][20] + signed_kernel[2][4] ~^ image[8][21] + signed_kernel[3][0] ~^ image[9][17] + signed_kernel[3][1] ~^ image[9][18] + signed_kernel[3][2] ~^ image[9][19] + signed_kernel[3][3] ~^ image[9][20] + signed_kernel[3][4] ~^ image[9][21] + signed_kernel[4][0] ~^ image[10][17] + signed_kernel[4][1] ~^ image[10][18] + signed_kernel[4][2] ~^ image[10][19] + signed_kernel[4][3] ~^ image[10][20] + signed_kernel[4][4] ~^ image[10][21];
assign xor_sum[6][18] = signed_kernel[0][0] ~^ image[6][18] + signed_kernel[0][1] ~^ image[6][19] + signed_kernel[0][2] ~^ image[6][20] + signed_kernel[0][3] ~^ image[6][21] + signed_kernel[0][4] ~^ image[6][22] + signed_kernel[1][0] ~^ image[7][18] + signed_kernel[1][1] ~^ image[7][19] + signed_kernel[1][2] ~^ image[7][20] + signed_kernel[1][3] ~^ image[7][21] + signed_kernel[1][4] ~^ image[7][22] + signed_kernel[2][0] ~^ image[8][18] + signed_kernel[2][1] ~^ image[8][19] + signed_kernel[2][2] ~^ image[8][20] + signed_kernel[2][3] ~^ image[8][21] + signed_kernel[2][4] ~^ image[8][22] + signed_kernel[3][0] ~^ image[9][18] + signed_kernel[3][1] ~^ image[9][19] + signed_kernel[3][2] ~^ image[9][20] + signed_kernel[3][3] ~^ image[9][21] + signed_kernel[3][4] ~^ image[9][22] + signed_kernel[4][0] ~^ image[10][18] + signed_kernel[4][1] ~^ image[10][19] + signed_kernel[4][2] ~^ image[10][20] + signed_kernel[4][3] ~^ image[10][21] + signed_kernel[4][4] ~^ image[10][22];
assign xor_sum[6][19] = signed_kernel[0][0] ~^ image[6][19] + signed_kernel[0][1] ~^ image[6][20] + signed_kernel[0][2] ~^ image[6][21] + signed_kernel[0][3] ~^ image[6][22] + signed_kernel[0][4] ~^ image[6][23] + signed_kernel[1][0] ~^ image[7][19] + signed_kernel[1][1] ~^ image[7][20] + signed_kernel[1][2] ~^ image[7][21] + signed_kernel[1][3] ~^ image[7][22] + signed_kernel[1][4] ~^ image[7][23] + signed_kernel[2][0] ~^ image[8][19] + signed_kernel[2][1] ~^ image[8][20] + signed_kernel[2][2] ~^ image[8][21] + signed_kernel[2][3] ~^ image[8][22] + signed_kernel[2][4] ~^ image[8][23] + signed_kernel[3][0] ~^ image[9][19] + signed_kernel[3][1] ~^ image[9][20] + signed_kernel[3][2] ~^ image[9][21] + signed_kernel[3][3] ~^ image[9][22] + signed_kernel[3][4] ~^ image[9][23] + signed_kernel[4][0] ~^ image[10][19] + signed_kernel[4][1] ~^ image[10][20] + signed_kernel[4][2] ~^ image[10][21] + signed_kernel[4][3] ~^ image[10][22] + signed_kernel[4][4] ~^ image[10][23];
assign xor_sum[6][20] = signed_kernel[0][0] ~^ image[6][20] + signed_kernel[0][1] ~^ image[6][21] + signed_kernel[0][2] ~^ image[6][22] + signed_kernel[0][3] ~^ image[6][23] + signed_kernel[0][4] ~^ image[6][24] + signed_kernel[1][0] ~^ image[7][20] + signed_kernel[1][1] ~^ image[7][21] + signed_kernel[1][2] ~^ image[7][22] + signed_kernel[1][3] ~^ image[7][23] + signed_kernel[1][4] ~^ image[7][24] + signed_kernel[2][0] ~^ image[8][20] + signed_kernel[2][1] ~^ image[8][21] + signed_kernel[2][2] ~^ image[8][22] + signed_kernel[2][3] ~^ image[8][23] + signed_kernel[2][4] ~^ image[8][24] + signed_kernel[3][0] ~^ image[9][20] + signed_kernel[3][1] ~^ image[9][21] + signed_kernel[3][2] ~^ image[9][22] + signed_kernel[3][3] ~^ image[9][23] + signed_kernel[3][4] ~^ image[9][24] + signed_kernel[4][0] ~^ image[10][20] + signed_kernel[4][1] ~^ image[10][21] + signed_kernel[4][2] ~^ image[10][22] + signed_kernel[4][3] ~^ image[10][23] + signed_kernel[4][4] ~^ image[10][24];
assign xor_sum[6][21] = signed_kernel[0][0] ~^ image[6][21] + signed_kernel[0][1] ~^ image[6][22] + signed_kernel[0][2] ~^ image[6][23] + signed_kernel[0][3] ~^ image[6][24] + signed_kernel[0][4] ~^ image[6][25] + signed_kernel[1][0] ~^ image[7][21] + signed_kernel[1][1] ~^ image[7][22] + signed_kernel[1][2] ~^ image[7][23] + signed_kernel[1][3] ~^ image[7][24] + signed_kernel[1][4] ~^ image[7][25] + signed_kernel[2][0] ~^ image[8][21] + signed_kernel[2][1] ~^ image[8][22] + signed_kernel[2][2] ~^ image[8][23] + signed_kernel[2][3] ~^ image[8][24] + signed_kernel[2][4] ~^ image[8][25] + signed_kernel[3][0] ~^ image[9][21] + signed_kernel[3][1] ~^ image[9][22] + signed_kernel[3][2] ~^ image[9][23] + signed_kernel[3][3] ~^ image[9][24] + signed_kernel[3][4] ~^ image[9][25] + signed_kernel[4][0] ~^ image[10][21] + signed_kernel[4][1] ~^ image[10][22] + signed_kernel[4][2] ~^ image[10][23] + signed_kernel[4][3] ~^ image[10][24] + signed_kernel[4][4] ~^ image[10][25];
assign xor_sum[6][22] = signed_kernel[0][0] ~^ image[6][22] + signed_kernel[0][1] ~^ image[6][23] + signed_kernel[0][2] ~^ image[6][24] + signed_kernel[0][3] ~^ image[6][25] + signed_kernel[0][4] ~^ image[6][26] + signed_kernel[1][0] ~^ image[7][22] + signed_kernel[1][1] ~^ image[7][23] + signed_kernel[1][2] ~^ image[7][24] + signed_kernel[1][3] ~^ image[7][25] + signed_kernel[1][4] ~^ image[7][26] + signed_kernel[2][0] ~^ image[8][22] + signed_kernel[2][1] ~^ image[8][23] + signed_kernel[2][2] ~^ image[8][24] + signed_kernel[2][3] ~^ image[8][25] + signed_kernel[2][4] ~^ image[8][26] + signed_kernel[3][0] ~^ image[9][22] + signed_kernel[3][1] ~^ image[9][23] + signed_kernel[3][2] ~^ image[9][24] + signed_kernel[3][3] ~^ image[9][25] + signed_kernel[3][4] ~^ image[9][26] + signed_kernel[4][0] ~^ image[10][22] + signed_kernel[4][1] ~^ image[10][23] + signed_kernel[4][2] ~^ image[10][24] + signed_kernel[4][3] ~^ image[10][25] + signed_kernel[4][4] ~^ image[10][26];
assign xor_sum[6][23] = signed_kernel[0][0] ~^ image[6][23] + signed_kernel[0][1] ~^ image[6][24] + signed_kernel[0][2] ~^ image[6][25] + signed_kernel[0][3] ~^ image[6][26] + signed_kernel[0][4] ~^ image[6][27] + signed_kernel[1][0] ~^ image[7][23] + signed_kernel[1][1] ~^ image[7][24] + signed_kernel[1][2] ~^ image[7][25] + signed_kernel[1][3] ~^ image[7][26] + signed_kernel[1][4] ~^ image[7][27] + signed_kernel[2][0] ~^ image[8][23] + signed_kernel[2][1] ~^ image[8][24] + signed_kernel[2][2] ~^ image[8][25] + signed_kernel[2][3] ~^ image[8][26] + signed_kernel[2][4] ~^ image[8][27] + signed_kernel[3][0] ~^ image[9][23] + signed_kernel[3][1] ~^ image[9][24] + signed_kernel[3][2] ~^ image[9][25] + signed_kernel[3][3] ~^ image[9][26] + signed_kernel[3][4] ~^ image[9][27] + signed_kernel[4][0] ~^ image[10][23] + signed_kernel[4][1] ~^ image[10][24] + signed_kernel[4][2] ~^ image[10][25] + signed_kernel[4][3] ~^ image[10][26] + signed_kernel[4][4] ~^ image[10][27];
assign xor_sum[7][0] = signed_kernel[0][0] ~^ image[7][0] + signed_kernel[0][1] ~^ image[7][1] + signed_kernel[0][2] ~^ image[7][2] + signed_kernel[0][3] ~^ image[7][3] + signed_kernel[0][4] ~^ image[7][4] + signed_kernel[1][0] ~^ image[8][0] + signed_kernel[1][1] ~^ image[8][1] + signed_kernel[1][2] ~^ image[8][2] + signed_kernel[1][3] ~^ image[8][3] + signed_kernel[1][4] ~^ image[8][4] + signed_kernel[2][0] ~^ image[9][0] + signed_kernel[2][1] ~^ image[9][1] + signed_kernel[2][2] ~^ image[9][2] + signed_kernel[2][3] ~^ image[9][3] + signed_kernel[2][4] ~^ image[9][4] + signed_kernel[3][0] ~^ image[10][0] + signed_kernel[3][1] ~^ image[10][1] + signed_kernel[3][2] ~^ image[10][2] + signed_kernel[3][3] ~^ image[10][3] + signed_kernel[3][4] ~^ image[10][4] + signed_kernel[4][0] ~^ image[11][0] + signed_kernel[4][1] ~^ image[11][1] + signed_kernel[4][2] ~^ image[11][2] + signed_kernel[4][3] ~^ image[11][3] + signed_kernel[4][4] ~^ image[11][4];
assign xor_sum[7][1] = signed_kernel[0][0] ~^ image[7][1] + signed_kernel[0][1] ~^ image[7][2] + signed_kernel[0][2] ~^ image[7][3] + signed_kernel[0][3] ~^ image[7][4] + signed_kernel[0][4] ~^ image[7][5] + signed_kernel[1][0] ~^ image[8][1] + signed_kernel[1][1] ~^ image[8][2] + signed_kernel[1][2] ~^ image[8][3] + signed_kernel[1][3] ~^ image[8][4] + signed_kernel[1][4] ~^ image[8][5] + signed_kernel[2][0] ~^ image[9][1] + signed_kernel[2][1] ~^ image[9][2] + signed_kernel[2][2] ~^ image[9][3] + signed_kernel[2][3] ~^ image[9][4] + signed_kernel[2][4] ~^ image[9][5] + signed_kernel[3][0] ~^ image[10][1] + signed_kernel[3][1] ~^ image[10][2] + signed_kernel[3][2] ~^ image[10][3] + signed_kernel[3][3] ~^ image[10][4] + signed_kernel[3][4] ~^ image[10][5] + signed_kernel[4][0] ~^ image[11][1] + signed_kernel[4][1] ~^ image[11][2] + signed_kernel[4][2] ~^ image[11][3] + signed_kernel[4][3] ~^ image[11][4] + signed_kernel[4][4] ~^ image[11][5];
assign xor_sum[7][2] = signed_kernel[0][0] ~^ image[7][2] + signed_kernel[0][1] ~^ image[7][3] + signed_kernel[0][2] ~^ image[7][4] + signed_kernel[0][3] ~^ image[7][5] + signed_kernel[0][4] ~^ image[7][6] + signed_kernel[1][0] ~^ image[8][2] + signed_kernel[1][1] ~^ image[8][3] + signed_kernel[1][2] ~^ image[8][4] + signed_kernel[1][3] ~^ image[8][5] + signed_kernel[1][4] ~^ image[8][6] + signed_kernel[2][0] ~^ image[9][2] + signed_kernel[2][1] ~^ image[9][3] + signed_kernel[2][2] ~^ image[9][4] + signed_kernel[2][3] ~^ image[9][5] + signed_kernel[2][4] ~^ image[9][6] + signed_kernel[3][0] ~^ image[10][2] + signed_kernel[3][1] ~^ image[10][3] + signed_kernel[3][2] ~^ image[10][4] + signed_kernel[3][3] ~^ image[10][5] + signed_kernel[3][4] ~^ image[10][6] + signed_kernel[4][0] ~^ image[11][2] + signed_kernel[4][1] ~^ image[11][3] + signed_kernel[4][2] ~^ image[11][4] + signed_kernel[4][3] ~^ image[11][5] + signed_kernel[4][4] ~^ image[11][6];
assign xor_sum[7][3] = signed_kernel[0][0] ~^ image[7][3] + signed_kernel[0][1] ~^ image[7][4] + signed_kernel[0][2] ~^ image[7][5] + signed_kernel[0][3] ~^ image[7][6] + signed_kernel[0][4] ~^ image[7][7] + signed_kernel[1][0] ~^ image[8][3] + signed_kernel[1][1] ~^ image[8][4] + signed_kernel[1][2] ~^ image[8][5] + signed_kernel[1][3] ~^ image[8][6] + signed_kernel[1][4] ~^ image[8][7] + signed_kernel[2][0] ~^ image[9][3] + signed_kernel[2][1] ~^ image[9][4] + signed_kernel[2][2] ~^ image[9][5] + signed_kernel[2][3] ~^ image[9][6] + signed_kernel[2][4] ~^ image[9][7] + signed_kernel[3][0] ~^ image[10][3] + signed_kernel[3][1] ~^ image[10][4] + signed_kernel[3][2] ~^ image[10][5] + signed_kernel[3][3] ~^ image[10][6] + signed_kernel[3][4] ~^ image[10][7] + signed_kernel[4][0] ~^ image[11][3] + signed_kernel[4][1] ~^ image[11][4] + signed_kernel[4][2] ~^ image[11][5] + signed_kernel[4][3] ~^ image[11][6] + signed_kernel[4][4] ~^ image[11][7];
assign xor_sum[7][4] = signed_kernel[0][0] ~^ image[7][4] + signed_kernel[0][1] ~^ image[7][5] + signed_kernel[0][2] ~^ image[7][6] + signed_kernel[0][3] ~^ image[7][7] + signed_kernel[0][4] ~^ image[7][8] + signed_kernel[1][0] ~^ image[8][4] + signed_kernel[1][1] ~^ image[8][5] + signed_kernel[1][2] ~^ image[8][6] + signed_kernel[1][3] ~^ image[8][7] + signed_kernel[1][4] ~^ image[8][8] + signed_kernel[2][0] ~^ image[9][4] + signed_kernel[2][1] ~^ image[9][5] + signed_kernel[2][2] ~^ image[9][6] + signed_kernel[2][3] ~^ image[9][7] + signed_kernel[2][4] ~^ image[9][8] + signed_kernel[3][0] ~^ image[10][4] + signed_kernel[3][1] ~^ image[10][5] + signed_kernel[3][2] ~^ image[10][6] + signed_kernel[3][3] ~^ image[10][7] + signed_kernel[3][4] ~^ image[10][8] + signed_kernel[4][0] ~^ image[11][4] + signed_kernel[4][1] ~^ image[11][5] + signed_kernel[4][2] ~^ image[11][6] + signed_kernel[4][3] ~^ image[11][7] + signed_kernel[4][4] ~^ image[11][8];
assign xor_sum[7][5] = signed_kernel[0][0] ~^ image[7][5] + signed_kernel[0][1] ~^ image[7][6] + signed_kernel[0][2] ~^ image[7][7] + signed_kernel[0][3] ~^ image[7][8] + signed_kernel[0][4] ~^ image[7][9] + signed_kernel[1][0] ~^ image[8][5] + signed_kernel[1][1] ~^ image[8][6] + signed_kernel[1][2] ~^ image[8][7] + signed_kernel[1][3] ~^ image[8][8] + signed_kernel[1][4] ~^ image[8][9] + signed_kernel[2][0] ~^ image[9][5] + signed_kernel[2][1] ~^ image[9][6] + signed_kernel[2][2] ~^ image[9][7] + signed_kernel[2][3] ~^ image[9][8] + signed_kernel[2][4] ~^ image[9][9] + signed_kernel[3][0] ~^ image[10][5] + signed_kernel[3][1] ~^ image[10][6] + signed_kernel[3][2] ~^ image[10][7] + signed_kernel[3][3] ~^ image[10][8] + signed_kernel[3][4] ~^ image[10][9] + signed_kernel[4][0] ~^ image[11][5] + signed_kernel[4][1] ~^ image[11][6] + signed_kernel[4][2] ~^ image[11][7] + signed_kernel[4][3] ~^ image[11][8] + signed_kernel[4][4] ~^ image[11][9];
assign xor_sum[7][6] = signed_kernel[0][0] ~^ image[7][6] + signed_kernel[0][1] ~^ image[7][7] + signed_kernel[0][2] ~^ image[7][8] + signed_kernel[0][3] ~^ image[7][9] + signed_kernel[0][4] ~^ image[7][10] + signed_kernel[1][0] ~^ image[8][6] + signed_kernel[1][1] ~^ image[8][7] + signed_kernel[1][2] ~^ image[8][8] + signed_kernel[1][3] ~^ image[8][9] + signed_kernel[1][4] ~^ image[8][10] + signed_kernel[2][0] ~^ image[9][6] + signed_kernel[2][1] ~^ image[9][7] + signed_kernel[2][2] ~^ image[9][8] + signed_kernel[2][3] ~^ image[9][9] + signed_kernel[2][4] ~^ image[9][10] + signed_kernel[3][0] ~^ image[10][6] + signed_kernel[3][1] ~^ image[10][7] + signed_kernel[3][2] ~^ image[10][8] + signed_kernel[3][3] ~^ image[10][9] + signed_kernel[3][4] ~^ image[10][10] + signed_kernel[4][0] ~^ image[11][6] + signed_kernel[4][1] ~^ image[11][7] + signed_kernel[4][2] ~^ image[11][8] + signed_kernel[4][3] ~^ image[11][9] + signed_kernel[4][4] ~^ image[11][10];
assign xor_sum[7][7] = signed_kernel[0][0] ~^ image[7][7] + signed_kernel[0][1] ~^ image[7][8] + signed_kernel[0][2] ~^ image[7][9] + signed_kernel[0][3] ~^ image[7][10] + signed_kernel[0][4] ~^ image[7][11] + signed_kernel[1][0] ~^ image[8][7] + signed_kernel[1][1] ~^ image[8][8] + signed_kernel[1][2] ~^ image[8][9] + signed_kernel[1][3] ~^ image[8][10] + signed_kernel[1][4] ~^ image[8][11] + signed_kernel[2][0] ~^ image[9][7] + signed_kernel[2][1] ~^ image[9][8] + signed_kernel[2][2] ~^ image[9][9] + signed_kernel[2][3] ~^ image[9][10] + signed_kernel[2][4] ~^ image[9][11] + signed_kernel[3][0] ~^ image[10][7] + signed_kernel[3][1] ~^ image[10][8] + signed_kernel[3][2] ~^ image[10][9] + signed_kernel[3][3] ~^ image[10][10] + signed_kernel[3][4] ~^ image[10][11] + signed_kernel[4][0] ~^ image[11][7] + signed_kernel[4][1] ~^ image[11][8] + signed_kernel[4][2] ~^ image[11][9] + signed_kernel[4][3] ~^ image[11][10] + signed_kernel[4][4] ~^ image[11][11];
assign xor_sum[7][8] = signed_kernel[0][0] ~^ image[7][8] + signed_kernel[0][1] ~^ image[7][9] + signed_kernel[0][2] ~^ image[7][10] + signed_kernel[0][3] ~^ image[7][11] + signed_kernel[0][4] ~^ image[7][12] + signed_kernel[1][0] ~^ image[8][8] + signed_kernel[1][1] ~^ image[8][9] + signed_kernel[1][2] ~^ image[8][10] + signed_kernel[1][3] ~^ image[8][11] + signed_kernel[1][4] ~^ image[8][12] + signed_kernel[2][0] ~^ image[9][8] + signed_kernel[2][1] ~^ image[9][9] + signed_kernel[2][2] ~^ image[9][10] + signed_kernel[2][3] ~^ image[9][11] + signed_kernel[2][4] ~^ image[9][12] + signed_kernel[3][0] ~^ image[10][8] + signed_kernel[3][1] ~^ image[10][9] + signed_kernel[3][2] ~^ image[10][10] + signed_kernel[3][3] ~^ image[10][11] + signed_kernel[3][4] ~^ image[10][12] + signed_kernel[4][0] ~^ image[11][8] + signed_kernel[4][1] ~^ image[11][9] + signed_kernel[4][2] ~^ image[11][10] + signed_kernel[4][3] ~^ image[11][11] + signed_kernel[4][4] ~^ image[11][12];
assign xor_sum[7][9] = signed_kernel[0][0] ~^ image[7][9] + signed_kernel[0][1] ~^ image[7][10] + signed_kernel[0][2] ~^ image[7][11] + signed_kernel[0][3] ~^ image[7][12] + signed_kernel[0][4] ~^ image[7][13] + signed_kernel[1][0] ~^ image[8][9] + signed_kernel[1][1] ~^ image[8][10] + signed_kernel[1][2] ~^ image[8][11] + signed_kernel[1][3] ~^ image[8][12] + signed_kernel[1][4] ~^ image[8][13] + signed_kernel[2][0] ~^ image[9][9] + signed_kernel[2][1] ~^ image[9][10] + signed_kernel[2][2] ~^ image[9][11] + signed_kernel[2][3] ~^ image[9][12] + signed_kernel[2][4] ~^ image[9][13] + signed_kernel[3][0] ~^ image[10][9] + signed_kernel[3][1] ~^ image[10][10] + signed_kernel[3][2] ~^ image[10][11] + signed_kernel[3][3] ~^ image[10][12] + signed_kernel[3][4] ~^ image[10][13] + signed_kernel[4][0] ~^ image[11][9] + signed_kernel[4][1] ~^ image[11][10] + signed_kernel[4][2] ~^ image[11][11] + signed_kernel[4][3] ~^ image[11][12] + signed_kernel[4][4] ~^ image[11][13];
assign xor_sum[7][10] = signed_kernel[0][0] ~^ image[7][10] + signed_kernel[0][1] ~^ image[7][11] + signed_kernel[0][2] ~^ image[7][12] + signed_kernel[0][3] ~^ image[7][13] + signed_kernel[0][4] ~^ image[7][14] + signed_kernel[1][0] ~^ image[8][10] + signed_kernel[1][1] ~^ image[8][11] + signed_kernel[1][2] ~^ image[8][12] + signed_kernel[1][3] ~^ image[8][13] + signed_kernel[1][4] ~^ image[8][14] + signed_kernel[2][0] ~^ image[9][10] + signed_kernel[2][1] ~^ image[9][11] + signed_kernel[2][2] ~^ image[9][12] + signed_kernel[2][3] ~^ image[9][13] + signed_kernel[2][4] ~^ image[9][14] + signed_kernel[3][0] ~^ image[10][10] + signed_kernel[3][1] ~^ image[10][11] + signed_kernel[3][2] ~^ image[10][12] + signed_kernel[3][3] ~^ image[10][13] + signed_kernel[3][4] ~^ image[10][14] + signed_kernel[4][0] ~^ image[11][10] + signed_kernel[4][1] ~^ image[11][11] + signed_kernel[4][2] ~^ image[11][12] + signed_kernel[4][3] ~^ image[11][13] + signed_kernel[4][4] ~^ image[11][14];
assign xor_sum[7][11] = signed_kernel[0][0] ~^ image[7][11] + signed_kernel[0][1] ~^ image[7][12] + signed_kernel[0][2] ~^ image[7][13] + signed_kernel[0][3] ~^ image[7][14] + signed_kernel[0][4] ~^ image[7][15] + signed_kernel[1][0] ~^ image[8][11] + signed_kernel[1][1] ~^ image[8][12] + signed_kernel[1][2] ~^ image[8][13] + signed_kernel[1][3] ~^ image[8][14] + signed_kernel[1][4] ~^ image[8][15] + signed_kernel[2][0] ~^ image[9][11] + signed_kernel[2][1] ~^ image[9][12] + signed_kernel[2][2] ~^ image[9][13] + signed_kernel[2][3] ~^ image[9][14] + signed_kernel[2][4] ~^ image[9][15] + signed_kernel[3][0] ~^ image[10][11] + signed_kernel[3][1] ~^ image[10][12] + signed_kernel[3][2] ~^ image[10][13] + signed_kernel[3][3] ~^ image[10][14] + signed_kernel[3][4] ~^ image[10][15] + signed_kernel[4][0] ~^ image[11][11] + signed_kernel[4][1] ~^ image[11][12] + signed_kernel[4][2] ~^ image[11][13] + signed_kernel[4][3] ~^ image[11][14] + signed_kernel[4][4] ~^ image[11][15];
assign xor_sum[7][12] = signed_kernel[0][0] ~^ image[7][12] + signed_kernel[0][1] ~^ image[7][13] + signed_kernel[0][2] ~^ image[7][14] + signed_kernel[0][3] ~^ image[7][15] + signed_kernel[0][4] ~^ image[7][16] + signed_kernel[1][0] ~^ image[8][12] + signed_kernel[1][1] ~^ image[8][13] + signed_kernel[1][2] ~^ image[8][14] + signed_kernel[1][3] ~^ image[8][15] + signed_kernel[1][4] ~^ image[8][16] + signed_kernel[2][0] ~^ image[9][12] + signed_kernel[2][1] ~^ image[9][13] + signed_kernel[2][2] ~^ image[9][14] + signed_kernel[2][3] ~^ image[9][15] + signed_kernel[2][4] ~^ image[9][16] + signed_kernel[3][0] ~^ image[10][12] + signed_kernel[3][1] ~^ image[10][13] + signed_kernel[3][2] ~^ image[10][14] + signed_kernel[3][3] ~^ image[10][15] + signed_kernel[3][4] ~^ image[10][16] + signed_kernel[4][0] ~^ image[11][12] + signed_kernel[4][1] ~^ image[11][13] + signed_kernel[4][2] ~^ image[11][14] + signed_kernel[4][3] ~^ image[11][15] + signed_kernel[4][4] ~^ image[11][16];
assign xor_sum[7][13] = signed_kernel[0][0] ~^ image[7][13] + signed_kernel[0][1] ~^ image[7][14] + signed_kernel[0][2] ~^ image[7][15] + signed_kernel[0][3] ~^ image[7][16] + signed_kernel[0][4] ~^ image[7][17] + signed_kernel[1][0] ~^ image[8][13] + signed_kernel[1][1] ~^ image[8][14] + signed_kernel[1][2] ~^ image[8][15] + signed_kernel[1][3] ~^ image[8][16] + signed_kernel[1][4] ~^ image[8][17] + signed_kernel[2][0] ~^ image[9][13] + signed_kernel[2][1] ~^ image[9][14] + signed_kernel[2][2] ~^ image[9][15] + signed_kernel[2][3] ~^ image[9][16] + signed_kernel[2][4] ~^ image[9][17] + signed_kernel[3][0] ~^ image[10][13] + signed_kernel[3][1] ~^ image[10][14] + signed_kernel[3][2] ~^ image[10][15] + signed_kernel[3][3] ~^ image[10][16] + signed_kernel[3][4] ~^ image[10][17] + signed_kernel[4][0] ~^ image[11][13] + signed_kernel[4][1] ~^ image[11][14] + signed_kernel[4][2] ~^ image[11][15] + signed_kernel[4][3] ~^ image[11][16] + signed_kernel[4][4] ~^ image[11][17];
assign xor_sum[7][14] = signed_kernel[0][0] ~^ image[7][14] + signed_kernel[0][1] ~^ image[7][15] + signed_kernel[0][2] ~^ image[7][16] + signed_kernel[0][3] ~^ image[7][17] + signed_kernel[0][4] ~^ image[7][18] + signed_kernel[1][0] ~^ image[8][14] + signed_kernel[1][1] ~^ image[8][15] + signed_kernel[1][2] ~^ image[8][16] + signed_kernel[1][3] ~^ image[8][17] + signed_kernel[1][4] ~^ image[8][18] + signed_kernel[2][0] ~^ image[9][14] + signed_kernel[2][1] ~^ image[9][15] + signed_kernel[2][2] ~^ image[9][16] + signed_kernel[2][3] ~^ image[9][17] + signed_kernel[2][4] ~^ image[9][18] + signed_kernel[3][0] ~^ image[10][14] + signed_kernel[3][1] ~^ image[10][15] + signed_kernel[3][2] ~^ image[10][16] + signed_kernel[3][3] ~^ image[10][17] + signed_kernel[3][4] ~^ image[10][18] + signed_kernel[4][0] ~^ image[11][14] + signed_kernel[4][1] ~^ image[11][15] + signed_kernel[4][2] ~^ image[11][16] + signed_kernel[4][3] ~^ image[11][17] + signed_kernel[4][4] ~^ image[11][18];
assign xor_sum[7][15] = signed_kernel[0][0] ~^ image[7][15] + signed_kernel[0][1] ~^ image[7][16] + signed_kernel[0][2] ~^ image[7][17] + signed_kernel[0][3] ~^ image[7][18] + signed_kernel[0][4] ~^ image[7][19] + signed_kernel[1][0] ~^ image[8][15] + signed_kernel[1][1] ~^ image[8][16] + signed_kernel[1][2] ~^ image[8][17] + signed_kernel[1][3] ~^ image[8][18] + signed_kernel[1][4] ~^ image[8][19] + signed_kernel[2][0] ~^ image[9][15] + signed_kernel[2][1] ~^ image[9][16] + signed_kernel[2][2] ~^ image[9][17] + signed_kernel[2][3] ~^ image[9][18] + signed_kernel[2][4] ~^ image[9][19] + signed_kernel[3][0] ~^ image[10][15] + signed_kernel[3][1] ~^ image[10][16] + signed_kernel[3][2] ~^ image[10][17] + signed_kernel[3][3] ~^ image[10][18] + signed_kernel[3][4] ~^ image[10][19] + signed_kernel[4][0] ~^ image[11][15] + signed_kernel[4][1] ~^ image[11][16] + signed_kernel[4][2] ~^ image[11][17] + signed_kernel[4][3] ~^ image[11][18] + signed_kernel[4][4] ~^ image[11][19];
assign xor_sum[7][16] = signed_kernel[0][0] ~^ image[7][16] + signed_kernel[0][1] ~^ image[7][17] + signed_kernel[0][2] ~^ image[7][18] + signed_kernel[0][3] ~^ image[7][19] + signed_kernel[0][4] ~^ image[7][20] + signed_kernel[1][0] ~^ image[8][16] + signed_kernel[1][1] ~^ image[8][17] + signed_kernel[1][2] ~^ image[8][18] + signed_kernel[1][3] ~^ image[8][19] + signed_kernel[1][4] ~^ image[8][20] + signed_kernel[2][0] ~^ image[9][16] + signed_kernel[2][1] ~^ image[9][17] + signed_kernel[2][2] ~^ image[9][18] + signed_kernel[2][3] ~^ image[9][19] + signed_kernel[2][4] ~^ image[9][20] + signed_kernel[3][0] ~^ image[10][16] + signed_kernel[3][1] ~^ image[10][17] + signed_kernel[3][2] ~^ image[10][18] + signed_kernel[3][3] ~^ image[10][19] + signed_kernel[3][4] ~^ image[10][20] + signed_kernel[4][0] ~^ image[11][16] + signed_kernel[4][1] ~^ image[11][17] + signed_kernel[4][2] ~^ image[11][18] + signed_kernel[4][3] ~^ image[11][19] + signed_kernel[4][4] ~^ image[11][20];
assign xor_sum[7][17] = signed_kernel[0][0] ~^ image[7][17] + signed_kernel[0][1] ~^ image[7][18] + signed_kernel[0][2] ~^ image[7][19] + signed_kernel[0][3] ~^ image[7][20] + signed_kernel[0][4] ~^ image[7][21] + signed_kernel[1][0] ~^ image[8][17] + signed_kernel[1][1] ~^ image[8][18] + signed_kernel[1][2] ~^ image[8][19] + signed_kernel[1][3] ~^ image[8][20] + signed_kernel[1][4] ~^ image[8][21] + signed_kernel[2][0] ~^ image[9][17] + signed_kernel[2][1] ~^ image[9][18] + signed_kernel[2][2] ~^ image[9][19] + signed_kernel[2][3] ~^ image[9][20] + signed_kernel[2][4] ~^ image[9][21] + signed_kernel[3][0] ~^ image[10][17] + signed_kernel[3][1] ~^ image[10][18] + signed_kernel[3][2] ~^ image[10][19] + signed_kernel[3][3] ~^ image[10][20] + signed_kernel[3][4] ~^ image[10][21] + signed_kernel[4][0] ~^ image[11][17] + signed_kernel[4][1] ~^ image[11][18] + signed_kernel[4][2] ~^ image[11][19] + signed_kernel[4][3] ~^ image[11][20] + signed_kernel[4][4] ~^ image[11][21];
assign xor_sum[7][18] = signed_kernel[0][0] ~^ image[7][18] + signed_kernel[0][1] ~^ image[7][19] + signed_kernel[0][2] ~^ image[7][20] + signed_kernel[0][3] ~^ image[7][21] + signed_kernel[0][4] ~^ image[7][22] + signed_kernel[1][0] ~^ image[8][18] + signed_kernel[1][1] ~^ image[8][19] + signed_kernel[1][2] ~^ image[8][20] + signed_kernel[1][3] ~^ image[8][21] + signed_kernel[1][4] ~^ image[8][22] + signed_kernel[2][0] ~^ image[9][18] + signed_kernel[2][1] ~^ image[9][19] + signed_kernel[2][2] ~^ image[9][20] + signed_kernel[2][3] ~^ image[9][21] + signed_kernel[2][4] ~^ image[9][22] + signed_kernel[3][0] ~^ image[10][18] + signed_kernel[3][1] ~^ image[10][19] + signed_kernel[3][2] ~^ image[10][20] + signed_kernel[3][3] ~^ image[10][21] + signed_kernel[3][4] ~^ image[10][22] + signed_kernel[4][0] ~^ image[11][18] + signed_kernel[4][1] ~^ image[11][19] + signed_kernel[4][2] ~^ image[11][20] + signed_kernel[4][3] ~^ image[11][21] + signed_kernel[4][4] ~^ image[11][22];
assign xor_sum[7][19] = signed_kernel[0][0] ~^ image[7][19] + signed_kernel[0][1] ~^ image[7][20] + signed_kernel[0][2] ~^ image[7][21] + signed_kernel[0][3] ~^ image[7][22] + signed_kernel[0][4] ~^ image[7][23] + signed_kernel[1][0] ~^ image[8][19] + signed_kernel[1][1] ~^ image[8][20] + signed_kernel[1][2] ~^ image[8][21] + signed_kernel[1][3] ~^ image[8][22] + signed_kernel[1][4] ~^ image[8][23] + signed_kernel[2][0] ~^ image[9][19] + signed_kernel[2][1] ~^ image[9][20] + signed_kernel[2][2] ~^ image[9][21] + signed_kernel[2][3] ~^ image[9][22] + signed_kernel[2][4] ~^ image[9][23] + signed_kernel[3][0] ~^ image[10][19] + signed_kernel[3][1] ~^ image[10][20] + signed_kernel[3][2] ~^ image[10][21] + signed_kernel[3][3] ~^ image[10][22] + signed_kernel[3][4] ~^ image[10][23] + signed_kernel[4][0] ~^ image[11][19] + signed_kernel[4][1] ~^ image[11][20] + signed_kernel[4][2] ~^ image[11][21] + signed_kernel[4][3] ~^ image[11][22] + signed_kernel[4][4] ~^ image[11][23];
assign xor_sum[7][20] = signed_kernel[0][0] ~^ image[7][20] + signed_kernel[0][1] ~^ image[7][21] + signed_kernel[0][2] ~^ image[7][22] + signed_kernel[0][3] ~^ image[7][23] + signed_kernel[0][4] ~^ image[7][24] + signed_kernel[1][0] ~^ image[8][20] + signed_kernel[1][1] ~^ image[8][21] + signed_kernel[1][2] ~^ image[8][22] + signed_kernel[1][3] ~^ image[8][23] + signed_kernel[1][4] ~^ image[8][24] + signed_kernel[2][0] ~^ image[9][20] + signed_kernel[2][1] ~^ image[9][21] + signed_kernel[2][2] ~^ image[9][22] + signed_kernel[2][3] ~^ image[9][23] + signed_kernel[2][4] ~^ image[9][24] + signed_kernel[3][0] ~^ image[10][20] + signed_kernel[3][1] ~^ image[10][21] + signed_kernel[3][2] ~^ image[10][22] + signed_kernel[3][3] ~^ image[10][23] + signed_kernel[3][4] ~^ image[10][24] + signed_kernel[4][0] ~^ image[11][20] + signed_kernel[4][1] ~^ image[11][21] + signed_kernel[4][2] ~^ image[11][22] + signed_kernel[4][3] ~^ image[11][23] + signed_kernel[4][4] ~^ image[11][24];
assign xor_sum[7][21] = signed_kernel[0][0] ~^ image[7][21] + signed_kernel[0][1] ~^ image[7][22] + signed_kernel[0][2] ~^ image[7][23] + signed_kernel[0][3] ~^ image[7][24] + signed_kernel[0][4] ~^ image[7][25] + signed_kernel[1][0] ~^ image[8][21] + signed_kernel[1][1] ~^ image[8][22] + signed_kernel[1][2] ~^ image[8][23] + signed_kernel[1][3] ~^ image[8][24] + signed_kernel[1][4] ~^ image[8][25] + signed_kernel[2][0] ~^ image[9][21] + signed_kernel[2][1] ~^ image[9][22] + signed_kernel[2][2] ~^ image[9][23] + signed_kernel[2][3] ~^ image[9][24] + signed_kernel[2][4] ~^ image[9][25] + signed_kernel[3][0] ~^ image[10][21] + signed_kernel[3][1] ~^ image[10][22] + signed_kernel[3][2] ~^ image[10][23] + signed_kernel[3][3] ~^ image[10][24] + signed_kernel[3][4] ~^ image[10][25] + signed_kernel[4][0] ~^ image[11][21] + signed_kernel[4][1] ~^ image[11][22] + signed_kernel[4][2] ~^ image[11][23] + signed_kernel[4][3] ~^ image[11][24] + signed_kernel[4][4] ~^ image[11][25];
assign xor_sum[7][22] = signed_kernel[0][0] ~^ image[7][22] + signed_kernel[0][1] ~^ image[7][23] + signed_kernel[0][2] ~^ image[7][24] + signed_kernel[0][3] ~^ image[7][25] + signed_kernel[0][4] ~^ image[7][26] + signed_kernel[1][0] ~^ image[8][22] + signed_kernel[1][1] ~^ image[8][23] + signed_kernel[1][2] ~^ image[8][24] + signed_kernel[1][3] ~^ image[8][25] + signed_kernel[1][4] ~^ image[8][26] + signed_kernel[2][0] ~^ image[9][22] + signed_kernel[2][1] ~^ image[9][23] + signed_kernel[2][2] ~^ image[9][24] + signed_kernel[2][3] ~^ image[9][25] + signed_kernel[2][4] ~^ image[9][26] + signed_kernel[3][0] ~^ image[10][22] + signed_kernel[3][1] ~^ image[10][23] + signed_kernel[3][2] ~^ image[10][24] + signed_kernel[3][3] ~^ image[10][25] + signed_kernel[3][4] ~^ image[10][26] + signed_kernel[4][0] ~^ image[11][22] + signed_kernel[4][1] ~^ image[11][23] + signed_kernel[4][2] ~^ image[11][24] + signed_kernel[4][3] ~^ image[11][25] + signed_kernel[4][4] ~^ image[11][26];
assign xor_sum[7][23] = signed_kernel[0][0] ~^ image[7][23] + signed_kernel[0][1] ~^ image[7][24] + signed_kernel[0][2] ~^ image[7][25] + signed_kernel[0][3] ~^ image[7][26] + signed_kernel[0][4] ~^ image[7][27] + signed_kernel[1][0] ~^ image[8][23] + signed_kernel[1][1] ~^ image[8][24] + signed_kernel[1][2] ~^ image[8][25] + signed_kernel[1][3] ~^ image[8][26] + signed_kernel[1][4] ~^ image[8][27] + signed_kernel[2][0] ~^ image[9][23] + signed_kernel[2][1] ~^ image[9][24] + signed_kernel[2][2] ~^ image[9][25] + signed_kernel[2][3] ~^ image[9][26] + signed_kernel[2][4] ~^ image[9][27] + signed_kernel[3][0] ~^ image[10][23] + signed_kernel[3][1] ~^ image[10][24] + signed_kernel[3][2] ~^ image[10][25] + signed_kernel[3][3] ~^ image[10][26] + signed_kernel[3][4] ~^ image[10][27] + signed_kernel[4][0] ~^ image[11][23] + signed_kernel[4][1] ~^ image[11][24] + signed_kernel[4][2] ~^ image[11][25] + signed_kernel[4][3] ~^ image[11][26] + signed_kernel[4][4] ~^ image[11][27];
assign xor_sum[8][0] = signed_kernel[0][0] ~^ image[8][0] + signed_kernel[0][1] ~^ image[8][1] + signed_kernel[0][2] ~^ image[8][2] + signed_kernel[0][3] ~^ image[8][3] + signed_kernel[0][4] ~^ image[8][4] + signed_kernel[1][0] ~^ image[9][0] + signed_kernel[1][1] ~^ image[9][1] + signed_kernel[1][2] ~^ image[9][2] + signed_kernel[1][3] ~^ image[9][3] + signed_kernel[1][4] ~^ image[9][4] + signed_kernel[2][0] ~^ image[10][0] + signed_kernel[2][1] ~^ image[10][1] + signed_kernel[2][2] ~^ image[10][2] + signed_kernel[2][3] ~^ image[10][3] + signed_kernel[2][4] ~^ image[10][4] + signed_kernel[3][0] ~^ image[11][0] + signed_kernel[3][1] ~^ image[11][1] + signed_kernel[3][2] ~^ image[11][2] + signed_kernel[3][3] ~^ image[11][3] + signed_kernel[3][4] ~^ image[11][4] + signed_kernel[4][0] ~^ image[12][0] + signed_kernel[4][1] ~^ image[12][1] + signed_kernel[4][2] ~^ image[12][2] + signed_kernel[4][3] ~^ image[12][3] + signed_kernel[4][4] ~^ image[12][4];
assign xor_sum[8][1] = signed_kernel[0][0] ~^ image[8][1] + signed_kernel[0][1] ~^ image[8][2] + signed_kernel[0][2] ~^ image[8][3] + signed_kernel[0][3] ~^ image[8][4] + signed_kernel[0][4] ~^ image[8][5] + signed_kernel[1][0] ~^ image[9][1] + signed_kernel[1][1] ~^ image[9][2] + signed_kernel[1][2] ~^ image[9][3] + signed_kernel[1][3] ~^ image[9][4] + signed_kernel[1][4] ~^ image[9][5] + signed_kernel[2][0] ~^ image[10][1] + signed_kernel[2][1] ~^ image[10][2] + signed_kernel[2][2] ~^ image[10][3] + signed_kernel[2][3] ~^ image[10][4] + signed_kernel[2][4] ~^ image[10][5] + signed_kernel[3][0] ~^ image[11][1] + signed_kernel[3][1] ~^ image[11][2] + signed_kernel[3][2] ~^ image[11][3] + signed_kernel[3][3] ~^ image[11][4] + signed_kernel[3][4] ~^ image[11][5] + signed_kernel[4][0] ~^ image[12][1] + signed_kernel[4][1] ~^ image[12][2] + signed_kernel[4][2] ~^ image[12][3] + signed_kernel[4][3] ~^ image[12][4] + signed_kernel[4][4] ~^ image[12][5];
assign xor_sum[8][2] = signed_kernel[0][0] ~^ image[8][2] + signed_kernel[0][1] ~^ image[8][3] + signed_kernel[0][2] ~^ image[8][4] + signed_kernel[0][3] ~^ image[8][5] + signed_kernel[0][4] ~^ image[8][6] + signed_kernel[1][0] ~^ image[9][2] + signed_kernel[1][1] ~^ image[9][3] + signed_kernel[1][2] ~^ image[9][4] + signed_kernel[1][3] ~^ image[9][5] + signed_kernel[1][4] ~^ image[9][6] + signed_kernel[2][0] ~^ image[10][2] + signed_kernel[2][1] ~^ image[10][3] + signed_kernel[2][2] ~^ image[10][4] + signed_kernel[2][3] ~^ image[10][5] + signed_kernel[2][4] ~^ image[10][6] + signed_kernel[3][0] ~^ image[11][2] + signed_kernel[3][1] ~^ image[11][3] + signed_kernel[3][2] ~^ image[11][4] + signed_kernel[3][3] ~^ image[11][5] + signed_kernel[3][4] ~^ image[11][6] + signed_kernel[4][0] ~^ image[12][2] + signed_kernel[4][1] ~^ image[12][3] + signed_kernel[4][2] ~^ image[12][4] + signed_kernel[4][3] ~^ image[12][5] + signed_kernel[4][4] ~^ image[12][6];
assign xor_sum[8][3] = signed_kernel[0][0] ~^ image[8][3] + signed_kernel[0][1] ~^ image[8][4] + signed_kernel[0][2] ~^ image[8][5] + signed_kernel[0][3] ~^ image[8][6] + signed_kernel[0][4] ~^ image[8][7] + signed_kernel[1][0] ~^ image[9][3] + signed_kernel[1][1] ~^ image[9][4] + signed_kernel[1][2] ~^ image[9][5] + signed_kernel[1][3] ~^ image[9][6] + signed_kernel[1][4] ~^ image[9][7] + signed_kernel[2][0] ~^ image[10][3] + signed_kernel[2][1] ~^ image[10][4] + signed_kernel[2][2] ~^ image[10][5] + signed_kernel[2][3] ~^ image[10][6] + signed_kernel[2][4] ~^ image[10][7] + signed_kernel[3][0] ~^ image[11][3] + signed_kernel[3][1] ~^ image[11][4] + signed_kernel[3][2] ~^ image[11][5] + signed_kernel[3][3] ~^ image[11][6] + signed_kernel[3][4] ~^ image[11][7] + signed_kernel[4][0] ~^ image[12][3] + signed_kernel[4][1] ~^ image[12][4] + signed_kernel[4][2] ~^ image[12][5] + signed_kernel[4][3] ~^ image[12][6] + signed_kernel[4][4] ~^ image[12][7];
assign xor_sum[8][4] = signed_kernel[0][0] ~^ image[8][4] + signed_kernel[0][1] ~^ image[8][5] + signed_kernel[0][2] ~^ image[8][6] + signed_kernel[0][3] ~^ image[8][7] + signed_kernel[0][4] ~^ image[8][8] + signed_kernel[1][0] ~^ image[9][4] + signed_kernel[1][1] ~^ image[9][5] + signed_kernel[1][2] ~^ image[9][6] + signed_kernel[1][3] ~^ image[9][7] + signed_kernel[1][4] ~^ image[9][8] + signed_kernel[2][0] ~^ image[10][4] + signed_kernel[2][1] ~^ image[10][5] + signed_kernel[2][2] ~^ image[10][6] + signed_kernel[2][3] ~^ image[10][7] + signed_kernel[2][4] ~^ image[10][8] + signed_kernel[3][0] ~^ image[11][4] + signed_kernel[3][1] ~^ image[11][5] + signed_kernel[3][2] ~^ image[11][6] + signed_kernel[3][3] ~^ image[11][7] + signed_kernel[3][4] ~^ image[11][8] + signed_kernel[4][0] ~^ image[12][4] + signed_kernel[4][1] ~^ image[12][5] + signed_kernel[4][2] ~^ image[12][6] + signed_kernel[4][3] ~^ image[12][7] + signed_kernel[4][4] ~^ image[12][8];
assign xor_sum[8][5] = signed_kernel[0][0] ~^ image[8][5] + signed_kernel[0][1] ~^ image[8][6] + signed_kernel[0][2] ~^ image[8][7] + signed_kernel[0][3] ~^ image[8][8] + signed_kernel[0][4] ~^ image[8][9] + signed_kernel[1][0] ~^ image[9][5] + signed_kernel[1][1] ~^ image[9][6] + signed_kernel[1][2] ~^ image[9][7] + signed_kernel[1][3] ~^ image[9][8] + signed_kernel[1][4] ~^ image[9][9] + signed_kernel[2][0] ~^ image[10][5] + signed_kernel[2][1] ~^ image[10][6] + signed_kernel[2][2] ~^ image[10][7] + signed_kernel[2][3] ~^ image[10][8] + signed_kernel[2][4] ~^ image[10][9] + signed_kernel[3][0] ~^ image[11][5] + signed_kernel[3][1] ~^ image[11][6] + signed_kernel[3][2] ~^ image[11][7] + signed_kernel[3][3] ~^ image[11][8] + signed_kernel[3][4] ~^ image[11][9] + signed_kernel[4][0] ~^ image[12][5] + signed_kernel[4][1] ~^ image[12][6] + signed_kernel[4][2] ~^ image[12][7] + signed_kernel[4][3] ~^ image[12][8] + signed_kernel[4][4] ~^ image[12][9];
assign xor_sum[8][6] = signed_kernel[0][0] ~^ image[8][6] + signed_kernel[0][1] ~^ image[8][7] + signed_kernel[0][2] ~^ image[8][8] + signed_kernel[0][3] ~^ image[8][9] + signed_kernel[0][4] ~^ image[8][10] + signed_kernel[1][0] ~^ image[9][6] + signed_kernel[1][1] ~^ image[9][7] + signed_kernel[1][2] ~^ image[9][8] + signed_kernel[1][3] ~^ image[9][9] + signed_kernel[1][4] ~^ image[9][10] + signed_kernel[2][0] ~^ image[10][6] + signed_kernel[2][1] ~^ image[10][7] + signed_kernel[2][2] ~^ image[10][8] + signed_kernel[2][3] ~^ image[10][9] + signed_kernel[2][4] ~^ image[10][10] + signed_kernel[3][0] ~^ image[11][6] + signed_kernel[3][1] ~^ image[11][7] + signed_kernel[3][2] ~^ image[11][8] + signed_kernel[3][3] ~^ image[11][9] + signed_kernel[3][4] ~^ image[11][10] + signed_kernel[4][0] ~^ image[12][6] + signed_kernel[4][1] ~^ image[12][7] + signed_kernel[4][2] ~^ image[12][8] + signed_kernel[4][3] ~^ image[12][9] + signed_kernel[4][4] ~^ image[12][10];
assign xor_sum[8][7] = signed_kernel[0][0] ~^ image[8][7] + signed_kernel[0][1] ~^ image[8][8] + signed_kernel[0][2] ~^ image[8][9] + signed_kernel[0][3] ~^ image[8][10] + signed_kernel[0][4] ~^ image[8][11] + signed_kernel[1][0] ~^ image[9][7] + signed_kernel[1][1] ~^ image[9][8] + signed_kernel[1][2] ~^ image[9][9] + signed_kernel[1][3] ~^ image[9][10] + signed_kernel[1][4] ~^ image[9][11] + signed_kernel[2][0] ~^ image[10][7] + signed_kernel[2][1] ~^ image[10][8] + signed_kernel[2][2] ~^ image[10][9] + signed_kernel[2][3] ~^ image[10][10] + signed_kernel[2][4] ~^ image[10][11] + signed_kernel[3][0] ~^ image[11][7] + signed_kernel[3][1] ~^ image[11][8] + signed_kernel[3][2] ~^ image[11][9] + signed_kernel[3][3] ~^ image[11][10] + signed_kernel[3][4] ~^ image[11][11] + signed_kernel[4][0] ~^ image[12][7] + signed_kernel[4][1] ~^ image[12][8] + signed_kernel[4][2] ~^ image[12][9] + signed_kernel[4][3] ~^ image[12][10] + signed_kernel[4][4] ~^ image[12][11];
assign xor_sum[8][8] = signed_kernel[0][0] ~^ image[8][8] + signed_kernel[0][1] ~^ image[8][9] + signed_kernel[0][2] ~^ image[8][10] + signed_kernel[0][3] ~^ image[8][11] + signed_kernel[0][4] ~^ image[8][12] + signed_kernel[1][0] ~^ image[9][8] + signed_kernel[1][1] ~^ image[9][9] + signed_kernel[1][2] ~^ image[9][10] + signed_kernel[1][3] ~^ image[9][11] + signed_kernel[1][4] ~^ image[9][12] + signed_kernel[2][0] ~^ image[10][8] + signed_kernel[2][1] ~^ image[10][9] + signed_kernel[2][2] ~^ image[10][10] + signed_kernel[2][3] ~^ image[10][11] + signed_kernel[2][4] ~^ image[10][12] + signed_kernel[3][0] ~^ image[11][8] + signed_kernel[3][1] ~^ image[11][9] + signed_kernel[3][2] ~^ image[11][10] + signed_kernel[3][3] ~^ image[11][11] + signed_kernel[3][4] ~^ image[11][12] + signed_kernel[4][0] ~^ image[12][8] + signed_kernel[4][1] ~^ image[12][9] + signed_kernel[4][2] ~^ image[12][10] + signed_kernel[4][3] ~^ image[12][11] + signed_kernel[4][4] ~^ image[12][12];
assign xor_sum[8][9] = signed_kernel[0][0] ~^ image[8][9] + signed_kernel[0][1] ~^ image[8][10] + signed_kernel[0][2] ~^ image[8][11] + signed_kernel[0][3] ~^ image[8][12] + signed_kernel[0][4] ~^ image[8][13] + signed_kernel[1][0] ~^ image[9][9] + signed_kernel[1][1] ~^ image[9][10] + signed_kernel[1][2] ~^ image[9][11] + signed_kernel[1][3] ~^ image[9][12] + signed_kernel[1][4] ~^ image[9][13] + signed_kernel[2][0] ~^ image[10][9] + signed_kernel[2][1] ~^ image[10][10] + signed_kernel[2][2] ~^ image[10][11] + signed_kernel[2][3] ~^ image[10][12] + signed_kernel[2][4] ~^ image[10][13] + signed_kernel[3][0] ~^ image[11][9] + signed_kernel[3][1] ~^ image[11][10] + signed_kernel[3][2] ~^ image[11][11] + signed_kernel[3][3] ~^ image[11][12] + signed_kernel[3][4] ~^ image[11][13] + signed_kernel[4][0] ~^ image[12][9] + signed_kernel[4][1] ~^ image[12][10] + signed_kernel[4][2] ~^ image[12][11] + signed_kernel[4][3] ~^ image[12][12] + signed_kernel[4][4] ~^ image[12][13];
assign xor_sum[8][10] = signed_kernel[0][0] ~^ image[8][10] + signed_kernel[0][1] ~^ image[8][11] + signed_kernel[0][2] ~^ image[8][12] + signed_kernel[0][3] ~^ image[8][13] + signed_kernel[0][4] ~^ image[8][14] + signed_kernel[1][0] ~^ image[9][10] + signed_kernel[1][1] ~^ image[9][11] + signed_kernel[1][2] ~^ image[9][12] + signed_kernel[1][3] ~^ image[9][13] + signed_kernel[1][4] ~^ image[9][14] + signed_kernel[2][0] ~^ image[10][10] + signed_kernel[2][1] ~^ image[10][11] + signed_kernel[2][2] ~^ image[10][12] + signed_kernel[2][3] ~^ image[10][13] + signed_kernel[2][4] ~^ image[10][14] + signed_kernel[3][0] ~^ image[11][10] + signed_kernel[3][1] ~^ image[11][11] + signed_kernel[3][2] ~^ image[11][12] + signed_kernel[3][3] ~^ image[11][13] + signed_kernel[3][4] ~^ image[11][14] + signed_kernel[4][0] ~^ image[12][10] + signed_kernel[4][1] ~^ image[12][11] + signed_kernel[4][2] ~^ image[12][12] + signed_kernel[4][3] ~^ image[12][13] + signed_kernel[4][4] ~^ image[12][14];
assign xor_sum[8][11] = signed_kernel[0][0] ~^ image[8][11] + signed_kernel[0][1] ~^ image[8][12] + signed_kernel[0][2] ~^ image[8][13] + signed_kernel[0][3] ~^ image[8][14] + signed_kernel[0][4] ~^ image[8][15] + signed_kernel[1][0] ~^ image[9][11] + signed_kernel[1][1] ~^ image[9][12] + signed_kernel[1][2] ~^ image[9][13] + signed_kernel[1][3] ~^ image[9][14] + signed_kernel[1][4] ~^ image[9][15] + signed_kernel[2][0] ~^ image[10][11] + signed_kernel[2][1] ~^ image[10][12] + signed_kernel[2][2] ~^ image[10][13] + signed_kernel[2][3] ~^ image[10][14] + signed_kernel[2][4] ~^ image[10][15] + signed_kernel[3][0] ~^ image[11][11] + signed_kernel[3][1] ~^ image[11][12] + signed_kernel[3][2] ~^ image[11][13] + signed_kernel[3][3] ~^ image[11][14] + signed_kernel[3][4] ~^ image[11][15] + signed_kernel[4][0] ~^ image[12][11] + signed_kernel[4][1] ~^ image[12][12] + signed_kernel[4][2] ~^ image[12][13] + signed_kernel[4][3] ~^ image[12][14] + signed_kernel[4][4] ~^ image[12][15];
assign xor_sum[8][12] = signed_kernel[0][0] ~^ image[8][12] + signed_kernel[0][1] ~^ image[8][13] + signed_kernel[0][2] ~^ image[8][14] + signed_kernel[0][3] ~^ image[8][15] + signed_kernel[0][4] ~^ image[8][16] + signed_kernel[1][0] ~^ image[9][12] + signed_kernel[1][1] ~^ image[9][13] + signed_kernel[1][2] ~^ image[9][14] + signed_kernel[1][3] ~^ image[9][15] + signed_kernel[1][4] ~^ image[9][16] + signed_kernel[2][0] ~^ image[10][12] + signed_kernel[2][1] ~^ image[10][13] + signed_kernel[2][2] ~^ image[10][14] + signed_kernel[2][3] ~^ image[10][15] + signed_kernel[2][4] ~^ image[10][16] + signed_kernel[3][0] ~^ image[11][12] + signed_kernel[3][1] ~^ image[11][13] + signed_kernel[3][2] ~^ image[11][14] + signed_kernel[3][3] ~^ image[11][15] + signed_kernel[3][4] ~^ image[11][16] + signed_kernel[4][0] ~^ image[12][12] + signed_kernel[4][1] ~^ image[12][13] + signed_kernel[4][2] ~^ image[12][14] + signed_kernel[4][3] ~^ image[12][15] + signed_kernel[4][4] ~^ image[12][16];
assign xor_sum[8][13] = signed_kernel[0][0] ~^ image[8][13] + signed_kernel[0][1] ~^ image[8][14] + signed_kernel[0][2] ~^ image[8][15] + signed_kernel[0][3] ~^ image[8][16] + signed_kernel[0][4] ~^ image[8][17] + signed_kernel[1][0] ~^ image[9][13] + signed_kernel[1][1] ~^ image[9][14] + signed_kernel[1][2] ~^ image[9][15] + signed_kernel[1][3] ~^ image[9][16] + signed_kernel[1][4] ~^ image[9][17] + signed_kernel[2][0] ~^ image[10][13] + signed_kernel[2][1] ~^ image[10][14] + signed_kernel[2][2] ~^ image[10][15] + signed_kernel[2][3] ~^ image[10][16] + signed_kernel[2][4] ~^ image[10][17] + signed_kernel[3][0] ~^ image[11][13] + signed_kernel[3][1] ~^ image[11][14] + signed_kernel[3][2] ~^ image[11][15] + signed_kernel[3][3] ~^ image[11][16] + signed_kernel[3][4] ~^ image[11][17] + signed_kernel[4][0] ~^ image[12][13] + signed_kernel[4][1] ~^ image[12][14] + signed_kernel[4][2] ~^ image[12][15] + signed_kernel[4][3] ~^ image[12][16] + signed_kernel[4][4] ~^ image[12][17];
assign xor_sum[8][14] = signed_kernel[0][0] ~^ image[8][14] + signed_kernel[0][1] ~^ image[8][15] + signed_kernel[0][2] ~^ image[8][16] + signed_kernel[0][3] ~^ image[8][17] + signed_kernel[0][4] ~^ image[8][18] + signed_kernel[1][0] ~^ image[9][14] + signed_kernel[1][1] ~^ image[9][15] + signed_kernel[1][2] ~^ image[9][16] + signed_kernel[1][3] ~^ image[9][17] + signed_kernel[1][4] ~^ image[9][18] + signed_kernel[2][0] ~^ image[10][14] + signed_kernel[2][1] ~^ image[10][15] + signed_kernel[2][2] ~^ image[10][16] + signed_kernel[2][3] ~^ image[10][17] + signed_kernel[2][4] ~^ image[10][18] + signed_kernel[3][0] ~^ image[11][14] + signed_kernel[3][1] ~^ image[11][15] + signed_kernel[3][2] ~^ image[11][16] + signed_kernel[3][3] ~^ image[11][17] + signed_kernel[3][4] ~^ image[11][18] + signed_kernel[4][0] ~^ image[12][14] + signed_kernel[4][1] ~^ image[12][15] + signed_kernel[4][2] ~^ image[12][16] + signed_kernel[4][3] ~^ image[12][17] + signed_kernel[4][4] ~^ image[12][18];
assign xor_sum[8][15] = signed_kernel[0][0] ~^ image[8][15] + signed_kernel[0][1] ~^ image[8][16] + signed_kernel[0][2] ~^ image[8][17] + signed_kernel[0][3] ~^ image[8][18] + signed_kernel[0][4] ~^ image[8][19] + signed_kernel[1][0] ~^ image[9][15] + signed_kernel[1][1] ~^ image[9][16] + signed_kernel[1][2] ~^ image[9][17] + signed_kernel[1][3] ~^ image[9][18] + signed_kernel[1][4] ~^ image[9][19] + signed_kernel[2][0] ~^ image[10][15] + signed_kernel[2][1] ~^ image[10][16] + signed_kernel[2][2] ~^ image[10][17] + signed_kernel[2][3] ~^ image[10][18] + signed_kernel[2][4] ~^ image[10][19] + signed_kernel[3][0] ~^ image[11][15] + signed_kernel[3][1] ~^ image[11][16] + signed_kernel[3][2] ~^ image[11][17] + signed_kernel[3][3] ~^ image[11][18] + signed_kernel[3][4] ~^ image[11][19] + signed_kernel[4][0] ~^ image[12][15] + signed_kernel[4][1] ~^ image[12][16] + signed_kernel[4][2] ~^ image[12][17] + signed_kernel[4][3] ~^ image[12][18] + signed_kernel[4][4] ~^ image[12][19];
assign xor_sum[8][16] = signed_kernel[0][0] ~^ image[8][16] + signed_kernel[0][1] ~^ image[8][17] + signed_kernel[0][2] ~^ image[8][18] + signed_kernel[0][3] ~^ image[8][19] + signed_kernel[0][4] ~^ image[8][20] + signed_kernel[1][0] ~^ image[9][16] + signed_kernel[1][1] ~^ image[9][17] + signed_kernel[1][2] ~^ image[9][18] + signed_kernel[1][3] ~^ image[9][19] + signed_kernel[1][4] ~^ image[9][20] + signed_kernel[2][0] ~^ image[10][16] + signed_kernel[2][1] ~^ image[10][17] + signed_kernel[2][2] ~^ image[10][18] + signed_kernel[2][3] ~^ image[10][19] + signed_kernel[2][4] ~^ image[10][20] + signed_kernel[3][0] ~^ image[11][16] + signed_kernel[3][1] ~^ image[11][17] + signed_kernel[3][2] ~^ image[11][18] + signed_kernel[3][3] ~^ image[11][19] + signed_kernel[3][4] ~^ image[11][20] + signed_kernel[4][0] ~^ image[12][16] + signed_kernel[4][1] ~^ image[12][17] + signed_kernel[4][2] ~^ image[12][18] + signed_kernel[4][3] ~^ image[12][19] + signed_kernel[4][4] ~^ image[12][20];
assign xor_sum[8][17] = signed_kernel[0][0] ~^ image[8][17] + signed_kernel[0][1] ~^ image[8][18] + signed_kernel[0][2] ~^ image[8][19] + signed_kernel[0][3] ~^ image[8][20] + signed_kernel[0][4] ~^ image[8][21] + signed_kernel[1][0] ~^ image[9][17] + signed_kernel[1][1] ~^ image[9][18] + signed_kernel[1][2] ~^ image[9][19] + signed_kernel[1][3] ~^ image[9][20] + signed_kernel[1][4] ~^ image[9][21] + signed_kernel[2][0] ~^ image[10][17] + signed_kernel[2][1] ~^ image[10][18] + signed_kernel[2][2] ~^ image[10][19] + signed_kernel[2][3] ~^ image[10][20] + signed_kernel[2][4] ~^ image[10][21] + signed_kernel[3][0] ~^ image[11][17] + signed_kernel[3][1] ~^ image[11][18] + signed_kernel[3][2] ~^ image[11][19] + signed_kernel[3][3] ~^ image[11][20] + signed_kernel[3][4] ~^ image[11][21] + signed_kernel[4][0] ~^ image[12][17] + signed_kernel[4][1] ~^ image[12][18] + signed_kernel[4][2] ~^ image[12][19] + signed_kernel[4][3] ~^ image[12][20] + signed_kernel[4][4] ~^ image[12][21];
assign xor_sum[8][18] = signed_kernel[0][0] ~^ image[8][18] + signed_kernel[0][1] ~^ image[8][19] + signed_kernel[0][2] ~^ image[8][20] + signed_kernel[0][3] ~^ image[8][21] + signed_kernel[0][4] ~^ image[8][22] + signed_kernel[1][0] ~^ image[9][18] + signed_kernel[1][1] ~^ image[9][19] + signed_kernel[1][2] ~^ image[9][20] + signed_kernel[1][3] ~^ image[9][21] + signed_kernel[1][4] ~^ image[9][22] + signed_kernel[2][0] ~^ image[10][18] + signed_kernel[2][1] ~^ image[10][19] + signed_kernel[2][2] ~^ image[10][20] + signed_kernel[2][3] ~^ image[10][21] + signed_kernel[2][4] ~^ image[10][22] + signed_kernel[3][0] ~^ image[11][18] + signed_kernel[3][1] ~^ image[11][19] + signed_kernel[3][2] ~^ image[11][20] + signed_kernel[3][3] ~^ image[11][21] + signed_kernel[3][4] ~^ image[11][22] + signed_kernel[4][0] ~^ image[12][18] + signed_kernel[4][1] ~^ image[12][19] + signed_kernel[4][2] ~^ image[12][20] + signed_kernel[4][3] ~^ image[12][21] + signed_kernel[4][4] ~^ image[12][22];
assign xor_sum[8][19] = signed_kernel[0][0] ~^ image[8][19] + signed_kernel[0][1] ~^ image[8][20] + signed_kernel[0][2] ~^ image[8][21] + signed_kernel[0][3] ~^ image[8][22] + signed_kernel[0][4] ~^ image[8][23] + signed_kernel[1][0] ~^ image[9][19] + signed_kernel[1][1] ~^ image[9][20] + signed_kernel[1][2] ~^ image[9][21] + signed_kernel[1][3] ~^ image[9][22] + signed_kernel[1][4] ~^ image[9][23] + signed_kernel[2][0] ~^ image[10][19] + signed_kernel[2][1] ~^ image[10][20] + signed_kernel[2][2] ~^ image[10][21] + signed_kernel[2][3] ~^ image[10][22] + signed_kernel[2][4] ~^ image[10][23] + signed_kernel[3][0] ~^ image[11][19] + signed_kernel[3][1] ~^ image[11][20] + signed_kernel[3][2] ~^ image[11][21] + signed_kernel[3][3] ~^ image[11][22] + signed_kernel[3][4] ~^ image[11][23] + signed_kernel[4][0] ~^ image[12][19] + signed_kernel[4][1] ~^ image[12][20] + signed_kernel[4][2] ~^ image[12][21] + signed_kernel[4][3] ~^ image[12][22] + signed_kernel[4][4] ~^ image[12][23];
assign xor_sum[8][20] = signed_kernel[0][0] ~^ image[8][20] + signed_kernel[0][1] ~^ image[8][21] + signed_kernel[0][2] ~^ image[8][22] + signed_kernel[0][3] ~^ image[8][23] + signed_kernel[0][4] ~^ image[8][24] + signed_kernel[1][0] ~^ image[9][20] + signed_kernel[1][1] ~^ image[9][21] + signed_kernel[1][2] ~^ image[9][22] + signed_kernel[1][3] ~^ image[9][23] + signed_kernel[1][4] ~^ image[9][24] + signed_kernel[2][0] ~^ image[10][20] + signed_kernel[2][1] ~^ image[10][21] + signed_kernel[2][2] ~^ image[10][22] + signed_kernel[2][3] ~^ image[10][23] + signed_kernel[2][4] ~^ image[10][24] + signed_kernel[3][0] ~^ image[11][20] + signed_kernel[3][1] ~^ image[11][21] + signed_kernel[3][2] ~^ image[11][22] + signed_kernel[3][3] ~^ image[11][23] + signed_kernel[3][4] ~^ image[11][24] + signed_kernel[4][0] ~^ image[12][20] + signed_kernel[4][1] ~^ image[12][21] + signed_kernel[4][2] ~^ image[12][22] + signed_kernel[4][3] ~^ image[12][23] + signed_kernel[4][4] ~^ image[12][24];
assign xor_sum[8][21] = signed_kernel[0][0] ~^ image[8][21] + signed_kernel[0][1] ~^ image[8][22] + signed_kernel[0][2] ~^ image[8][23] + signed_kernel[0][3] ~^ image[8][24] + signed_kernel[0][4] ~^ image[8][25] + signed_kernel[1][0] ~^ image[9][21] + signed_kernel[1][1] ~^ image[9][22] + signed_kernel[1][2] ~^ image[9][23] + signed_kernel[1][3] ~^ image[9][24] + signed_kernel[1][4] ~^ image[9][25] + signed_kernel[2][0] ~^ image[10][21] + signed_kernel[2][1] ~^ image[10][22] + signed_kernel[2][2] ~^ image[10][23] + signed_kernel[2][3] ~^ image[10][24] + signed_kernel[2][4] ~^ image[10][25] + signed_kernel[3][0] ~^ image[11][21] + signed_kernel[3][1] ~^ image[11][22] + signed_kernel[3][2] ~^ image[11][23] + signed_kernel[3][3] ~^ image[11][24] + signed_kernel[3][4] ~^ image[11][25] + signed_kernel[4][0] ~^ image[12][21] + signed_kernel[4][1] ~^ image[12][22] + signed_kernel[4][2] ~^ image[12][23] + signed_kernel[4][3] ~^ image[12][24] + signed_kernel[4][4] ~^ image[12][25];
assign xor_sum[8][22] = signed_kernel[0][0] ~^ image[8][22] + signed_kernel[0][1] ~^ image[8][23] + signed_kernel[0][2] ~^ image[8][24] + signed_kernel[0][3] ~^ image[8][25] + signed_kernel[0][4] ~^ image[8][26] + signed_kernel[1][0] ~^ image[9][22] + signed_kernel[1][1] ~^ image[9][23] + signed_kernel[1][2] ~^ image[9][24] + signed_kernel[1][3] ~^ image[9][25] + signed_kernel[1][4] ~^ image[9][26] + signed_kernel[2][0] ~^ image[10][22] + signed_kernel[2][1] ~^ image[10][23] + signed_kernel[2][2] ~^ image[10][24] + signed_kernel[2][3] ~^ image[10][25] + signed_kernel[2][4] ~^ image[10][26] + signed_kernel[3][0] ~^ image[11][22] + signed_kernel[3][1] ~^ image[11][23] + signed_kernel[3][2] ~^ image[11][24] + signed_kernel[3][3] ~^ image[11][25] + signed_kernel[3][4] ~^ image[11][26] + signed_kernel[4][0] ~^ image[12][22] + signed_kernel[4][1] ~^ image[12][23] + signed_kernel[4][2] ~^ image[12][24] + signed_kernel[4][3] ~^ image[12][25] + signed_kernel[4][4] ~^ image[12][26];
assign xor_sum[8][23] = signed_kernel[0][0] ~^ image[8][23] + signed_kernel[0][1] ~^ image[8][24] + signed_kernel[0][2] ~^ image[8][25] + signed_kernel[0][3] ~^ image[8][26] + signed_kernel[0][4] ~^ image[8][27] + signed_kernel[1][0] ~^ image[9][23] + signed_kernel[1][1] ~^ image[9][24] + signed_kernel[1][2] ~^ image[9][25] + signed_kernel[1][3] ~^ image[9][26] + signed_kernel[1][4] ~^ image[9][27] + signed_kernel[2][0] ~^ image[10][23] + signed_kernel[2][1] ~^ image[10][24] + signed_kernel[2][2] ~^ image[10][25] + signed_kernel[2][3] ~^ image[10][26] + signed_kernel[2][4] ~^ image[10][27] + signed_kernel[3][0] ~^ image[11][23] + signed_kernel[3][1] ~^ image[11][24] + signed_kernel[3][2] ~^ image[11][25] + signed_kernel[3][3] ~^ image[11][26] + signed_kernel[3][4] ~^ image[11][27] + signed_kernel[4][0] ~^ image[12][23] + signed_kernel[4][1] ~^ image[12][24] + signed_kernel[4][2] ~^ image[12][25] + signed_kernel[4][3] ~^ image[12][26] + signed_kernel[4][4] ~^ image[12][27];
assign xor_sum[9][0] = signed_kernel[0][0] ~^ image[9][0] + signed_kernel[0][1] ~^ image[9][1] + signed_kernel[0][2] ~^ image[9][2] + signed_kernel[0][3] ~^ image[9][3] + signed_kernel[0][4] ~^ image[9][4] + signed_kernel[1][0] ~^ image[10][0] + signed_kernel[1][1] ~^ image[10][1] + signed_kernel[1][2] ~^ image[10][2] + signed_kernel[1][3] ~^ image[10][3] + signed_kernel[1][4] ~^ image[10][4] + signed_kernel[2][0] ~^ image[11][0] + signed_kernel[2][1] ~^ image[11][1] + signed_kernel[2][2] ~^ image[11][2] + signed_kernel[2][3] ~^ image[11][3] + signed_kernel[2][4] ~^ image[11][4] + signed_kernel[3][0] ~^ image[12][0] + signed_kernel[3][1] ~^ image[12][1] + signed_kernel[3][2] ~^ image[12][2] + signed_kernel[3][3] ~^ image[12][3] + signed_kernel[3][4] ~^ image[12][4] + signed_kernel[4][0] ~^ image[13][0] + signed_kernel[4][1] ~^ image[13][1] + signed_kernel[4][2] ~^ image[13][2] + signed_kernel[4][3] ~^ image[13][3] + signed_kernel[4][4] ~^ image[13][4];
assign xor_sum[9][1] = signed_kernel[0][0] ~^ image[9][1] + signed_kernel[0][1] ~^ image[9][2] + signed_kernel[0][2] ~^ image[9][3] + signed_kernel[0][3] ~^ image[9][4] + signed_kernel[0][4] ~^ image[9][5] + signed_kernel[1][0] ~^ image[10][1] + signed_kernel[1][1] ~^ image[10][2] + signed_kernel[1][2] ~^ image[10][3] + signed_kernel[1][3] ~^ image[10][4] + signed_kernel[1][4] ~^ image[10][5] + signed_kernel[2][0] ~^ image[11][1] + signed_kernel[2][1] ~^ image[11][2] + signed_kernel[2][2] ~^ image[11][3] + signed_kernel[2][3] ~^ image[11][4] + signed_kernel[2][4] ~^ image[11][5] + signed_kernel[3][0] ~^ image[12][1] + signed_kernel[3][1] ~^ image[12][2] + signed_kernel[3][2] ~^ image[12][3] + signed_kernel[3][3] ~^ image[12][4] + signed_kernel[3][4] ~^ image[12][5] + signed_kernel[4][0] ~^ image[13][1] + signed_kernel[4][1] ~^ image[13][2] + signed_kernel[4][2] ~^ image[13][3] + signed_kernel[4][3] ~^ image[13][4] + signed_kernel[4][4] ~^ image[13][5];
assign xor_sum[9][2] = signed_kernel[0][0] ~^ image[9][2] + signed_kernel[0][1] ~^ image[9][3] + signed_kernel[0][2] ~^ image[9][4] + signed_kernel[0][3] ~^ image[9][5] + signed_kernel[0][4] ~^ image[9][6] + signed_kernel[1][0] ~^ image[10][2] + signed_kernel[1][1] ~^ image[10][3] + signed_kernel[1][2] ~^ image[10][4] + signed_kernel[1][3] ~^ image[10][5] + signed_kernel[1][4] ~^ image[10][6] + signed_kernel[2][0] ~^ image[11][2] + signed_kernel[2][1] ~^ image[11][3] + signed_kernel[2][2] ~^ image[11][4] + signed_kernel[2][3] ~^ image[11][5] + signed_kernel[2][4] ~^ image[11][6] + signed_kernel[3][0] ~^ image[12][2] + signed_kernel[3][1] ~^ image[12][3] + signed_kernel[3][2] ~^ image[12][4] + signed_kernel[3][3] ~^ image[12][5] + signed_kernel[3][4] ~^ image[12][6] + signed_kernel[4][0] ~^ image[13][2] + signed_kernel[4][1] ~^ image[13][3] + signed_kernel[4][2] ~^ image[13][4] + signed_kernel[4][3] ~^ image[13][5] + signed_kernel[4][4] ~^ image[13][6];
assign xor_sum[9][3] = signed_kernel[0][0] ~^ image[9][3] + signed_kernel[0][1] ~^ image[9][4] + signed_kernel[0][2] ~^ image[9][5] + signed_kernel[0][3] ~^ image[9][6] + signed_kernel[0][4] ~^ image[9][7] + signed_kernel[1][0] ~^ image[10][3] + signed_kernel[1][1] ~^ image[10][4] + signed_kernel[1][2] ~^ image[10][5] + signed_kernel[1][3] ~^ image[10][6] + signed_kernel[1][4] ~^ image[10][7] + signed_kernel[2][0] ~^ image[11][3] + signed_kernel[2][1] ~^ image[11][4] + signed_kernel[2][2] ~^ image[11][5] + signed_kernel[2][3] ~^ image[11][6] + signed_kernel[2][4] ~^ image[11][7] + signed_kernel[3][0] ~^ image[12][3] + signed_kernel[3][1] ~^ image[12][4] + signed_kernel[3][2] ~^ image[12][5] + signed_kernel[3][3] ~^ image[12][6] + signed_kernel[3][4] ~^ image[12][7] + signed_kernel[4][0] ~^ image[13][3] + signed_kernel[4][1] ~^ image[13][4] + signed_kernel[4][2] ~^ image[13][5] + signed_kernel[4][3] ~^ image[13][6] + signed_kernel[4][4] ~^ image[13][7];
assign xor_sum[9][4] = signed_kernel[0][0] ~^ image[9][4] + signed_kernel[0][1] ~^ image[9][5] + signed_kernel[0][2] ~^ image[9][6] + signed_kernel[0][3] ~^ image[9][7] + signed_kernel[0][4] ~^ image[9][8] + signed_kernel[1][0] ~^ image[10][4] + signed_kernel[1][1] ~^ image[10][5] + signed_kernel[1][2] ~^ image[10][6] + signed_kernel[1][3] ~^ image[10][7] + signed_kernel[1][4] ~^ image[10][8] + signed_kernel[2][0] ~^ image[11][4] + signed_kernel[2][1] ~^ image[11][5] + signed_kernel[2][2] ~^ image[11][6] + signed_kernel[2][3] ~^ image[11][7] + signed_kernel[2][4] ~^ image[11][8] + signed_kernel[3][0] ~^ image[12][4] + signed_kernel[3][1] ~^ image[12][5] + signed_kernel[3][2] ~^ image[12][6] + signed_kernel[3][3] ~^ image[12][7] + signed_kernel[3][4] ~^ image[12][8] + signed_kernel[4][0] ~^ image[13][4] + signed_kernel[4][1] ~^ image[13][5] + signed_kernel[4][2] ~^ image[13][6] + signed_kernel[4][3] ~^ image[13][7] + signed_kernel[4][4] ~^ image[13][8];
assign xor_sum[9][5] = signed_kernel[0][0] ~^ image[9][5] + signed_kernel[0][1] ~^ image[9][6] + signed_kernel[0][2] ~^ image[9][7] + signed_kernel[0][3] ~^ image[9][8] + signed_kernel[0][4] ~^ image[9][9] + signed_kernel[1][0] ~^ image[10][5] + signed_kernel[1][1] ~^ image[10][6] + signed_kernel[1][2] ~^ image[10][7] + signed_kernel[1][3] ~^ image[10][8] + signed_kernel[1][4] ~^ image[10][9] + signed_kernel[2][0] ~^ image[11][5] + signed_kernel[2][1] ~^ image[11][6] + signed_kernel[2][2] ~^ image[11][7] + signed_kernel[2][3] ~^ image[11][8] + signed_kernel[2][4] ~^ image[11][9] + signed_kernel[3][0] ~^ image[12][5] + signed_kernel[3][1] ~^ image[12][6] + signed_kernel[3][2] ~^ image[12][7] + signed_kernel[3][3] ~^ image[12][8] + signed_kernel[3][4] ~^ image[12][9] + signed_kernel[4][0] ~^ image[13][5] + signed_kernel[4][1] ~^ image[13][6] + signed_kernel[4][2] ~^ image[13][7] + signed_kernel[4][3] ~^ image[13][8] + signed_kernel[4][4] ~^ image[13][9];
assign xor_sum[9][6] = signed_kernel[0][0] ~^ image[9][6] + signed_kernel[0][1] ~^ image[9][7] + signed_kernel[0][2] ~^ image[9][8] + signed_kernel[0][3] ~^ image[9][9] + signed_kernel[0][4] ~^ image[9][10] + signed_kernel[1][0] ~^ image[10][6] + signed_kernel[1][1] ~^ image[10][7] + signed_kernel[1][2] ~^ image[10][8] + signed_kernel[1][3] ~^ image[10][9] + signed_kernel[1][4] ~^ image[10][10] + signed_kernel[2][0] ~^ image[11][6] + signed_kernel[2][1] ~^ image[11][7] + signed_kernel[2][2] ~^ image[11][8] + signed_kernel[2][3] ~^ image[11][9] + signed_kernel[2][4] ~^ image[11][10] + signed_kernel[3][0] ~^ image[12][6] + signed_kernel[3][1] ~^ image[12][7] + signed_kernel[3][2] ~^ image[12][8] + signed_kernel[3][3] ~^ image[12][9] + signed_kernel[3][4] ~^ image[12][10] + signed_kernel[4][0] ~^ image[13][6] + signed_kernel[4][1] ~^ image[13][7] + signed_kernel[4][2] ~^ image[13][8] + signed_kernel[4][3] ~^ image[13][9] + signed_kernel[4][4] ~^ image[13][10];
assign xor_sum[9][7] = signed_kernel[0][0] ~^ image[9][7] + signed_kernel[0][1] ~^ image[9][8] + signed_kernel[0][2] ~^ image[9][9] + signed_kernel[0][3] ~^ image[9][10] + signed_kernel[0][4] ~^ image[9][11] + signed_kernel[1][0] ~^ image[10][7] + signed_kernel[1][1] ~^ image[10][8] + signed_kernel[1][2] ~^ image[10][9] + signed_kernel[1][3] ~^ image[10][10] + signed_kernel[1][4] ~^ image[10][11] + signed_kernel[2][0] ~^ image[11][7] + signed_kernel[2][1] ~^ image[11][8] + signed_kernel[2][2] ~^ image[11][9] + signed_kernel[2][3] ~^ image[11][10] + signed_kernel[2][4] ~^ image[11][11] + signed_kernel[3][0] ~^ image[12][7] + signed_kernel[3][1] ~^ image[12][8] + signed_kernel[3][2] ~^ image[12][9] + signed_kernel[3][3] ~^ image[12][10] + signed_kernel[3][4] ~^ image[12][11] + signed_kernel[4][0] ~^ image[13][7] + signed_kernel[4][1] ~^ image[13][8] + signed_kernel[4][2] ~^ image[13][9] + signed_kernel[4][3] ~^ image[13][10] + signed_kernel[4][4] ~^ image[13][11];
assign xor_sum[9][8] = signed_kernel[0][0] ~^ image[9][8] + signed_kernel[0][1] ~^ image[9][9] + signed_kernel[0][2] ~^ image[9][10] + signed_kernel[0][3] ~^ image[9][11] + signed_kernel[0][4] ~^ image[9][12] + signed_kernel[1][0] ~^ image[10][8] + signed_kernel[1][1] ~^ image[10][9] + signed_kernel[1][2] ~^ image[10][10] + signed_kernel[1][3] ~^ image[10][11] + signed_kernel[1][4] ~^ image[10][12] + signed_kernel[2][0] ~^ image[11][8] + signed_kernel[2][1] ~^ image[11][9] + signed_kernel[2][2] ~^ image[11][10] + signed_kernel[2][3] ~^ image[11][11] + signed_kernel[2][4] ~^ image[11][12] + signed_kernel[3][0] ~^ image[12][8] + signed_kernel[3][1] ~^ image[12][9] + signed_kernel[3][2] ~^ image[12][10] + signed_kernel[3][3] ~^ image[12][11] + signed_kernel[3][4] ~^ image[12][12] + signed_kernel[4][0] ~^ image[13][8] + signed_kernel[4][1] ~^ image[13][9] + signed_kernel[4][2] ~^ image[13][10] + signed_kernel[4][3] ~^ image[13][11] + signed_kernel[4][4] ~^ image[13][12];
assign xor_sum[9][9] = signed_kernel[0][0] ~^ image[9][9] + signed_kernel[0][1] ~^ image[9][10] + signed_kernel[0][2] ~^ image[9][11] + signed_kernel[0][3] ~^ image[9][12] + signed_kernel[0][4] ~^ image[9][13] + signed_kernel[1][0] ~^ image[10][9] + signed_kernel[1][1] ~^ image[10][10] + signed_kernel[1][2] ~^ image[10][11] + signed_kernel[1][3] ~^ image[10][12] + signed_kernel[1][4] ~^ image[10][13] + signed_kernel[2][0] ~^ image[11][9] + signed_kernel[2][1] ~^ image[11][10] + signed_kernel[2][2] ~^ image[11][11] + signed_kernel[2][3] ~^ image[11][12] + signed_kernel[2][4] ~^ image[11][13] + signed_kernel[3][0] ~^ image[12][9] + signed_kernel[3][1] ~^ image[12][10] + signed_kernel[3][2] ~^ image[12][11] + signed_kernel[3][3] ~^ image[12][12] + signed_kernel[3][4] ~^ image[12][13] + signed_kernel[4][0] ~^ image[13][9] + signed_kernel[4][1] ~^ image[13][10] + signed_kernel[4][2] ~^ image[13][11] + signed_kernel[4][3] ~^ image[13][12] + signed_kernel[4][4] ~^ image[13][13];
assign xor_sum[9][10] = signed_kernel[0][0] ~^ image[9][10] + signed_kernel[0][1] ~^ image[9][11] + signed_kernel[0][2] ~^ image[9][12] + signed_kernel[0][3] ~^ image[9][13] + signed_kernel[0][4] ~^ image[9][14] + signed_kernel[1][0] ~^ image[10][10] + signed_kernel[1][1] ~^ image[10][11] + signed_kernel[1][2] ~^ image[10][12] + signed_kernel[1][3] ~^ image[10][13] + signed_kernel[1][4] ~^ image[10][14] + signed_kernel[2][0] ~^ image[11][10] + signed_kernel[2][1] ~^ image[11][11] + signed_kernel[2][2] ~^ image[11][12] + signed_kernel[2][3] ~^ image[11][13] + signed_kernel[2][4] ~^ image[11][14] + signed_kernel[3][0] ~^ image[12][10] + signed_kernel[3][1] ~^ image[12][11] + signed_kernel[3][2] ~^ image[12][12] + signed_kernel[3][3] ~^ image[12][13] + signed_kernel[3][4] ~^ image[12][14] + signed_kernel[4][0] ~^ image[13][10] + signed_kernel[4][1] ~^ image[13][11] + signed_kernel[4][2] ~^ image[13][12] + signed_kernel[4][3] ~^ image[13][13] + signed_kernel[4][4] ~^ image[13][14];
assign xor_sum[9][11] = signed_kernel[0][0] ~^ image[9][11] + signed_kernel[0][1] ~^ image[9][12] + signed_kernel[0][2] ~^ image[9][13] + signed_kernel[0][3] ~^ image[9][14] + signed_kernel[0][4] ~^ image[9][15] + signed_kernel[1][0] ~^ image[10][11] + signed_kernel[1][1] ~^ image[10][12] + signed_kernel[1][2] ~^ image[10][13] + signed_kernel[1][3] ~^ image[10][14] + signed_kernel[1][4] ~^ image[10][15] + signed_kernel[2][0] ~^ image[11][11] + signed_kernel[2][1] ~^ image[11][12] + signed_kernel[2][2] ~^ image[11][13] + signed_kernel[2][3] ~^ image[11][14] + signed_kernel[2][4] ~^ image[11][15] + signed_kernel[3][0] ~^ image[12][11] + signed_kernel[3][1] ~^ image[12][12] + signed_kernel[3][2] ~^ image[12][13] + signed_kernel[3][3] ~^ image[12][14] + signed_kernel[3][4] ~^ image[12][15] + signed_kernel[4][0] ~^ image[13][11] + signed_kernel[4][1] ~^ image[13][12] + signed_kernel[4][2] ~^ image[13][13] + signed_kernel[4][3] ~^ image[13][14] + signed_kernel[4][4] ~^ image[13][15];
assign xor_sum[9][12] = signed_kernel[0][0] ~^ image[9][12] + signed_kernel[0][1] ~^ image[9][13] + signed_kernel[0][2] ~^ image[9][14] + signed_kernel[0][3] ~^ image[9][15] + signed_kernel[0][4] ~^ image[9][16] + signed_kernel[1][0] ~^ image[10][12] + signed_kernel[1][1] ~^ image[10][13] + signed_kernel[1][2] ~^ image[10][14] + signed_kernel[1][3] ~^ image[10][15] + signed_kernel[1][4] ~^ image[10][16] + signed_kernel[2][0] ~^ image[11][12] + signed_kernel[2][1] ~^ image[11][13] + signed_kernel[2][2] ~^ image[11][14] + signed_kernel[2][3] ~^ image[11][15] + signed_kernel[2][4] ~^ image[11][16] + signed_kernel[3][0] ~^ image[12][12] + signed_kernel[3][1] ~^ image[12][13] + signed_kernel[3][2] ~^ image[12][14] + signed_kernel[3][3] ~^ image[12][15] + signed_kernel[3][4] ~^ image[12][16] + signed_kernel[4][0] ~^ image[13][12] + signed_kernel[4][1] ~^ image[13][13] + signed_kernel[4][2] ~^ image[13][14] + signed_kernel[4][3] ~^ image[13][15] + signed_kernel[4][4] ~^ image[13][16];
assign xor_sum[9][13] = signed_kernel[0][0] ~^ image[9][13] + signed_kernel[0][1] ~^ image[9][14] + signed_kernel[0][2] ~^ image[9][15] + signed_kernel[0][3] ~^ image[9][16] + signed_kernel[0][4] ~^ image[9][17] + signed_kernel[1][0] ~^ image[10][13] + signed_kernel[1][1] ~^ image[10][14] + signed_kernel[1][2] ~^ image[10][15] + signed_kernel[1][3] ~^ image[10][16] + signed_kernel[1][4] ~^ image[10][17] + signed_kernel[2][0] ~^ image[11][13] + signed_kernel[2][1] ~^ image[11][14] + signed_kernel[2][2] ~^ image[11][15] + signed_kernel[2][3] ~^ image[11][16] + signed_kernel[2][4] ~^ image[11][17] + signed_kernel[3][0] ~^ image[12][13] + signed_kernel[3][1] ~^ image[12][14] + signed_kernel[3][2] ~^ image[12][15] + signed_kernel[3][3] ~^ image[12][16] + signed_kernel[3][4] ~^ image[12][17] + signed_kernel[4][0] ~^ image[13][13] + signed_kernel[4][1] ~^ image[13][14] + signed_kernel[4][2] ~^ image[13][15] + signed_kernel[4][3] ~^ image[13][16] + signed_kernel[4][4] ~^ image[13][17];
assign xor_sum[9][14] = signed_kernel[0][0] ~^ image[9][14] + signed_kernel[0][1] ~^ image[9][15] + signed_kernel[0][2] ~^ image[9][16] + signed_kernel[0][3] ~^ image[9][17] + signed_kernel[0][4] ~^ image[9][18] + signed_kernel[1][0] ~^ image[10][14] + signed_kernel[1][1] ~^ image[10][15] + signed_kernel[1][2] ~^ image[10][16] + signed_kernel[1][3] ~^ image[10][17] + signed_kernel[1][4] ~^ image[10][18] + signed_kernel[2][0] ~^ image[11][14] + signed_kernel[2][1] ~^ image[11][15] + signed_kernel[2][2] ~^ image[11][16] + signed_kernel[2][3] ~^ image[11][17] + signed_kernel[2][4] ~^ image[11][18] + signed_kernel[3][0] ~^ image[12][14] + signed_kernel[3][1] ~^ image[12][15] + signed_kernel[3][2] ~^ image[12][16] + signed_kernel[3][3] ~^ image[12][17] + signed_kernel[3][4] ~^ image[12][18] + signed_kernel[4][0] ~^ image[13][14] + signed_kernel[4][1] ~^ image[13][15] + signed_kernel[4][2] ~^ image[13][16] + signed_kernel[4][3] ~^ image[13][17] + signed_kernel[4][4] ~^ image[13][18];
assign xor_sum[9][15] = signed_kernel[0][0] ~^ image[9][15] + signed_kernel[0][1] ~^ image[9][16] + signed_kernel[0][2] ~^ image[9][17] + signed_kernel[0][3] ~^ image[9][18] + signed_kernel[0][4] ~^ image[9][19] + signed_kernel[1][0] ~^ image[10][15] + signed_kernel[1][1] ~^ image[10][16] + signed_kernel[1][2] ~^ image[10][17] + signed_kernel[1][3] ~^ image[10][18] + signed_kernel[1][4] ~^ image[10][19] + signed_kernel[2][0] ~^ image[11][15] + signed_kernel[2][1] ~^ image[11][16] + signed_kernel[2][2] ~^ image[11][17] + signed_kernel[2][3] ~^ image[11][18] + signed_kernel[2][4] ~^ image[11][19] + signed_kernel[3][0] ~^ image[12][15] + signed_kernel[3][1] ~^ image[12][16] + signed_kernel[3][2] ~^ image[12][17] + signed_kernel[3][3] ~^ image[12][18] + signed_kernel[3][4] ~^ image[12][19] + signed_kernel[4][0] ~^ image[13][15] + signed_kernel[4][1] ~^ image[13][16] + signed_kernel[4][2] ~^ image[13][17] + signed_kernel[4][3] ~^ image[13][18] + signed_kernel[4][4] ~^ image[13][19];
assign xor_sum[9][16] = signed_kernel[0][0] ~^ image[9][16] + signed_kernel[0][1] ~^ image[9][17] + signed_kernel[0][2] ~^ image[9][18] + signed_kernel[0][3] ~^ image[9][19] + signed_kernel[0][4] ~^ image[9][20] + signed_kernel[1][0] ~^ image[10][16] + signed_kernel[1][1] ~^ image[10][17] + signed_kernel[1][2] ~^ image[10][18] + signed_kernel[1][3] ~^ image[10][19] + signed_kernel[1][4] ~^ image[10][20] + signed_kernel[2][0] ~^ image[11][16] + signed_kernel[2][1] ~^ image[11][17] + signed_kernel[2][2] ~^ image[11][18] + signed_kernel[2][3] ~^ image[11][19] + signed_kernel[2][4] ~^ image[11][20] + signed_kernel[3][0] ~^ image[12][16] + signed_kernel[3][1] ~^ image[12][17] + signed_kernel[3][2] ~^ image[12][18] + signed_kernel[3][3] ~^ image[12][19] + signed_kernel[3][4] ~^ image[12][20] + signed_kernel[4][0] ~^ image[13][16] + signed_kernel[4][1] ~^ image[13][17] + signed_kernel[4][2] ~^ image[13][18] + signed_kernel[4][3] ~^ image[13][19] + signed_kernel[4][4] ~^ image[13][20];
assign xor_sum[9][17] = signed_kernel[0][0] ~^ image[9][17] + signed_kernel[0][1] ~^ image[9][18] + signed_kernel[0][2] ~^ image[9][19] + signed_kernel[0][3] ~^ image[9][20] + signed_kernel[0][4] ~^ image[9][21] + signed_kernel[1][0] ~^ image[10][17] + signed_kernel[1][1] ~^ image[10][18] + signed_kernel[1][2] ~^ image[10][19] + signed_kernel[1][3] ~^ image[10][20] + signed_kernel[1][4] ~^ image[10][21] + signed_kernel[2][0] ~^ image[11][17] + signed_kernel[2][1] ~^ image[11][18] + signed_kernel[2][2] ~^ image[11][19] + signed_kernel[2][3] ~^ image[11][20] + signed_kernel[2][4] ~^ image[11][21] + signed_kernel[3][0] ~^ image[12][17] + signed_kernel[3][1] ~^ image[12][18] + signed_kernel[3][2] ~^ image[12][19] + signed_kernel[3][3] ~^ image[12][20] + signed_kernel[3][4] ~^ image[12][21] + signed_kernel[4][0] ~^ image[13][17] + signed_kernel[4][1] ~^ image[13][18] + signed_kernel[4][2] ~^ image[13][19] + signed_kernel[4][3] ~^ image[13][20] + signed_kernel[4][4] ~^ image[13][21];
assign xor_sum[9][18] = signed_kernel[0][0] ~^ image[9][18] + signed_kernel[0][1] ~^ image[9][19] + signed_kernel[0][2] ~^ image[9][20] + signed_kernel[0][3] ~^ image[9][21] + signed_kernel[0][4] ~^ image[9][22] + signed_kernel[1][0] ~^ image[10][18] + signed_kernel[1][1] ~^ image[10][19] + signed_kernel[1][2] ~^ image[10][20] + signed_kernel[1][3] ~^ image[10][21] + signed_kernel[1][4] ~^ image[10][22] + signed_kernel[2][0] ~^ image[11][18] + signed_kernel[2][1] ~^ image[11][19] + signed_kernel[2][2] ~^ image[11][20] + signed_kernel[2][3] ~^ image[11][21] + signed_kernel[2][4] ~^ image[11][22] + signed_kernel[3][0] ~^ image[12][18] + signed_kernel[3][1] ~^ image[12][19] + signed_kernel[3][2] ~^ image[12][20] + signed_kernel[3][3] ~^ image[12][21] + signed_kernel[3][4] ~^ image[12][22] + signed_kernel[4][0] ~^ image[13][18] + signed_kernel[4][1] ~^ image[13][19] + signed_kernel[4][2] ~^ image[13][20] + signed_kernel[4][3] ~^ image[13][21] + signed_kernel[4][4] ~^ image[13][22];
assign xor_sum[9][19] = signed_kernel[0][0] ~^ image[9][19] + signed_kernel[0][1] ~^ image[9][20] + signed_kernel[0][2] ~^ image[9][21] + signed_kernel[0][3] ~^ image[9][22] + signed_kernel[0][4] ~^ image[9][23] + signed_kernel[1][0] ~^ image[10][19] + signed_kernel[1][1] ~^ image[10][20] + signed_kernel[1][2] ~^ image[10][21] + signed_kernel[1][3] ~^ image[10][22] + signed_kernel[1][4] ~^ image[10][23] + signed_kernel[2][0] ~^ image[11][19] + signed_kernel[2][1] ~^ image[11][20] + signed_kernel[2][2] ~^ image[11][21] + signed_kernel[2][3] ~^ image[11][22] + signed_kernel[2][4] ~^ image[11][23] + signed_kernel[3][0] ~^ image[12][19] + signed_kernel[3][1] ~^ image[12][20] + signed_kernel[3][2] ~^ image[12][21] + signed_kernel[3][3] ~^ image[12][22] + signed_kernel[3][4] ~^ image[12][23] + signed_kernel[4][0] ~^ image[13][19] + signed_kernel[4][1] ~^ image[13][20] + signed_kernel[4][2] ~^ image[13][21] + signed_kernel[4][3] ~^ image[13][22] + signed_kernel[4][4] ~^ image[13][23];
assign xor_sum[9][20] = signed_kernel[0][0] ~^ image[9][20] + signed_kernel[0][1] ~^ image[9][21] + signed_kernel[0][2] ~^ image[9][22] + signed_kernel[0][3] ~^ image[9][23] + signed_kernel[0][4] ~^ image[9][24] + signed_kernel[1][0] ~^ image[10][20] + signed_kernel[1][1] ~^ image[10][21] + signed_kernel[1][2] ~^ image[10][22] + signed_kernel[1][3] ~^ image[10][23] + signed_kernel[1][4] ~^ image[10][24] + signed_kernel[2][0] ~^ image[11][20] + signed_kernel[2][1] ~^ image[11][21] + signed_kernel[2][2] ~^ image[11][22] + signed_kernel[2][3] ~^ image[11][23] + signed_kernel[2][4] ~^ image[11][24] + signed_kernel[3][0] ~^ image[12][20] + signed_kernel[3][1] ~^ image[12][21] + signed_kernel[3][2] ~^ image[12][22] + signed_kernel[3][3] ~^ image[12][23] + signed_kernel[3][4] ~^ image[12][24] + signed_kernel[4][0] ~^ image[13][20] + signed_kernel[4][1] ~^ image[13][21] + signed_kernel[4][2] ~^ image[13][22] + signed_kernel[4][3] ~^ image[13][23] + signed_kernel[4][4] ~^ image[13][24];
assign xor_sum[9][21] = signed_kernel[0][0] ~^ image[9][21] + signed_kernel[0][1] ~^ image[9][22] + signed_kernel[0][2] ~^ image[9][23] + signed_kernel[0][3] ~^ image[9][24] + signed_kernel[0][4] ~^ image[9][25] + signed_kernel[1][0] ~^ image[10][21] + signed_kernel[1][1] ~^ image[10][22] + signed_kernel[1][2] ~^ image[10][23] + signed_kernel[1][3] ~^ image[10][24] + signed_kernel[1][4] ~^ image[10][25] + signed_kernel[2][0] ~^ image[11][21] + signed_kernel[2][1] ~^ image[11][22] + signed_kernel[2][2] ~^ image[11][23] + signed_kernel[2][3] ~^ image[11][24] + signed_kernel[2][4] ~^ image[11][25] + signed_kernel[3][0] ~^ image[12][21] + signed_kernel[3][1] ~^ image[12][22] + signed_kernel[3][2] ~^ image[12][23] + signed_kernel[3][3] ~^ image[12][24] + signed_kernel[3][4] ~^ image[12][25] + signed_kernel[4][0] ~^ image[13][21] + signed_kernel[4][1] ~^ image[13][22] + signed_kernel[4][2] ~^ image[13][23] + signed_kernel[4][3] ~^ image[13][24] + signed_kernel[4][4] ~^ image[13][25];
assign xor_sum[9][22] = signed_kernel[0][0] ~^ image[9][22] + signed_kernel[0][1] ~^ image[9][23] + signed_kernel[0][2] ~^ image[9][24] + signed_kernel[0][3] ~^ image[9][25] + signed_kernel[0][4] ~^ image[9][26] + signed_kernel[1][0] ~^ image[10][22] + signed_kernel[1][1] ~^ image[10][23] + signed_kernel[1][2] ~^ image[10][24] + signed_kernel[1][3] ~^ image[10][25] + signed_kernel[1][4] ~^ image[10][26] + signed_kernel[2][0] ~^ image[11][22] + signed_kernel[2][1] ~^ image[11][23] + signed_kernel[2][2] ~^ image[11][24] + signed_kernel[2][3] ~^ image[11][25] + signed_kernel[2][4] ~^ image[11][26] + signed_kernel[3][0] ~^ image[12][22] + signed_kernel[3][1] ~^ image[12][23] + signed_kernel[3][2] ~^ image[12][24] + signed_kernel[3][3] ~^ image[12][25] + signed_kernel[3][4] ~^ image[12][26] + signed_kernel[4][0] ~^ image[13][22] + signed_kernel[4][1] ~^ image[13][23] + signed_kernel[4][2] ~^ image[13][24] + signed_kernel[4][3] ~^ image[13][25] + signed_kernel[4][4] ~^ image[13][26];
assign xor_sum[9][23] = signed_kernel[0][0] ~^ image[9][23] + signed_kernel[0][1] ~^ image[9][24] + signed_kernel[0][2] ~^ image[9][25] + signed_kernel[0][3] ~^ image[9][26] + signed_kernel[0][4] ~^ image[9][27] + signed_kernel[1][0] ~^ image[10][23] + signed_kernel[1][1] ~^ image[10][24] + signed_kernel[1][2] ~^ image[10][25] + signed_kernel[1][3] ~^ image[10][26] + signed_kernel[1][4] ~^ image[10][27] + signed_kernel[2][0] ~^ image[11][23] + signed_kernel[2][1] ~^ image[11][24] + signed_kernel[2][2] ~^ image[11][25] + signed_kernel[2][3] ~^ image[11][26] + signed_kernel[2][4] ~^ image[11][27] + signed_kernel[3][0] ~^ image[12][23] + signed_kernel[3][1] ~^ image[12][24] + signed_kernel[3][2] ~^ image[12][25] + signed_kernel[3][3] ~^ image[12][26] + signed_kernel[3][4] ~^ image[12][27] + signed_kernel[4][0] ~^ image[13][23] + signed_kernel[4][1] ~^ image[13][24] + signed_kernel[4][2] ~^ image[13][25] + signed_kernel[4][3] ~^ image[13][26] + signed_kernel[4][4] ~^ image[13][27];
assign xor_sum[10][0] = signed_kernel[0][0] ~^ image[10][0] + signed_kernel[0][1] ~^ image[10][1] + signed_kernel[0][2] ~^ image[10][2] + signed_kernel[0][3] ~^ image[10][3] + signed_kernel[0][4] ~^ image[10][4] + signed_kernel[1][0] ~^ image[11][0] + signed_kernel[1][1] ~^ image[11][1] + signed_kernel[1][2] ~^ image[11][2] + signed_kernel[1][3] ~^ image[11][3] + signed_kernel[1][4] ~^ image[11][4] + signed_kernel[2][0] ~^ image[12][0] + signed_kernel[2][1] ~^ image[12][1] + signed_kernel[2][2] ~^ image[12][2] + signed_kernel[2][3] ~^ image[12][3] + signed_kernel[2][4] ~^ image[12][4] + signed_kernel[3][0] ~^ image[13][0] + signed_kernel[3][1] ~^ image[13][1] + signed_kernel[3][2] ~^ image[13][2] + signed_kernel[3][3] ~^ image[13][3] + signed_kernel[3][4] ~^ image[13][4] + signed_kernel[4][0] ~^ image[14][0] + signed_kernel[4][1] ~^ image[14][1] + signed_kernel[4][2] ~^ image[14][2] + signed_kernel[4][3] ~^ image[14][3] + signed_kernel[4][4] ~^ image[14][4];
assign xor_sum[10][1] = signed_kernel[0][0] ~^ image[10][1] + signed_kernel[0][1] ~^ image[10][2] + signed_kernel[0][2] ~^ image[10][3] + signed_kernel[0][3] ~^ image[10][4] + signed_kernel[0][4] ~^ image[10][5] + signed_kernel[1][0] ~^ image[11][1] + signed_kernel[1][1] ~^ image[11][2] + signed_kernel[1][2] ~^ image[11][3] + signed_kernel[1][3] ~^ image[11][4] + signed_kernel[1][4] ~^ image[11][5] + signed_kernel[2][0] ~^ image[12][1] + signed_kernel[2][1] ~^ image[12][2] + signed_kernel[2][2] ~^ image[12][3] + signed_kernel[2][3] ~^ image[12][4] + signed_kernel[2][4] ~^ image[12][5] + signed_kernel[3][0] ~^ image[13][1] + signed_kernel[3][1] ~^ image[13][2] + signed_kernel[3][2] ~^ image[13][3] + signed_kernel[3][3] ~^ image[13][4] + signed_kernel[3][4] ~^ image[13][5] + signed_kernel[4][0] ~^ image[14][1] + signed_kernel[4][1] ~^ image[14][2] + signed_kernel[4][2] ~^ image[14][3] + signed_kernel[4][3] ~^ image[14][4] + signed_kernel[4][4] ~^ image[14][5];
assign xor_sum[10][2] = signed_kernel[0][0] ~^ image[10][2] + signed_kernel[0][1] ~^ image[10][3] + signed_kernel[0][2] ~^ image[10][4] + signed_kernel[0][3] ~^ image[10][5] + signed_kernel[0][4] ~^ image[10][6] + signed_kernel[1][0] ~^ image[11][2] + signed_kernel[1][1] ~^ image[11][3] + signed_kernel[1][2] ~^ image[11][4] + signed_kernel[1][3] ~^ image[11][5] + signed_kernel[1][4] ~^ image[11][6] + signed_kernel[2][0] ~^ image[12][2] + signed_kernel[2][1] ~^ image[12][3] + signed_kernel[2][2] ~^ image[12][4] + signed_kernel[2][3] ~^ image[12][5] + signed_kernel[2][4] ~^ image[12][6] + signed_kernel[3][0] ~^ image[13][2] + signed_kernel[3][1] ~^ image[13][3] + signed_kernel[3][2] ~^ image[13][4] + signed_kernel[3][3] ~^ image[13][5] + signed_kernel[3][4] ~^ image[13][6] + signed_kernel[4][0] ~^ image[14][2] + signed_kernel[4][1] ~^ image[14][3] + signed_kernel[4][2] ~^ image[14][4] + signed_kernel[4][3] ~^ image[14][5] + signed_kernel[4][4] ~^ image[14][6];
assign xor_sum[10][3] = signed_kernel[0][0] ~^ image[10][3] + signed_kernel[0][1] ~^ image[10][4] + signed_kernel[0][2] ~^ image[10][5] + signed_kernel[0][3] ~^ image[10][6] + signed_kernel[0][4] ~^ image[10][7] + signed_kernel[1][0] ~^ image[11][3] + signed_kernel[1][1] ~^ image[11][4] + signed_kernel[1][2] ~^ image[11][5] + signed_kernel[1][3] ~^ image[11][6] + signed_kernel[1][4] ~^ image[11][7] + signed_kernel[2][0] ~^ image[12][3] + signed_kernel[2][1] ~^ image[12][4] + signed_kernel[2][2] ~^ image[12][5] + signed_kernel[2][3] ~^ image[12][6] + signed_kernel[2][4] ~^ image[12][7] + signed_kernel[3][0] ~^ image[13][3] + signed_kernel[3][1] ~^ image[13][4] + signed_kernel[3][2] ~^ image[13][5] + signed_kernel[3][3] ~^ image[13][6] + signed_kernel[3][4] ~^ image[13][7] + signed_kernel[4][0] ~^ image[14][3] + signed_kernel[4][1] ~^ image[14][4] + signed_kernel[4][2] ~^ image[14][5] + signed_kernel[4][3] ~^ image[14][6] + signed_kernel[4][4] ~^ image[14][7];
assign xor_sum[10][4] = signed_kernel[0][0] ~^ image[10][4] + signed_kernel[0][1] ~^ image[10][5] + signed_kernel[0][2] ~^ image[10][6] + signed_kernel[0][3] ~^ image[10][7] + signed_kernel[0][4] ~^ image[10][8] + signed_kernel[1][0] ~^ image[11][4] + signed_kernel[1][1] ~^ image[11][5] + signed_kernel[1][2] ~^ image[11][6] + signed_kernel[1][3] ~^ image[11][7] + signed_kernel[1][4] ~^ image[11][8] + signed_kernel[2][0] ~^ image[12][4] + signed_kernel[2][1] ~^ image[12][5] + signed_kernel[2][2] ~^ image[12][6] + signed_kernel[2][3] ~^ image[12][7] + signed_kernel[2][4] ~^ image[12][8] + signed_kernel[3][0] ~^ image[13][4] + signed_kernel[3][1] ~^ image[13][5] + signed_kernel[3][2] ~^ image[13][6] + signed_kernel[3][3] ~^ image[13][7] + signed_kernel[3][4] ~^ image[13][8] + signed_kernel[4][0] ~^ image[14][4] + signed_kernel[4][1] ~^ image[14][5] + signed_kernel[4][2] ~^ image[14][6] + signed_kernel[4][3] ~^ image[14][7] + signed_kernel[4][4] ~^ image[14][8];
assign xor_sum[10][5] = signed_kernel[0][0] ~^ image[10][5] + signed_kernel[0][1] ~^ image[10][6] + signed_kernel[0][2] ~^ image[10][7] + signed_kernel[0][3] ~^ image[10][8] + signed_kernel[0][4] ~^ image[10][9] + signed_kernel[1][0] ~^ image[11][5] + signed_kernel[1][1] ~^ image[11][6] + signed_kernel[1][2] ~^ image[11][7] + signed_kernel[1][3] ~^ image[11][8] + signed_kernel[1][4] ~^ image[11][9] + signed_kernel[2][0] ~^ image[12][5] + signed_kernel[2][1] ~^ image[12][6] + signed_kernel[2][2] ~^ image[12][7] + signed_kernel[2][3] ~^ image[12][8] + signed_kernel[2][4] ~^ image[12][9] + signed_kernel[3][0] ~^ image[13][5] + signed_kernel[3][1] ~^ image[13][6] + signed_kernel[3][2] ~^ image[13][7] + signed_kernel[3][3] ~^ image[13][8] + signed_kernel[3][4] ~^ image[13][9] + signed_kernel[4][0] ~^ image[14][5] + signed_kernel[4][1] ~^ image[14][6] + signed_kernel[4][2] ~^ image[14][7] + signed_kernel[4][3] ~^ image[14][8] + signed_kernel[4][4] ~^ image[14][9];
assign xor_sum[10][6] = signed_kernel[0][0] ~^ image[10][6] + signed_kernel[0][1] ~^ image[10][7] + signed_kernel[0][2] ~^ image[10][8] + signed_kernel[0][3] ~^ image[10][9] + signed_kernel[0][4] ~^ image[10][10] + signed_kernel[1][0] ~^ image[11][6] + signed_kernel[1][1] ~^ image[11][7] + signed_kernel[1][2] ~^ image[11][8] + signed_kernel[1][3] ~^ image[11][9] + signed_kernel[1][4] ~^ image[11][10] + signed_kernel[2][0] ~^ image[12][6] + signed_kernel[2][1] ~^ image[12][7] + signed_kernel[2][2] ~^ image[12][8] + signed_kernel[2][3] ~^ image[12][9] + signed_kernel[2][4] ~^ image[12][10] + signed_kernel[3][0] ~^ image[13][6] + signed_kernel[3][1] ~^ image[13][7] + signed_kernel[3][2] ~^ image[13][8] + signed_kernel[3][3] ~^ image[13][9] + signed_kernel[3][4] ~^ image[13][10] + signed_kernel[4][0] ~^ image[14][6] + signed_kernel[4][1] ~^ image[14][7] + signed_kernel[4][2] ~^ image[14][8] + signed_kernel[4][3] ~^ image[14][9] + signed_kernel[4][4] ~^ image[14][10];
assign xor_sum[10][7] = signed_kernel[0][0] ~^ image[10][7] + signed_kernel[0][1] ~^ image[10][8] + signed_kernel[0][2] ~^ image[10][9] + signed_kernel[0][3] ~^ image[10][10] + signed_kernel[0][4] ~^ image[10][11] + signed_kernel[1][0] ~^ image[11][7] + signed_kernel[1][1] ~^ image[11][8] + signed_kernel[1][2] ~^ image[11][9] + signed_kernel[1][3] ~^ image[11][10] + signed_kernel[1][4] ~^ image[11][11] + signed_kernel[2][0] ~^ image[12][7] + signed_kernel[2][1] ~^ image[12][8] + signed_kernel[2][2] ~^ image[12][9] + signed_kernel[2][3] ~^ image[12][10] + signed_kernel[2][4] ~^ image[12][11] + signed_kernel[3][0] ~^ image[13][7] + signed_kernel[3][1] ~^ image[13][8] + signed_kernel[3][2] ~^ image[13][9] + signed_kernel[3][3] ~^ image[13][10] + signed_kernel[3][4] ~^ image[13][11] + signed_kernel[4][0] ~^ image[14][7] + signed_kernel[4][1] ~^ image[14][8] + signed_kernel[4][2] ~^ image[14][9] + signed_kernel[4][3] ~^ image[14][10] + signed_kernel[4][4] ~^ image[14][11];
assign xor_sum[10][8] = signed_kernel[0][0] ~^ image[10][8] + signed_kernel[0][1] ~^ image[10][9] + signed_kernel[0][2] ~^ image[10][10] + signed_kernel[0][3] ~^ image[10][11] + signed_kernel[0][4] ~^ image[10][12] + signed_kernel[1][0] ~^ image[11][8] + signed_kernel[1][1] ~^ image[11][9] + signed_kernel[1][2] ~^ image[11][10] + signed_kernel[1][3] ~^ image[11][11] + signed_kernel[1][4] ~^ image[11][12] + signed_kernel[2][0] ~^ image[12][8] + signed_kernel[2][1] ~^ image[12][9] + signed_kernel[2][2] ~^ image[12][10] + signed_kernel[2][3] ~^ image[12][11] + signed_kernel[2][4] ~^ image[12][12] + signed_kernel[3][0] ~^ image[13][8] + signed_kernel[3][1] ~^ image[13][9] + signed_kernel[3][2] ~^ image[13][10] + signed_kernel[3][3] ~^ image[13][11] + signed_kernel[3][4] ~^ image[13][12] + signed_kernel[4][0] ~^ image[14][8] + signed_kernel[4][1] ~^ image[14][9] + signed_kernel[4][2] ~^ image[14][10] + signed_kernel[4][3] ~^ image[14][11] + signed_kernel[4][4] ~^ image[14][12];
assign xor_sum[10][9] = signed_kernel[0][0] ~^ image[10][9] + signed_kernel[0][1] ~^ image[10][10] + signed_kernel[0][2] ~^ image[10][11] + signed_kernel[0][3] ~^ image[10][12] + signed_kernel[0][4] ~^ image[10][13] + signed_kernel[1][0] ~^ image[11][9] + signed_kernel[1][1] ~^ image[11][10] + signed_kernel[1][2] ~^ image[11][11] + signed_kernel[1][3] ~^ image[11][12] + signed_kernel[1][4] ~^ image[11][13] + signed_kernel[2][0] ~^ image[12][9] + signed_kernel[2][1] ~^ image[12][10] + signed_kernel[2][2] ~^ image[12][11] + signed_kernel[2][3] ~^ image[12][12] + signed_kernel[2][4] ~^ image[12][13] + signed_kernel[3][0] ~^ image[13][9] + signed_kernel[3][1] ~^ image[13][10] + signed_kernel[3][2] ~^ image[13][11] + signed_kernel[3][3] ~^ image[13][12] + signed_kernel[3][4] ~^ image[13][13] + signed_kernel[4][0] ~^ image[14][9] + signed_kernel[4][1] ~^ image[14][10] + signed_kernel[4][2] ~^ image[14][11] + signed_kernel[4][3] ~^ image[14][12] + signed_kernel[4][4] ~^ image[14][13];
assign xor_sum[10][10] = signed_kernel[0][0] ~^ image[10][10] + signed_kernel[0][1] ~^ image[10][11] + signed_kernel[0][2] ~^ image[10][12] + signed_kernel[0][3] ~^ image[10][13] + signed_kernel[0][4] ~^ image[10][14] + signed_kernel[1][0] ~^ image[11][10] + signed_kernel[1][1] ~^ image[11][11] + signed_kernel[1][2] ~^ image[11][12] + signed_kernel[1][3] ~^ image[11][13] + signed_kernel[1][4] ~^ image[11][14] + signed_kernel[2][0] ~^ image[12][10] + signed_kernel[2][1] ~^ image[12][11] + signed_kernel[2][2] ~^ image[12][12] + signed_kernel[2][3] ~^ image[12][13] + signed_kernel[2][4] ~^ image[12][14] + signed_kernel[3][0] ~^ image[13][10] + signed_kernel[3][1] ~^ image[13][11] + signed_kernel[3][2] ~^ image[13][12] + signed_kernel[3][3] ~^ image[13][13] + signed_kernel[3][4] ~^ image[13][14] + signed_kernel[4][0] ~^ image[14][10] + signed_kernel[4][1] ~^ image[14][11] + signed_kernel[4][2] ~^ image[14][12] + signed_kernel[4][3] ~^ image[14][13] + signed_kernel[4][4] ~^ image[14][14];
assign xor_sum[10][11] = signed_kernel[0][0] ~^ image[10][11] + signed_kernel[0][1] ~^ image[10][12] + signed_kernel[0][2] ~^ image[10][13] + signed_kernel[0][3] ~^ image[10][14] + signed_kernel[0][4] ~^ image[10][15] + signed_kernel[1][0] ~^ image[11][11] + signed_kernel[1][1] ~^ image[11][12] + signed_kernel[1][2] ~^ image[11][13] + signed_kernel[1][3] ~^ image[11][14] + signed_kernel[1][4] ~^ image[11][15] + signed_kernel[2][0] ~^ image[12][11] + signed_kernel[2][1] ~^ image[12][12] + signed_kernel[2][2] ~^ image[12][13] + signed_kernel[2][3] ~^ image[12][14] + signed_kernel[2][4] ~^ image[12][15] + signed_kernel[3][0] ~^ image[13][11] + signed_kernel[3][1] ~^ image[13][12] + signed_kernel[3][2] ~^ image[13][13] + signed_kernel[3][3] ~^ image[13][14] + signed_kernel[3][4] ~^ image[13][15] + signed_kernel[4][0] ~^ image[14][11] + signed_kernel[4][1] ~^ image[14][12] + signed_kernel[4][2] ~^ image[14][13] + signed_kernel[4][3] ~^ image[14][14] + signed_kernel[4][4] ~^ image[14][15];
assign xor_sum[10][12] = signed_kernel[0][0] ~^ image[10][12] + signed_kernel[0][1] ~^ image[10][13] + signed_kernel[0][2] ~^ image[10][14] + signed_kernel[0][3] ~^ image[10][15] + signed_kernel[0][4] ~^ image[10][16] + signed_kernel[1][0] ~^ image[11][12] + signed_kernel[1][1] ~^ image[11][13] + signed_kernel[1][2] ~^ image[11][14] + signed_kernel[1][3] ~^ image[11][15] + signed_kernel[1][4] ~^ image[11][16] + signed_kernel[2][0] ~^ image[12][12] + signed_kernel[2][1] ~^ image[12][13] + signed_kernel[2][2] ~^ image[12][14] + signed_kernel[2][3] ~^ image[12][15] + signed_kernel[2][4] ~^ image[12][16] + signed_kernel[3][0] ~^ image[13][12] + signed_kernel[3][1] ~^ image[13][13] + signed_kernel[3][2] ~^ image[13][14] + signed_kernel[3][3] ~^ image[13][15] + signed_kernel[3][4] ~^ image[13][16] + signed_kernel[4][0] ~^ image[14][12] + signed_kernel[4][1] ~^ image[14][13] + signed_kernel[4][2] ~^ image[14][14] + signed_kernel[4][3] ~^ image[14][15] + signed_kernel[4][4] ~^ image[14][16];
assign xor_sum[10][13] = signed_kernel[0][0] ~^ image[10][13] + signed_kernel[0][1] ~^ image[10][14] + signed_kernel[0][2] ~^ image[10][15] + signed_kernel[0][3] ~^ image[10][16] + signed_kernel[0][4] ~^ image[10][17] + signed_kernel[1][0] ~^ image[11][13] + signed_kernel[1][1] ~^ image[11][14] + signed_kernel[1][2] ~^ image[11][15] + signed_kernel[1][3] ~^ image[11][16] + signed_kernel[1][4] ~^ image[11][17] + signed_kernel[2][0] ~^ image[12][13] + signed_kernel[2][1] ~^ image[12][14] + signed_kernel[2][2] ~^ image[12][15] + signed_kernel[2][3] ~^ image[12][16] + signed_kernel[2][4] ~^ image[12][17] + signed_kernel[3][0] ~^ image[13][13] + signed_kernel[3][1] ~^ image[13][14] + signed_kernel[3][2] ~^ image[13][15] + signed_kernel[3][3] ~^ image[13][16] + signed_kernel[3][4] ~^ image[13][17] + signed_kernel[4][0] ~^ image[14][13] + signed_kernel[4][1] ~^ image[14][14] + signed_kernel[4][2] ~^ image[14][15] + signed_kernel[4][3] ~^ image[14][16] + signed_kernel[4][4] ~^ image[14][17];
assign xor_sum[10][14] = signed_kernel[0][0] ~^ image[10][14] + signed_kernel[0][1] ~^ image[10][15] + signed_kernel[0][2] ~^ image[10][16] + signed_kernel[0][3] ~^ image[10][17] + signed_kernel[0][4] ~^ image[10][18] + signed_kernel[1][0] ~^ image[11][14] + signed_kernel[1][1] ~^ image[11][15] + signed_kernel[1][2] ~^ image[11][16] + signed_kernel[1][3] ~^ image[11][17] + signed_kernel[1][4] ~^ image[11][18] + signed_kernel[2][0] ~^ image[12][14] + signed_kernel[2][1] ~^ image[12][15] + signed_kernel[2][2] ~^ image[12][16] + signed_kernel[2][3] ~^ image[12][17] + signed_kernel[2][4] ~^ image[12][18] + signed_kernel[3][0] ~^ image[13][14] + signed_kernel[3][1] ~^ image[13][15] + signed_kernel[3][2] ~^ image[13][16] + signed_kernel[3][3] ~^ image[13][17] + signed_kernel[3][4] ~^ image[13][18] + signed_kernel[4][0] ~^ image[14][14] + signed_kernel[4][1] ~^ image[14][15] + signed_kernel[4][2] ~^ image[14][16] + signed_kernel[4][3] ~^ image[14][17] + signed_kernel[4][4] ~^ image[14][18];
assign xor_sum[10][15] = signed_kernel[0][0] ~^ image[10][15] + signed_kernel[0][1] ~^ image[10][16] + signed_kernel[0][2] ~^ image[10][17] + signed_kernel[0][3] ~^ image[10][18] + signed_kernel[0][4] ~^ image[10][19] + signed_kernel[1][0] ~^ image[11][15] + signed_kernel[1][1] ~^ image[11][16] + signed_kernel[1][2] ~^ image[11][17] + signed_kernel[1][3] ~^ image[11][18] + signed_kernel[1][4] ~^ image[11][19] + signed_kernel[2][0] ~^ image[12][15] + signed_kernel[2][1] ~^ image[12][16] + signed_kernel[2][2] ~^ image[12][17] + signed_kernel[2][3] ~^ image[12][18] + signed_kernel[2][4] ~^ image[12][19] + signed_kernel[3][0] ~^ image[13][15] + signed_kernel[3][1] ~^ image[13][16] + signed_kernel[3][2] ~^ image[13][17] + signed_kernel[3][3] ~^ image[13][18] + signed_kernel[3][4] ~^ image[13][19] + signed_kernel[4][0] ~^ image[14][15] + signed_kernel[4][1] ~^ image[14][16] + signed_kernel[4][2] ~^ image[14][17] + signed_kernel[4][3] ~^ image[14][18] + signed_kernel[4][4] ~^ image[14][19];
assign xor_sum[10][16] = signed_kernel[0][0] ~^ image[10][16] + signed_kernel[0][1] ~^ image[10][17] + signed_kernel[0][2] ~^ image[10][18] + signed_kernel[0][3] ~^ image[10][19] + signed_kernel[0][4] ~^ image[10][20] + signed_kernel[1][0] ~^ image[11][16] + signed_kernel[1][1] ~^ image[11][17] + signed_kernel[1][2] ~^ image[11][18] + signed_kernel[1][3] ~^ image[11][19] + signed_kernel[1][4] ~^ image[11][20] + signed_kernel[2][0] ~^ image[12][16] + signed_kernel[2][1] ~^ image[12][17] + signed_kernel[2][2] ~^ image[12][18] + signed_kernel[2][3] ~^ image[12][19] + signed_kernel[2][4] ~^ image[12][20] + signed_kernel[3][0] ~^ image[13][16] + signed_kernel[3][1] ~^ image[13][17] + signed_kernel[3][2] ~^ image[13][18] + signed_kernel[3][3] ~^ image[13][19] + signed_kernel[3][4] ~^ image[13][20] + signed_kernel[4][0] ~^ image[14][16] + signed_kernel[4][1] ~^ image[14][17] + signed_kernel[4][2] ~^ image[14][18] + signed_kernel[4][3] ~^ image[14][19] + signed_kernel[4][4] ~^ image[14][20];
assign xor_sum[10][17] = signed_kernel[0][0] ~^ image[10][17] + signed_kernel[0][1] ~^ image[10][18] + signed_kernel[0][2] ~^ image[10][19] + signed_kernel[0][3] ~^ image[10][20] + signed_kernel[0][4] ~^ image[10][21] + signed_kernel[1][0] ~^ image[11][17] + signed_kernel[1][1] ~^ image[11][18] + signed_kernel[1][2] ~^ image[11][19] + signed_kernel[1][3] ~^ image[11][20] + signed_kernel[1][4] ~^ image[11][21] + signed_kernel[2][0] ~^ image[12][17] + signed_kernel[2][1] ~^ image[12][18] + signed_kernel[2][2] ~^ image[12][19] + signed_kernel[2][3] ~^ image[12][20] + signed_kernel[2][4] ~^ image[12][21] + signed_kernel[3][0] ~^ image[13][17] + signed_kernel[3][1] ~^ image[13][18] + signed_kernel[3][2] ~^ image[13][19] + signed_kernel[3][3] ~^ image[13][20] + signed_kernel[3][4] ~^ image[13][21] + signed_kernel[4][0] ~^ image[14][17] + signed_kernel[4][1] ~^ image[14][18] + signed_kernel[4][2] ~^ image[14][19] + signed_kernel[4][3] ~^ image[14][20] + signed_kernel[4][4] ~^ image[14][21];
assign xor_sum[10][18] = signed_kernel[0][0] ~^ image[10][18] + signed_kernel[0][1] ~^ image[10][19] + signed_kernel[0][2] ~^ image[10][20] + signed_kernel[0][3] ~^ image[10][21] + signed_kernel[0][4] ~^ image[10][22] + signed_kernel[1][0] ~^ image[11][18] + signed_kernel[1][1] ~^ image[11][19] + signed_kernel[1][2] ~^ image[11][20] + signed_kernel[1][3] ~^ image[11][21] + signed_kernel[1][4] ~^ image[11][22] + signed_kernel[2][0] ~^ image[12][18] + signed_kernel[2][1] ~^ image[12][19] + signed_kernel[2][2] ~^ image[12][20] + signed_kernel[2][3] ~^ image[12][21] + signed_kernel[2][4] ~^ image[12][22] + signed_kernel[3][0] ~^ image[13][18] + signed_kernel[3][1] ~^ image[13][19] + signed_kernel[3][2] ~^ image[13][20] + signed_kernel[3][3] ~^ image[13][21] + signed_kernel[3][4] ~^ image[13][22] + signed_kernel[4][0] ~^ image[14][18] + signed_kernel[4][1] ~^ image[14][19] + signed_kernel[4][2] ~^ image[14][20] + signed_kernel[4][3] ~^ image[14][21] + signed_kernel[4][4] ~^ image[14][22];
assign xor_sum[10][19] = signed_kernel[0][0] ~^ image[10][19] + signed_kernel[0][1] ~^ image[10][20] + signed_kernel[0][2] ~^ image[10][21] + signed_kernel[0][3] ~^ image[10][22] + signed_kernel[0][4] ~^ image[10][23] + signed_kernel[1][0] ~^ image[11][19] + signed_kernel[1][1] ~^ image[11][20] + signed_kernel[1][2] ~^ image[11][21] + signed_kernel[1][3] ~^ image[11][22] + signed_kernel[1][4] ~^ image[11][23] + signed_kernel[2][0] ~^ image[12][19] + signed_kernel[2][1] ~^ image[12][20] + signed_kernel[2][2] ~^ image[12][21] + signed_kernel[2][3] ~^ image[12][22] + signed_kernel[2][4] ~^ image[12][23] + signed_kernel[3][0] ~^ image[13][19] + signed_kernel[3][1] ~^ image[13][20] + signed_kernel[3][2] ~^ image[13][21] + signed_kernel[3][3] ~^ image[13][22] + signed_kernel[3][4] ~^ image[13][23] + signed_kernel[4][0] ~^ image[14][19] + signed_kernel[4][1] ~^ image[14][20] + signed_kernel[4][2] ~^ image[14][21] + signed_kernel[4][3] ~^ image[14][22] + signed_kernel[4][4] ~^ image[14][23];
assign xor_sum[10][20] = signed_kernel[0][0] ~^ image[10][20] + signed_kernel[0][1] ~^ image[10][21] + signed_kernel[0][2] ~^ image[10][22] + signed_kernel[0][3] ~^ image[10][23] + signed_kernel[0][4] ~^ image[10][24] + signed_kernel[1][0] ~^ image[11][20] + signed_kernel[1][1] ~^ image[11][21] + signed_kernel[1][2] ~^ image[11][22] + signed_kernel[1][3] ~^ image[11][23] + signed_kernel[1][4] ~^ image[11][24] + signed_kernel[2][0] ~^ image[12][20] + signed_kernel[2][1] ~^ image[12][21] + signed_kernel[2][2] ~^ image[12][22] + signed_kernel[2][3] ~^ image[12][23] + signed_kernel[2][4] ~^ image[12][24] + signed_kernel[3][0] ~^ image[13][20] + signed_kernel[3][1] ~^ image[13][21] + signed_kernel[3][2] ~^ image[13][22] + signed_kernel[3][3] ~^ image[13][23] + signed_kernel[3][4] ~^ image[13][24] + signed_kernel[4][0] ~^ image[14][20] + signed_kernel[4][1] ~^ image[14][21] + signed_kernel[4][2] ~^ image[14][22] + signed_kernel[4][3] ~^ image[14][23] + signed_kernel[4][4] ~^ image[14][24];
assign xor_sum[10][21] = signed_kernel[0][0] ~^ image[10][21] + signed_kernel[0][1] ~^ image[10][22] + signed_kernel[0][2] ~^ image[10][23] + signed_kernel[0][3] ~^ image[10][24] + signed_kernel[0][4] ~^ image[10][25] + signed_kernel[1][0] ~^ image[11][21] + signed_kernel[1][1] ~^ image[11][22] + signed_kernel[1][2] ~^ image[11][23] + signed_kernel[1][3] ~^ image[11][24] + signed_kernel[1][4] ~^ image[11][25] + signed_kernel[2][0] ~^ image[12][21] + signed_kernel[2][1] ~^ image[12][22] + signed_kernel[2][2] ~^ image[12][23] + signed_kernel[2][3] ~^ image[12][24] + signed_kernel[2][4] ~^ image[12][25] + signed_kernel[3][0] ~^ image[13][21] + signed_kernel[3][1] ~^ image[13][22] + signed_kernel[3][2] ~^ image[13][23] + signed_kernel[3][3] ~^ image[13][24] + signed_kernel[3][4] ~^ image[13][25] + signed_kernel[4][0] ~^ image[14][21] + signed_kernel[4][1] ~^ image[14][22] + signed_kernel[4][2] ~^ image[14][23] + signed_kernel[4][3] ~^ image[14][24] + signed_kernel[4][4] ~^ image[14][25];
assign xor_sum[10][22] = signed_kernel[0][0] ~^ image[10][22] + signed_kernel[0][1] ~^ image[10][23] + signed_kernel[0][2] ~^ image[10][24] + signed_kernel[0][3] ~^ image[10][25] + signed_kernel[0][4] ~^ image[10][26] + signed_kernel[1][0] ~^ image[11][22] + signed_kernel[1][1] ~^ image[11][23] + signed_kernel[1][2] ~^ image[11][24] + signed_kernel[1][3] ~^ image[11][25] + signed_kernel[1][4] ~^ image[11][26] + signed_kernel[2][0] ~^ image[12][22] + signed_kernel[2][1] ~^ image[12][23] + signed_kernel[2][2] ~^ image[12][24] + signed_kernel[2][3] ~^ image[12][25] + signed_kernel[2][4] ~^ image[12][26] + signed_kernel[3][0] ~^ image[13][22] + signed_kernel[3][1] ~^ image[13][23] + signed_kernel[3][2] ~^ image[13][24] + signed_kernel[3][3] ~^ image[13][25] + signed_kernel[3][4] ~^ image[13][26] + signed_kernel[4][0] ~^ image[14][22] + signed_kernel[4][1] ~^ image[14][23] + signed_kernel[4][2] ~^ image[14][24] + signed_kernel[4][3] ~^ image[14][25] + signed_kernel[4][4] ~^ image[14][26];
assign xor_sum[10][23] = signed_kernel[0][0] ~^ image[10][23] + signed_kernel[0][1] ~^ image[10][24] + signed_kernel[0][2] ~^ image[10][25] + signed_kernel[0][3] ~^ image[10][26] + signed_kernel[0][4] ~^ image[10][27] + signed_kernel[1][0] ~^ image[11][23] + signed_kernel[1][1] ~^ image[11][24] + signed_kernel[1][2] ~^ image[11][25] + signed_kernel[1][3] ~^ image[11][26] + signed_kernel[1][4] ~^ image[11][27] + signed_kernel[2][0] ~^ image[12][23] + signed_kernel[2][1] ~^ image[12][24] + signed_kernel[2][2] ~^ image[12][25] + signed_kernel[2][3] ~^ image[12][26] + signed_kernel[2][4] ~^ image[12][27] + signed_kernel[3][0] ~^ image[13][23] + signed_kernel[3][1] ~^ image[13][24] + signed_kernel[3][2] ~^ image[13][25] + signed_kernel[3][3] ~^ image[13][26] + signed_kernel[3][4] ~^ image[13][27] + signed_kernel[4][0] ~^ image[14][23] + signed_kernel[4][1] ~^ image[14][24] + signed_kernel[4][2] ~^ image[14][25] + signed_kernel[4][3] ~^ image[14][26] + signed_kernel[4][4] ~^ image[14][27];
assign xor_sum[11][0] = signed_kernel[0][0] ~^ image[11][0] + signed_kernel[0][1] ~^ image[11][1] + signed_kernel[0][2] ~^ image[11][2] + signed_kernel[0][3] ~^ image[11][3] + signed_kernel[0][4] ~^ image[11][4] + signed_kernel[1][0] ~^ image[12][0] + signed_kernel[1][1] ~^ image[12][1] + signed_kernel[1][2] ~^ image[12][2] + signed_kernel[1][3] ~^ image[12][3] + signed_kernel[1][4] ~^ image[12][4] + signed_kernel[2][0] ~^ image[13][0] + signed_kernel[2][1] ~^ image[13][1] + signed_kernel[2][2] ~^ image[13][2] + signed_kernel[2][3] ~^ image[13][3] + signed_kernel[2][4] ~^ image[13][4] + signed_kernel[3][0] ~^ image[14][0] + signed_kernel[3][1] ~^ image[14][1] + signed_kernel[3][2] ~^ image[14][2] + signed_kernel[3][3] ~^ image[14][3] + signed_kernel[3][4] ~^ image[14][4] + signed_kernel[4][0] ~^ image[15][0] + signed_kernel[4][1] ~^ image[15][1] + signed_kernel[4][2] ~^ image[15][2] + signed_kernel[4][3] ~^ image[15][3] + signed_kernel[4][4] ~^ image[15][4];
assign xor_sum[11][1] = signed_kernel[0][0] ~^ image[11][1] + signed_kernel[0][1] ~^ image[11][2] + signed_kernel[0][2] ~^ image[11][3] + signed_kernel[0][3] ~^ image[11][4] + signed_kernel[0][4] ~^ image[11][5] + signed_kernel[1][0] ~^ image[12][1] + signed_kernel[1][1] ~^ image[12][2] + signed_kernel[1][2] ~^ image[12][3] + signed_kernel[1][3] ~^ image[12][4] + signed_kernel[1][4] ~^ image[12][5] + signed_kernel[2][0] ~^ image[13][1] + signed_kernel[2][1] ~^ image[13][2] + signed_kernel[2][2] ~^ image[13][3] + signed_kernel[2][3] ~^ image[13][4] + signed_kernel[2][4] ~^ image[13][5] + signed_kernel[3][0] ~^ image[14][1] + signed_kernel[3][1] ~^ image[14][2] + signed_kernel[3][2] ~^ image[14][3] + signed_kernel[3][3] ~^ image[14][4] + signed_kernel[3][4] ~^ image[14][5] + signed_kernel[4][0] ~^ image[15][1] + signed_kernel[4][1] ~^ image[15][2] + signed_kernel[4][2] ~^ image[15][3] + signed_kernel[4][3] ~^ image[15][4] + signed_kernel[4][4] ~^ image[15][5];
assign xor_sum[11][2] = signed_kernel[0][0] ~^ image[11][2] + signed_kernel[0][1] ~^ image[11][3] + signed_kernel[0][2] ~^ image[11][4] + signed_kernel[0][3] ~^ image[11][5] + signed_kernel[0][4] ~^ image[11][6] + signed_kernel[1][0] ~^ image[12][2] + signed_kernel[1][1] ~^ image[12][3] + signed_kernel[1][2] ~^ image[12][4] + signed_kernel[1][3] ~^ image[12][5] + signed_kernel[1][4] ~^ image[12][6] + signed_kernel[2][0] ~^ image[13][2] + signed_kernel[2][1] ~^ image[13][3] + signed_kernel[2][2] ~^ image[13][4] + signed_kernel[2][3] ~^ image[13][5] + signed_kernel[2][4] ~^ image[13][6] + signed_kernel[3][0] ~^ image[14][2] + signed_kernel[3][1] ~^ image[14][3] + signed_kernel[3][2] ~^ image[14][4] + signed_kernel[3][3] ~^ image[14][5] + signed_kernel[3][4] ~^ image[14][6] + signed_kernel[4][0] ~^ image[15][2] + signed_kernel[4][1] ~^ image[15][3] + signed_kernel[4][2] ~^ image[15][4] + signed_kernel[4][3] ~^ image[15][5] + signed_kernel[4][4] ~^ image[15][6];
assign xor_sum[11][3] = signed_kernel[0][0] ~^ image[11][3] + signed_kernel[0][1] ~^ image[11][4] + signed_kernel[0][2] ~^ image[11][5] + signed_kernel[0][3] ~^ image[11][6] + signed_kernel[0][4] ~^ image[11][7] + signed_kernel[1][0] ~^ image[12][3] + signed_kernel[1][1] ~^ image[12][4] + signed_kernel[1][2] ~^ image[12][5] + signed_kernel[1][3] ~^ image[12][6] + signed_kernel[1][4] ~^ image[12][7] + signed_kernel[2][0] ~^ image[13][3] + signed_kernel[2][1] ~^ image[13][4] + signed_kernel[2][2] ~^ image[13][5] + signed_kernel[2][3] ~^ image[13][6] + signed_kernel[2][4] ~^ image[13][7] + signed_kernel[3][0] ~^ image[14][3] + signed_kernel[3][1] ~^ image[14][4] + signed_kernel[3][2] ~^ image[14][5] + signed_kernel[3][3] ~^ image[14][6] + signed_kernel[3][4] ~^ image[14][7] + signed_kernel[4][0] ~^ image[15][3] + signed_kernel[4][1] ~^ image[15][4] + signed_kernel[4][2] ~^ image[15][5] + signed_kernel[4][3] ~^ image[15][6] + signed_kernel[4][4] ~^ image[15][7];
assign xor_sum[11][4] = signed_kernel[0][0] ~^ image[11][4] + signed_kernel[0][1] ~^ image[11][5] + signed_kernel[0][2] ~^ image[11][6] + signed_kernel[0][3] ~^ image[11][7] + signed_kernel[0][4] ~^ image[11][8] + signed_kernel[1][0] ~^ image[12][4] + signed_kernel[1][1] ~^ image[12][5] + signed_kernel[1][2] ~^ image[12][6] + signed_kernel[1][3] ~^ image[12][7] + signed_kernel[1][4] ~^ image[12][8] + signed_kernel[2][0] ~^ image[13][4] + signed_kernel[2][1] ~^ image[13][5] + signed_kernel[2][2] ~^ image[13][6] + signed_kernel[2][3] ~^ image[13][7] + signed_kernel[2][4] ~^ image[13][8] + signed_kernel[3][0] ~^ image[14][4] + signed_kernel[3][1] ~^ image[14][5] + signed_kernel[3][2] ~^ image[14][6] + signed_kernel[3][3] ~^ image[14][7] + signed_kernel[3][4] ~^ image[14][8] + signed_kernel[4][0] ~^ image[15][4] + signed_kernel[4][1] ~^ image[15][5] + signed_kernel[4][2] ~^ image[15][6] + signed_kernel[4][3] ~^ image[15][7] + signed_kernel[4][4] ~^ image[15][8];
assign xor_sum[11][5] = signed_kernel[0][0] ~^ image[11][5] + signed_kernel[0][1] ~^ image[11][6] + signed_kernel[0][2] ~^ image[11][7] + signed_kernel[0][3] ~^ image[11][8] + signed_kernel[0][4] ~^ image[11][9] + signed_kernel[1][0] ~^ image[12][5] + signed_kernel[1][1] ~^ image[12][6] + signed_kernel[1][2] ~^ image[12][7] + signed_kernel[1][3] ~^ image[12][8] + signed_kernel[1][4] ~^ image[12][9] + signed_kernel[2][0] ~^ image[13][5] + signed_kernel[2][1] ~^ image[13][6] + signed_kernel[2][2] ~^ image[13][7] + signed_kernel[2][3] ~^ image[13][8] + signed_kernel[2][4] ~^ image[13][9] + signed_kernel[3][0] ~^ image[14][5] + signed_kernel[3][1] ~^ image[14][6] + signed_kernel[3][2] ~^ image[14][7] + signed_kernel[3][3] ~^ image[14][8] + signed_kernel[3][4] ~^ image[14][9] + signed_kernel[4][0] ~^ image[15][5] + signed_kernel[4][1] ~^ image[15][6] + signed_kernel[4][2] ~^ image[15][7] + signed_kernel[4][3] ~^ image[15][8] + signed_kernel[4][4] ~^ image[15][9];
assign xor_sum[11][6] = signed_kernel[0][0] ~^ image[11][6] + signed_kernel[0][1] ~^ image[11][7] + signed_kernel[0][2] ~^ image[11][8] + signed_kernel[0][3] ~^ image[11][9] + signed_kernel[0][4] ~^ image[11][10] + signed_kernel[1][0] ~^ image[12][6] + signed_kernel[1][1] ~^ image[12][7] + signed_kernel[1][2] ~^ image[12][8] + signed_kernel[1][3] ~^ image[12][9] + signed_kernel[1][4] ~^ image[12][10] + signed_kernel[2][0] ~^ image[13][6] + signed_kernel[2][1] ~^ image[13][7] + signed_kernel[2][2] ~^ image[13][8] + signed_kernel[2][3] ~^ image[13][9] + signed_kernel[2][4] ~^ image[13][10] + signed_kernel[3][0] ~^ image[14][6] + signed_kernel[3][1] ~^ image[14][7] + signed_kernel[3][2] ~^ image[14][8] + signed_kernel[3][3] ~^ image[14][9] + signed_kernel[3][4] ~^ image[14][10] + signed_kernel[4][0] ~^ image[15][6] + signed_kernel[4][1] ~^ image[15][7] + signed_kernel[4][2] ~^ image[15][8] + signed_kernel[4][3] ~^ image[15][9] + signed_kernel[4][4] ~^ image[15][10];
assign xor_sum[11][7] = signed_kernel[0][0] ~^ image[11][7] + signed_kernel[0][1] ~^ image[11][8] + signed_kernel[0][2] ~^ image[11][9] + signed_kernel[0][3] ~^ image[11][10] + signed_kernel[0][4] ~^ image[11][11] + signed_kernel[1][0] ~^ image[12][7] + signed_kernel[1][1] ~^ image[12][8] + signed_kernel[1][2] ~^ image[12][9] + signed_kernel[1][3] ~^ image[12][10] + signed_kernel[1][4] ~^ image[12][11] + signed_kernel[2][0] ~^ image[13][7] + signed_kernel[2][1] ~^ image[13][8] + signed_kernel[2][2] ~^ image[13][9] + signed_kernel[2][3] ~^ image[13][10] + signed_kernel[2][4] ~^ image[13][11] + signed_kernel[3][0] ~^ image[14][7] + signed_kernel[3][1] ~^ image[14][8] + signed_kernel[3][2] ~^ image[14][9] + signed_kernel[3][3] ~^ image[14][10] + signed_kernel[3][4] ~^ image[14][11] + signed_kernel[4][0] ~^ image[15][7] + signed_kernel[4][1] ~^ image[15][8] + signed_kernel[4][2] ~^ image[15][9] + signed_kernel[4][3] ~^ image[15][10] + signed_kernel[4][4] ~^ image[15][11];
assign xor_sum[11][8] = signed_kernel[0][0] ~^ image[11][8] + signed_kernel[0][1] ~^ image[11][9] + signed_kernel[0][2] ~^ image[11][10] + signed_kernel[0][3] ~^ image[11][11] + signed_kernel[0][4] ~^ image[11][12] + signed_kernel[1][0] ~^ image[12][8] + signed_kernel[1][1] ~^ image[12][9] + signed_kernel[1][2] ~^ image[12][10] + signed_kernel[1][3] ~^ image[12][11] + signed_kernel[1][4] ~^ image[12][12] + signed_kernel[2][0] ~^ image[13][8] + signed_kernel[2][1] ~^ image[13][9] + signed_kernel[2][2] ~^ image[13][10] + signed_kernel[2][3] ~^ image[13][11] + signed_kernel[2][4] ~^ image[13][12] + signed_kernel[3][0] ~^ image[14][8] + signed_kernel[3][1] ~^ image[14][9] + signed_kernel[3][2] ~^ image[14][10] + signed_kernel[3][3] ~^ image[14][11] + signed_kernel[3][4] ~^ image[14][12] + signed_kernel[4][0] ~^ image[15][8] + signed_kernel[4][1] ~^ image[15][9] + signed_kernel[4][2] ~^ image[15][10] + signed_kernel[4][3] ~^ image[15][11] + signed_kernel[4][4] ~^ image[15][12];
assign xor_sum[11][9] = signed_kernel[0][0] ~^ image[11][9] + signed_kernel[0][1] ~^ image[11][10] + signed_kernel[0][2] ~^ image[11][11] + signed_kernel[0][3] ~^ image[11][12] + signed_kernel[0][4] ~^ image[11][13] + signed_kernel[1][0] ~^ image[12][9] + signed_kernel[1][1] ~^ image[12][10] + signed_kernel[1][2] ~^ image[12][11] + signed_kernel[1][3] ~^ image[12][12] + signed_kernel[1][4] ~^ image[12][13] + signed_kernel[2][0] ~^ image[13][9] + signed_kernel[2][1] ~^ image[13][10] + signed_kernel[2][2] ~^ image[13][11] + signed_kernel[2][3] ~^ image[13][12] + signed_kernel[2][4] ~^ image[13][13] + signed_kernel[3][0] ~^ image[14][9] + signed_kernel[3][1] ~^ image[14][10] + signed_kernel[3][2] ~^ image[14][11] + signed_kernel[3][3] ~^ image[14][12] + signed_kernel[3][4] ~^ image[14][13] + signed_kernel[4][0] ~^ image[15][9] + signed_kernel[4][1] ~^ image[15][10] + signed_kernel[4][2] ~^ image[15][11] + signed_kernel[4][3] ~^ image[15][12] + signed_kernel[4][4] ~^ image[15][13];
assign xor_sum[11][10] = signed_kernel[0][0] ~^ image[11][10] + signed_kernel[0][1] ~^ image[11][11] + signed_kernel[0][2] ~^ image[11][12] + signed_kernel[0][3] ~^ image[11][13] + signed_kernel[0][4] ~^ image[11][14] + signed_kernel[1][0] ~^ image[12][10] + signed_kernel[1][1] ~^ image[12][11] + signed_kernel[1][2] ~^ image[12][12] + signed_kernel[1][3] ~^ image[12][13] + signed_kernel[1][4] ~^ image[12][14] + signed_kernel[2][0] ~^ image[13][10] + signed_kernel[2][1] ~^ image[13][11] + signed_kernel[2][2] ~^ image[13][12] + signed_kernel[2][3] ~^ image[13][13] + signed_kernel[2][4] ~^ image[13][14] + signed_kernel[3][0] ~^ image[14][10] + signed_kernel[3][1] ~^ image[14][11] + signed_kernel[3][2] ~^ image[14][12] + signed_kernel[3][3] ~^ image[14][13] + signed_kernel[3][4] ~^ image[14][14] + signed_kernel[4][0] ~^ image[15][10] + signed_kernel[4][1] ~^ image[15][11] + signed_kernel[4][2] ~^ image[15][12] + signed_kernel[4][3] ~^ image[15][13] + signed_kernel[4][4] ~^ image[15][14];
assign xor_sum[11][11] = signed_kernel[0][0] ~^ image[11][11] + signed_kernel[0][1] ~^ image[11][12] + signed_kernel[0][2] ~^ image[11][13] + signed_kernel[0][3] ~^ image[11][14] + signed_kernel[0][4] ~^ image[11][15] + signed_kernel[1][0] ~^ image[12][11] + signed_kernel[1][1] ~^ image[12][12] + signed_kernel[1][2] ~^ image[12][13] + signed_kernel[1][3] ~^ image[12][14] + signed_kernel[1][4] ~^ image[12][15] + signed_kernel[2][0] ~^ image[13][11] + signed_kernel[2][1] ~^ image[13][12] + signed_kernel[2][2] ~^ image[13][13] + signed_kernel[2][3] ~^ image[13][14] + signed_kernel[2][4] ~^ image[13][15] + signed_kernel[3][0] ~^ image[14][11] + signed_kernel[3][1] ~^ image[14][12] + signed_kernel[3][2] ~^ image[14][13] + signed_kernel[3][3] ~^ image[14][14] + signed_kernel[3][4] ~^ image[14][15] + signed_kernel[4][0] ~^ image[15][11] + signed_kernel[4][1] ~^ image[15][12] + signed_kernel[4][2] ~^ image[15][13] + signed_kernel[4][3] ~^ image[15][14] + signed_kernel[4][4] ~^ image[15][15];
assign xor_sum[11][12] = signed_kernel[0][0] ~^ image[11][12] + signed_kernel[0][1] ~^ image[11][13] + signed_kernel[0][2] ~^ image[11][14] + signed_kernel[0][3] ~^ image[11][15] + signed_kernel[0][4] ~^ image[11][16] + signed_kernel[1][0] ~^ image[12][12] + signed_kernel[1][1] ~^ image[12][13] + signed_kernel[1][2] ~^ image[12][14] + signed_kernel[1][3] ~^ image[12][15] + signed_kernel[1][4] ~^ image[12][16] + signed_kernel[2][0] ~^ image[13][12] + signed_kernel[2][1] ~^ image[13][13] + signed_kernel[2][2] ~^ image[13][14] + signed_kernel[2][3] ~^ image[13][15] + signed_kernel[2][4] ~^ image[13][16] + signed_kernel[3][0] ~^ image[14][12] + signed_kernel[3][1] ~^ image[14][13] + signed_kernel[3][2] ~^ image[14][14] + signed_kernel[3][3] ~^ image[14][15] + signed_kernel[3][4] ~^ image[14][16] + signed_kernel[4][0] ~^ image[15][12] + signed_kernel[4][1] ~^ image[15][13] + signed_kernel[4][2] ~^ image[15][14] + signed_kernel[4][3] ~^ image[15][15] + signed_kernel[4][4] ~^ image[15][16];
assign xor_sum[11][13] = signed_kernel[0][0] ~^ image[11][13] + signed_kernel[0][1] ~^ image[11][14] + signed_kernel[0][2] ~^ image[11][15] + signed_kernel[0][3] ~^ image[11][16] + signed_kernel[0][4] ~^ image[11][17] + signed_kernel[1][0] ~^ image[12][13] + signed_kernel[1][1] ~^ image[12][14] + signed_kernel[1][2] ~^ image[12][15] + signed_kernel[1][3] ~^ image[12][16] + signed_kernel[1][4] ~^ image[12][17] + signed_kernel[2][0] ~^ image[13][13] + signed_kernel[2][1] ~^ image[13][14] + signed_kernel[2][2] ~^ image[13][15] + signed_kernel[2][3] ~^ image[13][16] + signed_kernel[2][4] ~^ image[13][17] + signed_kernel[3][0] ~^ image[14][13] + signed_kernel[3][1] ~^ image[14][14] + signed_kernel[3][2] ~^ image[14][15] + signed_kernel[3][3] ~^ image[14][16] + signed_kernel[3][4] ~^ image[14][17] + signed_kernel[4][0] ~^ image[15][13] + signed_kernel[4][1] ~^ image[15][14] + signed_kernel[4][2] ~^ image[15][15] + signed_kernel[4][3] ~^ image[15][16] + signed_kernel[4][4] ~^ image[15][17];
assign xor_sum[11][14] = signed_kernel[0][0] ~^ image[11][14] + signed_kernel[0][1] ~^ image[11][15] + signed_kernel[0][2] ~^ image[11][16] + signed_kernel[0][3] ~^ image[11][17] + signed_kernel[0][4] ~^ image[11][18] + signed_kernel[1][0] ~^ image[12][14] + signed_kernel[1][1] ~^ image[12][15] + signed_kernel[1][2] ~^ image[12][16] + signed_kernel[1][3] ~^ image[12][17] + signed_kernel[1][4] ~^ image[12][18] + signed_kernel[2][0] ~^ image[13][14] + signed_kernel[2][1] ~^ image[13][15] + signed_kernel[2][2] ~^ image[13][16] + signed_kernel[2][3] ~^ image[13][17] + signed_kernel[2][4] ~^ image[13][18] + signed_kernel[3][0] ~^ image[14][14] + signed_kernel[3][1] ~^ image[14][15] + signed_kernel[3][2] ~^ image[14][16] + signed_kernel[3][3] ~^ image[14][17] + signed_kernel[3][4] ~^ image[14][18] + signed_kernel[4][0] ~^ image[15][14] + signed_kernel[4][1] ~^ image[15][15] + signed_kernel[4][2] ~^ image[15][16] + signed_kernel[4][3] ~^ image[15][17] + signed_kernel[4][4] ~^ image[15][18];
assign xor_sum[11][15] = signed_kernel[0][0] ~^ image[11][15] + signed_kernel[0][1] ~^ image[11][16] + signed_kernel[0][2] ~^ image[11][17] + signed_kernel[0][3] ~^ image[11][18] + signed_kernel[0][4] ~^ image[11][19] + signed_kernel[1][0] ~^ image[12][15] + signed_kernel[1][1] ~^ image[12][16] + signed_kernel[1][2] ~^ image[12][17] + signed_kernel[1][3] ~^ image[12][18] + signed_kernel[1][4] ~^ image[12][19] + signed_kernel[2][0] ~^ image[13][15] + signed_kernel[2][1] ~^ image[13][16] + signed_kernel[2][2] ~^ image[13][17] + signed_kernel[2][3] ~^ image[13][18] + signed_kernel[2][4] ~^ image[13][19] + signed_kernel[3][0] ~^ image[14][15] + signed_kernel[3][1] ~^ image[14][16] + signed_kernel[3][2] ~^ image[14][17] + signed_kernel[3][3] ~^ image[14][18] + signed_kernel[3][4] ~^ image[14][19] + signed_kernel[4][0] ~^ image[15][15] + signed_kernel[4][1] ~^ image[15][16] + signed_kernel[4][2] ~^ image[15][17] + signed_kernel[4][3] ~^ image[15][18] + signed_kernel[4][4] ~^ image[15][19];
assign xor_sum[11][16] = signed_kernel[0][0] ~^ image[11][16] + signed_kernel[0][1] ~^ image[11][17] + signed_kernel[0][2] ~^ image[11][18] + signed_kernel[0][3] ~^ image[11][19] + signed_kernel[0][4] ~^ image[11][20] + signed_kernel[1][0] ~^ image[12][16] + signed_kernel[1][1] ~^ image[12][17] + signed_kernel[1][2] ~^ image[12][18] + signed_kernel[1][3] ~^ image[12][19] + signed_kernel[1][4] ~^ image[12][20] + signed_kernel[2][0] ~^ image[13][16] + signed_kernel[2][1] ~^ image[13][17] + signed_kernel[2][2] ~^ image[13][18] + signed_kernel[2][3] ~^ image[13][19] + signed_kernel[2][4] ~^ image[13][20] + signed_kernel[3][0] ~^ image[14][16] + signed_kernel[3][1] ~^ image[14][17] + signed_kernel[3][2] ~^ image[14][18] + signed_kernel[3][3] ~^ image[14][19] + signed_kernel[3][4] ~^ image[14][20] + signed_kernel[4][0] ~^ image[15][16] + signed_kernel[4][1] ~^ image[15][17] + signed_kernel[4][2] ~^ image[15][18] + signed_kernel[4][3] ~^ image[15][19] + signed_kernel[4][4] ~^ image[15][20];
assign xor_sum[11][17] = signed_kernel[0][0] ~^ image[11][17] + signed_kernel[0][1] ~^ image[11][18] + signed_kernel[0][2] ~^ image[11][19] + signed_kernel[0][3] ~^ image[11][20] + signed_kernel[0][4] ~^ image[11][21] + signed_kernel[1][0] ~^ image[12][17] + signed_kernel[1][1] ~^ image[12][18] + signed_kernel[1][2] ~^ image[12][19] + signed_kernel[1][3] ~^ image[12][20] + signed_kernel[1][4] ~^ image[12][21] + signed_kernel[2][0] ~^ image[13][17] + signed_kernel[2][1] ~^ image[13][18] + signed_kernel[2][2] ~^ image[13][19] + signed_kernel[2][3] ~^ image[13][20] + signed_kernel[2][4] ~^ image[13][21] + signed_kernel[3][0] ~^ image[14][17] + signed_kernel[3][1] ~^ image[14][18] + signed_kernel[3][2] ~^ image[14][19] + signed_kernel[3][3] ~^ image[14][20] + signed_kernel[3][4] ~^ image[14][21] + signed_kernel[4][0] ~^ image[15][17] + signed_kernel[4][1] ~^ image[15][18] + signed_kernel[4][2] ~^ image[15][19] + signed_kernel[4][3] ~^ image[15][20] + signed_kernel[4][4] ~^ image[15][21];
assign xor_sum[11][18] = signed_kernel[0][0] ~^ image[11][18] + signed_kernel[0][1] ~^ image[11][19] + signed_kernel[0][2] ~^ image[11][20] + signed_kernel[0][3] ~^ image[11][21] + signed_kernel[0][4] ~^ image[11][22] + signed_kernel[1][0] ~^ image[12][18] + signed_kernel[1][1] ~^ image[12][19] + signed_kernel[1][2] ~^ image[12][20] + signed_kernel[1][3] ~^ image[12][21] + signed_kernel[1][4] ~^ image[12][22] + signed_kernel[2][0] ~^ image[13][18] + signed_kernel[2][1] ~^ image[13][19] + signed_kernel[2][2] ~^ image[13][20] + signed_kernel[2][3] ~^ image[13][21] + signed_kernel[2][4] ~^ image[13][22] + signed_kernel[3][0] ~^ image[14][18] + signed_kernel[3][1] ~^ image[14][19] + signed_kernel[3][2] ~^ image[14][20] + signed_kernel[3][3] ~^ image[14][21] + signed_kernel[3][4] ~^ image[14][22] + signed_kernel[4][0] ~^ image[15][18] + signed_kernel[4][1] ~^ image[15][19] + signed_kernel[4][2] ~^ image[15][20] + signed_kernel[4][3] ~^ image[15][21] + signed_kernel[4][4] ~^ image[15][22];
assign xor_sum[11][19] = signed_kernel[0][0] ~^ image[11][19] + signed_kernel[0][1] ~^ image[11][20] + signed_kernel[0][2] ~^ image[11][21] + signed_kernel[0][3] ~^ image[11][22] + signed_kernel[0][4] ~^ image[11][23] + signed_kernel[1][0] ~^ image[12][19] + signed_kernel[1][1] ~^ image[12][20] + signed_kernel[1][2] ~^ image[12][21] + signed_kernel[1][3] ~^ image[12][22] + signed_kernel[1][4] ~^ image[12][23] + signed_kernel[2][0] ~^ image[13][19] + signed_kernel[2][1] ~^ image[13][20] + signed_kernel[2][2] ~^ image[13][21] + signed_kernel[2][3] ~^ image[13][22] + signed_kernel[2][4] ~^ image[13][23] + signed_kernel[3][0] ~^ image[14][19] + signed_kernel[3][1] ~^ image[14][20] + signed_kernel[3][2] ~^ image[14][21] + signed_kernel[3][3] ~^ image[14][22] + signed_kernel[3][4] ~^ image[14][23] + signed_kernel[4][0] ~^ image[15][19] + signed_kernel[4][1] ~^ image[15][20] + signed_kernel[4][2] ~^ image[15][21] + signed_kernel[4][3] ~^ image[15][22] + signed_kernel[4][4] ~^ image[15][23];
assign xor_sum[11][20] = signed_kernel[0][0] ~^ image[11][20] + signed_kernel[0][1] ~^ image[11][21] + signed_kernel[0][2] ~^ image[11][22] + signed_kernel[0][3] ~^ image[11][23] + signed_kernel[0][4] ~^ image[11][24] + signed_kernel[1][0] ~^ image[12][20] + signed_kernel[1][1] ~^ image[12][21] + signed_kernel[1][2] ~^ image[12][22] + signed_kernel[1][3] ~^ image[12][23] + signed_kernel[1][4] ~^ image[12][24] + signed_kernel[2][0] ~^ image[13][20] + signed_kernel[2][1] ~^ image[13][21] + signed_kernel[2][2] ~^ image[13][22] + signed_kernel[2][3] ~^ image[13][23] + signed_kernel[2][4] ~^ image[13][24] + signed_kernel[3][0] ~^ image[14][20] + signed_kernel[3][1] ~^ image[14][21] + signed_kernel[3][2] ~^ image[14][22] + signed_kernel[3][3] ~^ image[14][23] + signed_kernel[3][4] ~^ image[14][24] + signed_kernel[4][0] ~^ image[15][20] + signed_kernel[4][1] ~^ image[15][21] + signed_kernel[4][2] ~^ image[15][22] + signed_kernel[4][3] ~^ image[15][23] + signed_kernel[4][4] ~^ image[15][24];
assign xor_sum[11][21] = signed_kernel[0][0] ~^ image[11][21] + signed_kernel[0][1] ~^ image[11][22] + signed_kernel[0][2] ~^ image[11][23] + signed_kernel[0][3] ~^ image[11][24] + signed_kernel[0][4] ~^ image[11][25] + signed_kernel[1][0] ~^ image[12][21] + signed_kernel[1][1] ~^ image[12][22] + signed_kernel[1][2] ~^ image[12][23] + signed_kernel[1][3] ~^ image[12][24] + signed_kernel[1][4] ~^ image[12][25] + signed_kernel[2][0] ~^ image[13][21] + signed_kernel[2][1] ~^ image[13][22] + signed_kernel[2][2] ~^ image[13][23] + signed_kernel[2][3] ~^ image[13][24] + signed_kernel[2][4] ~^ image[13][25] + signed_kernel[3][0] ~^ image[14][21] + signed_kernel[3][1] ~^ image[14][22] + signed_kernel[3][2] ~^ image[14][23] + signed_kernel[3][3] ~^ image[14][24] + signed_kernel[3][4] ~^ image[14][25] + signed_kernel[4][0] ~^ image[15][21] + signed_kernel[4][1] ~^ image[15][22] + signed_kernel[4][2] ~^ image[15][23] + signed_kernel[4][3] ~^ image[15][24] + signed_kernel[4][4] ~^ image[15][25];
assign xor_sum[11][22] = signed_kernel[0][0] ~^ image[11][22] + signed_kernel[0][1] ~^ image[11][23] + signed_kernel[0][2] ~^ image[11][24] + signed_kernel[0][3] ~^ image[11][25] + signed_kernel[0][4] ~^ image[11][26] + signed_kernel[1][0] ~^ image[12][22] + signed_kernel[1][1] ~^ image[12][23] + signed_kernel[1][2] ~^ image[12][24] + signed_kernel[1][3] ~^ image[12][25] + signed_kernel[1][4] ~^ image[12][26] + signed_kernel[2][0] ~^ image[13][22] + signed_kernel[2][1] ~^ image[13][23] + signed_kernel[2][2] ~^ image[13][24] + signed_kernel[2][3] ~^ image[13][25] + signed_kernel[2][4] ~^ image[13][26] + signed_kernel[3][0] ~^ image[14][22] + signed_kernel[3][1] ~^ image[14][23] + signed_kernel[3][2] ~^ image[14][24] + signed_kernel[3][3] ~^ image[14][25] + signed_kernel[3][4] ~^ image[14][26] + signed_kernel[4][0] ~^ image[15][22] + signed_kernel[4][1] ~^ image[15][23] + signed_kernel[4][2] ~^ image[15][24] + signed_kernel[4][3] ~^ image[15][25] + signed_kernel[4][4] ~^ image[15][26];
assign xor_sum[11][23] = signed_kernel[0][0] ~^ image[11][23] + signed_kernel[0][1] ~^ image[11][24] + signed_kernel[0][2] ~^ image[11][25] + signed_kernel[0][3] ~^ image[11][26] + signed_kernel[0][4] ~^ image[11][27] + signed_kernel[1][0] ~^ image[12][23] + signed_kernel[1][1] ~^ image[12][24] + signed_kernel[1][2] ~^ image[12][25] + signed_kernel[1][3] ~^ image[12][26] + signed_kernel[1][4] ~^ image[12][27] + signed_kernel[2][0] ~^ image[13][23] + signed_kernel[2][1] ~^ image[13][24] + signed_kernel[2][2] ~^ image[13][25] + signed_kernel[2][3] ~^ image[13][26] + signed_kernel[2][4] ~^ image[13][27] + signed_kernel[3][0] ~^ image[14][23] + signed_kernel[3][1] ~^ image[14][24] + signed_kernel[3][2] ~^ image[14][25] + signed_kernel[3][3] ~^ image[14][26] + signed_kernel[3][4] ~^ image[14][27] + signed_kernel[4][0] ~^ image[15][23] + signed_kernel[4][1] ~^ image[15][24] + signed_kernel[4][2] ~^ image[15][25] + signed_kernel[4][3] ~^ image[15][26] + signed_kernel[4][4] ~^ image[15][27];
assign xor_sum[12][0] = signed_kernel[0][0] ~^ image[12][0] + signed_kernel[0][1] ~^ image[12][1] + signed_kernel[0][2] ~^ image[12][2] + signed_kernel[0][3] ~^ image[12][3] + signed_kernel[0][4] ~^ image[12][4] + signed_kernel[1][0] ~^ image[13][0] + signed_kernel[1][1] ~^ image[13][1] + signed_kernel[1][2] ~^ image[13][2] + signed_kernel[1][3] ~^ image[13][3] + signed_kernel[1][4] ~^ image[13][4] + signed_kernel[2][0] ~^ image[14][0] + signed_kernel[2][1] ~^ image[14][1] + signed_kernel[2][2] ~^ image[14][2] + signed_kernel[2][3] ~^ image[14][3] + signed_kernel[2][4] ~^ image[14][4] + signed_kernel[3][0] ~^ image[15][0] + signed_kernel[3][1] ~^ image[15][1] + signed_kernel[3][2] ~^ image[15][2] + signed_kernel[3][3] ~^ image[15][3] + signed_kernel[3][4] ~^ image[15][4] + signed_kernel[4][0] ~^ image[16][0] + signed_kernel[4][1] ~^ image[16][1] + signed_kernel[4][2] ~^ image[16][2] + signed_kernel[4][3] ~^ image[16][3] + signed_kernel[4][4] ~^ image[16][4];
assign xor_sum[12][1] = signed_kernel[0][0] ~^ image[12][1] + signed_kernel[0][1] ~^ image[12][2] + signed_kernel[0][2] ~^ image[12][3] + signed_kernel[0][3] ~^ image[12][4] + signed_kernel[0][4] ~^ image[12][5] + signed_kernel[1][0] ~^ image[13][1] + signed_kernel[1][1] ~^ image[13][2] + signed_kernel[1][2] ~^ image[13][3] + signed_kernel[1][3] ~^ image[13][4] + signed_kernel[1][4] ~^ image[13][5] + signed_kernel[2][0] ~^ image[14][1] + signed_kernel[2][1] ~^ image[14][2] + signed_kernel[2][2] ~^ image[14][3] + signed_kernel[2][3] ~^ image[14][4] + signed_kernel[2][4] ~^ image[14][5] + signed_kernel[3][0] ~^ image[15][1] + signed_kernel[3][1] ~^ image[15][2] + signed_kernel[3][2] ~^ image[15][3] + signed_kernel[3][3] ~^ image[15][4] + signed_kernel[3][4] ~^ image[15][5] + signed_kernel[4][0] ~^ image[16][1] + signed_kernel[4][1] ~^ image[16][2] + signed_kernel[4][2] ~^ image[16][3] + signed_kernel[4][3] ~^ image[16][4] + signed_kernel[4][4] ~^ image[16][5];
assign xor_sum[12][2] = signed_kernel[0][0] ~^ image[12][2] + signed_kernel[0][1] ~^ image[12][3] + signed_kernel[0][2] ~^ image[12][4] + signed_kernel[0][3] ~^ image[12][5] + signed_kernel[0][4] ~^ image[12][6] + signed_kernel[1][0] ~^ image[13][2] + signed_kernel[1][1] ~^ image[13][3] + signed_kernel[1][2] ~^ image[13][4] + signed_kernel[1][3] ~^ image[13][5] + signed_kernel[1][4] ~^ image[13][6] + signed_kernel[2][0] ~^ image[14][2] + signed_kernel[2][1] ~^ image[14][3] + signed_kernel[2][2] ~^ image[14][4] + signed_kernel[2][3] ~^ image[14][5] + signed_kernel[2][4] ~^ image[14][6] + signed_kernel[3][0] ~^ image[15][2] + signed_kernel[3][1] ~^ image[15][3] + signed_kernel[3][2] ~^ image[15][4] + signed_kernel[3][3] ~^ image[15][5] + signed_kernel[3][4] ~^ image[15][6] + signed_kernel[4][0] ~^ image[16][2] + signed_kernel[4][1] ~^ image[16][3] + signed_kernel[4][2] ~^ image[16][4] + signed_kernel[4][3] ~^ image[16][5] + signed_kernel[4][4] ~^ image[16][6];
assign xor_sum[12][3] = signed_kernel[0][0] ~^ image[12][3] + signed_kernel[0][1] ~^ image[12][4] + signed_kernel[0][2] ~^ image[12][5] + signed_kernel[0][3] ~^ image[12][6] + signed_kernel[0][4] ~^ image[12][7] + signed_kernel[1][0] ~^ image[13][3] + signed_kernel[1][1] ~^ image[13][4] + signed_kernel[1][2] ~^ image[13][5] + signed_kernel[1][3] ~^ image[13][6] + signed_kernel[1][4] ~^ image[13][7] + signed_kernel[2][0] ~^ image[14][3] + signed_kernel[2][1] ~^ image[14][4] + signed_kernel[2][2] ~^ image[14][5] + signed_kernel[2][3] ~^ image[14][6] + signed_kernel[2][4] ~^ image[14][7] + signed_kernel[3][0] ~^ image[15][3] + signed_kernel[3][1] ~^ image[15][4] + signed_kernel[3][2] ~^ image[15][5] + signed_kernel[3][3] ~^ image[15][6] + signed_kernel[3][4] ~^ image[15][7] + signed_kernel[4][0] ~^ image[16][3] + signed_kernel[4][1] ~^ image[16][4] + signed_kernel[4][2] ~^ image[16][5] + signed_kernel[4][3] ~^ image[16][6] + signed_kernel[4][4] ~^ image[16][7];
assign xor_sum[12][4] = signed_kernel[0][0] ~^ image[12][4] + signed_kernel[0][1] ~^ image[12][5] + signed_kernel[0][2] ~^ image[12][6] + signed_kernel[0][3] ~^ image[12][7] + signed_kernel[0][4] ~^ image[12][8] + signed_kernel[1][0] ~^ image[13][4] + signed_kernel[1][1] ~^ image[13][5] + signed_kernel[1][2] ~^ image[13][6] + signed_kernel[1][3] ~^ image[13][7] + signed_kernel[1][4] ~^ image[13][8] + signed_kernel[2][0] ~^ image[14][4] + signed_kernel[2][1] ~^ image[14][5] + signed_kernel[2][2] ~^ image[14][6] + signed_kernel[2][3] ~^ image[14][7] + signed_kernel[2][4] ~^ image[14][8] + signed_kernel[3][0] ~^ image[15][4] + signed_kernel[3][1] ~^ image[15][5] + signed_kernel[3][2] ~^ image[15][6] + signed_kernel[3][3] ~^ image[15][7] + signed_kernel[3][4] ~^ image[15][8] + signed_kernel[4][0] ~^ image[16][4] + signed_kernel[4][1] ~^ image[16][5] + signed_kernel[4][2] ~^ image[16][6] + signed_kernel[4][3] ~^ image[16][7] + signed_kernel[4][4] ~^ image[16][8];
assign xor_sum[12][5] = signed_kernel[0][0] ~^ image[12][5] + signed_kernel[0][1] ~^ image[12][6] + signed_kernel[0][2] ~^ image[12][7] + signed_kernel[0][3] ~^ image[12][8] + signed_kernel[0][4] ~^ image[12][9] + signed_kernel[1][0] ~^ image[13][5] + signed_kernel[1][1] ~^ image[13][6] + signed_kernel[1][2] ~^ image[13][7] + signed_kernel[1][3] ~^ image[13][8] + signed_kernel[1][4] ~^ image[13][9] + signed_kernel[2][0] ~^ image[14][5] + signed_kernel[2][1] ~^ image[14][6] + signed_kernel[2][2] ~^ image[14][7] + signed_kernel[2][3] ~^ image[14][8] + signed_kernel[2][4] ~^ image[14][9] + signed_kernel[3][0] ~^ image[15][5] + signed_kernel[3][1] ~^ image[15][6] + signed_kernel[3][2] ~^ image[15][7] + signed_kernel[3][3] ~^ image[15][8] + signed_kernel[3][4] ~^ image[15][9] + signed_kernel[4][0] ~^ image[16][5] + signed_kernel[4][1] ~^ image[16][6] + signed_kernel[4][2] ~^ image[16][7] + signed_kernel[4][3] ~^ image[16][8] + signed_kernel[4][4] ~^ image[16][9];
assign xor_sum[12][6] = signed_kernel[0][0] ~^ image[12][6] + signed_kernel[0][1] ~^ image[12][7] + signed_kernel[0][2] ~^ image[12][8] + signed_kernel[0][3] ~^ image[12][9] + signed_kernel[0][4] ~^ image[12][10] + signed_kernel[1][0] ~^ image[13][6] + signed_kernel[1][1] ~^ image[13][7] + signed_kernel[1][2] ~^ image[13][8] + signed_kernel[1][3] ~^ image[13][9] + signed_kernel[1][4] ~^ image[13][10] + signed_kernel[2][0] ~^ image[14][6] + signed_kernel[2][1] ~^ image[14][7] + signed_kernel[2][2] ~^ image[14][8] + signed_kernel[2][3] ~^ image[14][9] + signed_kernel[2][4] ~^ image[14][10] + signed_kernel[3][0] ~^ image[15][6] + signed_kernel[3][1] ~^ image[15][7] + signed_kernel[3][2] ~^ image[15][8] + signed_kernel[3][3] ~^ image[15][9] + signed_kernel[3][4] ~^ image[15][10] + signed_kernel[4][0] ~^ image[16][6] + signed_kernel[4][1] ~^ image[16][7] + signed_kernel[4][2] ~^ image[16][8] + signed_kernel[4][3] ~^ image[16][9] + signed_kernel[4][4] ~^ image[16][10];
assign xor_sum[12][7] = signed_kernel[0][0] ~^ image[12][7] + signed_kernel[0][1] ~^ image[12][8] + signed_kernel[0][2] ~^ image[12][9] + signed_kernel[0][3] ~^ image[12][10] + signed_kernel[0][4] ~^ image[12][11] + signed_kernel[1][0] ~^ image[13][7] + signed_kernel[1][1] ~^ image[13][8] + signed_kernel[1][2] ~^ image[13][9] + signed_kernel[1][3] ~^ image[13][10] + signed_kernel[1][4] ~^ image[13][11] + signed_kernel[2][0] ~^ image[14][7] + signed_kernel[2][1] ~^ image[14][8] + signed_kernel[2][2] ~^ image[14][9] + signed_kernel[2][3] ~^ image[14][10] + signed_kernel[2][4] ~^ image[14][11] + signed_kernel[3][0] ~^ image[15][7] + signed_kernel[3][1] ~^ image[15][8] + signed_kernel[3][2] ~^ image[15][9] + signed_kernel[3][3] ~^ image[15][10] + signed_kernel[3][4] ~^ image[15][11] + signed_kernel[4][0] ~^ image[16][7] + signed_kernel[4][1] ~^ image[16][8] + signed_kernel[4][2] ~^ image[16][9] + signed_kernel[4][3] ~^ image[16][10] + signed_kernel[4][4] ~^ image[16][11];
assign xor_sum[12][8] = signed_kernel[0][0] ~^ image[12][8] + signed_kernel[0][1] ~^ image[12][9] + signed_kernel[0][2] ~^ image[12][10] + signed_kernel[0][3] ~^ image[12][11] + signed_kernel[0][4] ~^ image[12][12] + signed_kernel[1][0] ~^ image[13][8] + signed_kernel[1][1] ~^ image[13][9] + signed_kernel[1][2] ~^ image[13][10] + signed_kernel[1][3] ~^ image[13][11] + signed_kernel[1][4] ~^ image[13][12] + signed_kernel[2][0] ~^ image[14][8] + signed_kernel[2][1] ~^ image[14][9] + signed_kernel[2][2] ~^ image[14][10] + signed_kernel[2][3] ~^ image[14][11] + signed_kernel[2][4] ~^ image[14][12] + signed_kernel[3][0] ~^ image[15][8] + signed_kernel[3][1] ~^ image[15][9] + signed_kernel[3][2] ~^ image[15][10] + signed_kernel[3][3] ~^ image[15][11] + signed_kernel[3][4] ~^ image[15][12] + signed_kernel[4][0] ~^ image[16][8] + signed_kernel[4][1] ~^ image[16][9] + signed_kernel[4][2] ~^ image[16][10] + signed_kernel[4][3] ~^ image[16][11] + signed_kernel[4][4] ~^ image[16][12];
assign xor_sum[12][9] = signed_kernel[0][0] ~^ image[12][9] + signed_kernel[0][1] ~^ image[12][10] + signed_kernel[0][2] ~^ image[12][11] + signed_kernel[0][3] ~^ image[12][12] + signed_kernel[0][4] ~^ image[12][13] + signed_kernel[1][0] ~^ image[13][9] + signed_kernel[1][1] ~^ image[13][10] + signed_kernel[1][2] ~^ image[13][11] + signed_kernel[1][3] ~^ image[13][12] + signed_kernel[1][4] ~^ image[13][13] + signed_kernel[2][0] ~^ image[14][9] + signed_kernel[2][1] ~^ image[14][10] + signed_kernel[2][2] ~^ image[14][11] + signed_kernel[2][3] ~^ image[14][12] + signed_kernel[2][4] ~^ image[14][13] + signed_kernel[3][0] ~^ image[15][9] + signed_kernel[3][1] ~^ image[15][10] + signed_kernel[3][2] ~^ image[15][11] + signed_kernel[3][3] ~^ image[15][12] + signed_kernel[3][4] ~^ image[15][13] + signed_kernel[4][0] ~^ image[16][9] + signed_kernel[4][1] ~^ image[16][10] + signed_kernel[4][2] ~^ image[16][11] + signed_kernel[4][3] ~^ image[16][12] + signed_kernel[4][4] ~^ image[16][13];
assign xor_sum[12][10] = signed_kernel[0][0] ~^ image[12][10] + signed_kernel[0][1] ~^ image[12][11] + signed_kernel[0][2] ~^ image[12][12] + signed_kernel[0][3] ~^ image[12][13] + signed_kernel[0][4] ~^ image[12][14] + signed_kernel[1][0] ~^ image[13][10] + signed_kernel[1][1] ~^ image[13][11] + signed_kernel[1][2] ~^ image[13][12] + signed_kernel[1][3] ~^ image[13][13] + signed_kernel[1][4] ~^ image[13][14] + signed_kernel[2][0] ~^ image[14][10] + signed_kernel[2][1] ~^ image[14][11] + signed_kernel[2][2] ~^ image[14][12] + signed_kernel[2][3] ~^ image[14][13] + signed_kernel[2][4] ~^ image[14][14] + signed_kernel[3][0] ~^ image[15][10] + signed_kernel[3][1] ~^ image[15][11] + signed_kernel[3][2] ~^ image[15][12] + signed_kernel[3][3] ~^ image[15][13] + signed_kernel[3][4] ~^ image[15][14] + signed_kernel[4][0] ~^ image[16][10] + signed_kernel[4][1] ~^ image[16][11] + signed_kernel[4][2] ~^ image[16][12] + signed_kernel[4][3] ~^ image[16][13] + signed_kernel[4][4] ~^ image[16][14];
assign xor_sum[12][11] = signed_kernel[0][0] ~^ image[12][11] + signed_kernel[0][1] ~^ image[12][12] + signed_kernel[0][2] ~^ image[12][13] + signed_kernel[0][3] ~^ image[12][14] + signed_kernel[0][4] ~^ image[12][15] + signed_kernel[1][0] ~^ image[13][11] + signed_kernel[1][1] ~^ image[13][12] + signed_kernel[1][2] ~^ image[13][13] + signed_kernel[1][3] ~^ image[13][14] + signed_kernel[1][4] ~^ image[13][15] + signed_kernel[2][0] ~^ image[14][11] + signed_kernel[2][1] ~^ image[14][12] + signed_kernel[2][2] ~^ image[14][13] + signed_kernel[2][3] ~^ image[14][14] + signed_kernel[2][4] ~^ image[14][15] + signed_kernel[3][0] ~^ image[15][11] + signed_kernel[3][1] ~^ image[15][12] + signed_kernel[3][2] ~^ image[15][13] + signed_kernel[3][3] ~^ image[15][14] + signed_kernel[3][4] ~^ image[15][15] + signed_kernel[4][0] ~^ image[16][11] + signed_kernel[4][1] ~^ image[16][12] + signed_kernel[4][2] ~^ image[16][13] + signed_kernel[4][3] ~^ image[16][14] + signed_kernel[4][4] ~^ image[16][15];
assign xor_sum[12][12] = signed_kernel[0][0] ~^ image[12][12] + signed_kernel[0][1] ~^ image[12][13] + signed_kernel[0][2] ~^ image[12][14] + signed_kernel[0][3] ~^ image[12][15] + signed_kernel[0][4] ~^ image[12][16] + signed_kernel[1][0] ~^ image[13][12] + signed_kernel[1][1] ~^ image[13][13] + signed_kernel[1][2] ~^ image[13][14] + signed_kernel[1][3] ~^ image[13][15] + signed_kernel[1][4] ~^ image[13][16] + signed_kernel[2][0] ~^ image[14][12] + signed_kernel[2][1] ~^ image[14][13] + signed_kernel[2][2] ~^ image[14][14] + signed_kernel[2][3] ~^ image[14][15] + signed_kernel[2][4] ~^ image[14][16] + signed_kernel[3][0] ~^ image[15][12] + signed_kernel[3][1] ~^ image[15][13] + signed_kernel[3][2] ~^ image[15][14] + signed_kernel[3][3] ~^ image[15][15] + signed_kernel[3][4] ~^ image[15][16] + signed_kernel[4][0] ~^ image[16][12] + signed_kernel[4][1] ~^ image[16][13] + signed_kernel[4][2] ~^ image[16][14] + signed_kernel[4][3] ~^ image[16][15] + signed_kernel[4][4] ~^ image[16][16];
assign xor_sum[12][13] = signed_kernel[0][0] ~^ image[12][13] + signed_kernel[0][1] ~^ image[12][14] + signed_kernel[0][2] ~^ image[12][15] + signed_kernel[0][3] ~^ image[12][16] + signed_kernel[0][4] ~^ image[12][17] + signed_kernel[1][0] ~^ image[13][13] + signed_kernel[1][1] ~^ image[13][14] + signed_kernel[1][2] ~^ image[13][15] + signed_kernel[1][3] ~^ image[13][16] + signed_kernel[1][4] ~^ image[13][17] + signed_kernel[2][0] ~^ image[14][13] + signed_kernel[2][1] ~^ image[14][14] + signed_kernel[2][2] ~^ image[14][15] + signed_kernel[2][3] ~^ image[14][16] + signed_kernel[2][4] ~^ image[14][17] + signed_kernel[3][0] ~^ image[15][13] + signed_kernel[3][1] ~^ image[15][14] + signed_kernel[3][2] ~^ image[15][15] + signed_kernel[3][3] ~^ image[15][16] + signed_kernel[3][4] ~^ image[15][17] + signed_kernel[4][0] ~^ image[16][13] + signed_kernel[4][1] ~^ image[16][14] + signed_kernel[4][2] ~^ image[16][15] + signed_kernel[4][3] ~^ image[16][16] + signed_kernel[4][4] ~^ image[16][17];
assign xor_sum[12][14] = signed_kernel[0][0] ~^ image[12][14] + signed_kernel[0][1] ~^ image[12][15] + signed_kernel[0][2] ~^ image[12][16] + signed_kernel[0][3] ~^ image[12][17] + signed_kernel[0][4] ~^ image[12][18] + signed_kernel[1][0] ~^ image[13][14] + signed_kernel[1][1] ~^ image[13][15] + signed_kernel[1][2] ~^ image[13][16] + signed_kernel[1][3] ~^ image[13][17] + signed_kernel[1][4] ~^ image[13][18] + signed_kernel[2][0] ~^ image[14][14] + signed_kernel[2][1] ~^ image[14][15] + signed_kernel[2][2] ~^ image[14][16] + signed_kernel[2][3] ~^ image[14][17] + signed_kernel[2][4] ~^ image[14][18] + signed_kernel[3][0] ~^ image[15][14] + signed_kernel[3][1] ~^ image[15][15] + signed_kernel[3][2] ~^ image[15][16] + signed_kernel[3][3] ~^ image[15][17] + signed_kernel[3][4] ~^ image[15][18] + signed_kernel[4][0] ~^ image[16][14] + signed_kernel[4][1] ~^ image[16][15] + signed_kernel[4][2] ~^ image[16][16] + signed_kernel[4][3] ~^ image[16][17] + signed_kernel[4][4] ~^ image[16][18];
assign xor_sum[12][15] = signed_kernel[0][0] ~^ image[12][15] + signed_kernel[0][1] ~^ image[12][16] + signed_kernel[0][2] ~^ image[12][17] + signed_kernel[0][3] ~^ image[12][18] + signed_kernel[0][4] ~^ image[12][19] + signed_kernel[1][0] ~^ image[13][15] + signed_kernel[1][1] ~^ image[13][16] + signed_kernel[1][2] ~^ image[13][17] + signed_kernel[1][3] ~^ image[13][18] + signed_kernel[1][4] ~^ image[13][19] + signed_kernel[2][0] ~^ image[14][15] + signed_kernel[2][1] ~^ image[14][16] + signed_kernel[2][2] ~^ image[14][17] + signed_kernel[2][3] ~^ image[14][18] + signed_kernel[2][4] ~^ image[14][19] + signed_kernel[3][0] ~^ image[15][15] + signed_kernel[3][1] ~^ image[15][16] + signed_kernel[3][2] ~^ image[15][17] + signed_kernel[3][3] ~^ image[15][18] + signed_kernel[3][4] ~^ image[15][19] + signed_kernel[4][0] ~^ image[16][15] + signed_kernel[4][1] ~^ image[16][16] + signed_kernel[4][2] ~^ image[16][17] + signed_kernel[4][3] ~^ image[16][18] + signed_kernel[4][4] ~^ image[16][19];
assign xor_sum[12][16] = signed_kernel[0][0] ~^ image[12][16] + signed_kernel[0][1] ~^ image[12][17] + signed_kernel[0][2] ~^ image[12][18] + signed_kernel[0][3] ~^ image[12][19] + signed_kernel[0][4] ~^ image[12][20] + signed_kernel[1][0] ~^ image[13][16] + signed_kernel[1][1] ~^ image[13][17] + signed_kernel[1][2] ~^ image[13][18] + signed_kernel[1][3] ~^ image[13][19] + signed_kernel[1][4] ~^ image[13][20] + signed_kernel[2][0] ~^ image[14][16] + signed_kernel[2][1] ~^ image[14][17] + signed_kernel[2][2] ~^ image[14][18] + signed_kernel[2][3] ~^ image[14][19] + signed_kernel[2][4] ~^ image[14][20] + signed_kernel[3][0] ~^ image[15][16] + signed_kernel[3][1] ~^ image[15][17] + signed_kernel[3][2] ~^ image[15][18] + signed_kernel[3][3] ~^ image[15][19] + signed_kernel[3][4] ~^ image[15][20] + signed_kernel[4][0] ~^ image[16][16] + signed_kernel[4][1] ~^ image[16][17] + signed_kernel[4][2] ~^ image[16][18] + signed_kernel[4][3] ~^ image[16][19] + signed_kernel[4][4] ~^ image[16][20];
assign xor_sum[12][17] = signed_kernel[0][0] ~^ image[12][17] + signed_kernel[0][1] ~^ image[12][18] + signed_kernel[0][2] ~^ image[12][19] + signed_kernel[0][3] ~^ image[12][20] + signed_kernel[0][4] ~^ image[12][21] + signed_kernel[1][0] ~^ image[13][17] + signed_kernel[1][1] ~^ image[13][18] + signed_kernel[1][2] ~^ image[13][19] + signed_kernel[1][3] ~^ image[13][20] + signed_kernel[1][4] ~^ image[13][21] + signed_kernel[2][0] ~^ image[14][17] + signed_kernel[2][1] ~^ image[14][18] + signed_kernel[2][2] ~^ image[14][19] + signed_kernel[2][3] ~^ image[14][20] + signed_kernel[2][4] ~^ image[14][21] + signed_kernel[3][0] ~^ image[15][17] + signed_kernel[3][1] ~^ image[15][18] + signed_kernel[3][2] ~^ image[15][19] + signed_kernel[3][3] ~^ image[15][20] + signed_kernel[3][4] ~^ image[15][21] + signed_kernel[4][0] ~^ image[16][17] + signed_kernel[4][1] ~^ image[16][18] + signed_kernel[4][2] ~^ image[16][19] + signed_kernel[4][3] ~^ image[16][20] + signed_kernel[4][4] ~^ image[16][21];
assign xor_sum[12][18] = signed_kernel[0][0] ~^ image[12][18] + signed_kernel[0][1] ~^ image[12][19] + signed_kernel[0][2] ~^ image[12][20] + signed_kernel[0][3] ~^ image[12][21] + signed_kernel[0][4] ~^ image[12][22] + signed_kernel[1][0] ~^ image[13][18] + signed_kernel[1][1] ~^ image[13][19] + signed_kernel[1][2] ~^ image[13][20] + signed_kernel[1][3] ~^ image[13][21] + signed_kernel[1][4] ~^ image[13][22] + signed_kernel[2][0] ~^ image[14][18] + signed_kernel[2][1] ~^ image[14][19] + signed_kernel[2][2] ~^ image[14][20] + signed_kernel[2][3] ~^ image[14][21] + signed_kernel[2][4] ~^ image[14][22] + signed_kernel[3][0] ~^ image[15][18] + signed_kernel[3][1] ~^ image[15][19] + signed_kernel[3][2] ~^ image[15][20] + signed_kernel[3][3] ~^ image[15][21] + signed_kernel[3][4] ~^ image[15][22] + signed_kernel[4][0] ~^ image[16][18] + signed_kernel[4][1] ~^ image[16][19] + signed_kernel[4][2] ~^ image[16][20] + signed_kernel[4][3] ~^ image[16][21] + signed_kernel[4][4] ~^ image[16][22];
assign xor_sum[12][19] = signed_kernel[0][0] ~^ image[12][19] + signed_kernel[0][1] ~^ image[12][20] + signed_kernel[0][2] ~^ image[12][21] + signed_kernel[0][3] ~^ image[12][22] + signed_kernel[0][4] ~^ image[12][23] + signed_kernel[1][0] ~^ image[13][19] + signed_kernel[1][1] ~^ image[13][20] + signed_kernel[1][2] ~^ image[13][21] + signed_kernel[1][3] ~^ image[13][22] + signed_kernel[1][4] ~^ image[13][23] + signed_kernel[2][0] ~^ image[14][19] + signed_kernel[2][1] ~^ image[14][20] + signed_kernel[2][2] ~^ image[14][21] + signed_kernel[2][3] ~^ image[14][22] + signed_kernel[2][4] ~^ image[14][23] + signed_kernel[3][0] ~^ image[15][19] + signed_kernel[3][1] ~^ image[15][20] + signed_kernel[3][2] ~^ image[15][21] + signed_kernel[3][3] ~^ image[15][22] + signed_kernel[3][4] ~^ image[15][23] + signed_kernel[4][0] ~^ image[16][19] + signed_kernel[4][1] ~^ image[16][20] + signed_kernel[4][2] ~^ image[16][21] + signed_kernel[4][3] ~^ image[16][22] + signed_kernel[4][4] ~^ image[16][23];
assign xor_sum[12][20] = signed_kernel[0][0] ~^ image[12][20] + signed_kernel[0][1] ~^ image[12][21] + signed_kernel[0][2] ~^ image[12][22] + signed_kernel[0][3] ~^ image[12][23] + signed_kernel[0][4] ~^ image[12][24] + signed_kernel[1][0] ~^ image[13][20] + signed_kernel[1][1] ~^ image[13][21] + signed_kernel[1][2] ~^ image[13][22] + signed_kernel[1][3] ~^ image[13][23] + signed_kernel[1][4] ~^ image[13][24] + signed_kernel[2][0] ~^ image[14][20] + signed_kernel[2][1] ~^ image[14][21] + signed_kernel[2][2] ~^ image[14][22] + signed_kernel[2][3] ~^ image[14][23] + signed_kernel[2][4] ~^ image[14][24] + signed_kernel[3][0] ~^ image[15][20] + signed_kernel[3][1] ~^ image[15][21] + signed_kernel[3][2] ~^ image[15][22] + signed_kernel[3][3] ~^ image[15][23] + signed_kernel[3][4] ~^ image[15][24] + signed_kernel[4][0] ~^ image[16][20] + signed_kernel[4][1] ~^ image[16][21] + signed_kernel[4][2] ~^ image[16][22] + signed_kernel[4][3] ~^ image[16][23] + signed_kernel[4][4] ~^ image[16][24];
assign xor_sum[12][21] = signed_kernel[0][0] ~^ image[12][21] + signed_kernel[0][1] ~^ image[12][22] + signed_kernel[0][2] ~^ image[12][23] + signed_kernel[0][3] ~^ image[12][24] + signed_kernel[0][4] ~^ image[12][25] + signed_kernel[1][0] ~^ image[13][21] + signed_kernel[1][1] ~^ image[13][22] + signed_kernel[1][2] ~^ image[13][23] + signed_kernel[1][3] ~^ image[13][24] + signed_kernel[1][4] ~^ image[13][25] + signed_kernel[2][0] ~^ image[14][21] + signed_kernel[2][1] ~^ image[14][22] + signed_kernel[2][2] ~^ image[14][23] + signed_kernel[2][3] ~^ image[14][24] + signed_kernel[2][4] ~^ image[14][25] + signed_kernel[3][0] ~^ image[15][21] + signed_kernel[3][1] ~^ image[15][22] + signed_kernel[3][2] ~^ image[15][23] + signed_kernel[3][3] ~^ image[15][24] + signed_kernel[3][4] ~^ image[15][25] + signed_kernel[4][0] ~^ image[16][21] + signed_kernel[4][1] ~^ image[16][22] + signed_kernel[4][2] ~^ image[16][23] + signed_kernel[4][3] ~^ image[16][24] + signed_kernel[4][4] ~^ image[16][25];
assign xor_sum[12][22] = signed_kernel[0][0] ~^ image[12][22] + signed_kernel[0][1] ~^ image[12][23] + signed_kernel[0][2] ~^ image[12][24] + signed_kernel[0][3] ~^ image[12][25] + signed_kernel[0][4] ~^ image[12][26] + signed_kernel[1][0] ~^ image[13][22] + signed_kernel[1][1] ~^ image[13][23] + signed_kernel[1][2] ~^ image[13][24] + signed_kernel[1][3] ~^ image[13][25] + signed_kernel[1][4] ~^ image[13][26] + signed_kernel[2][0] ~^ image[14][22] + signed_kernel[2][1] ~^ image[14][23] + signed_kernel[2][2] ~^ image[14][24] + signed_kernel[2][3] ~^ image[14][25] + signed_kernel[2][4] ~^ image[14][26] + signed_kernel[3][0] ~^ image[15][22] + signed_kernel[3][1] ~^ image[15][23] + signed_kernel[3][2] ~^ image[15][24] + signed_kernel[3][3] ~^ image[15][25] + signed_kernel[3][4] ~^ image[15][26] + signed_kernel[4][0] ~^ image[16][22] + signed_kernel[4][1] ~^ image[16][23] + signed_kernel[4][2] ~^ image[16][24] + signed_kernel[4][3] ~^ image[16][25] + signed_kernel[4][4] ~^ image[16][26];
assign xor_sum[12][23] = signed_kernel[0][0] ~^ image[12][23] + signed_kernel[0][1] ~^ image[12][24] + signed_kernel[0][2] ~^ image[12][25] + signed_kernel[0][3] ~^ image[12][26] + signed_kernel[0][4] ~^ image[12][27] + signed_kernel[1][0] ~^ image[13][23] + signed_kernel[1][1] ~^ image[13][24] + signed_kernel[1][2] ~^ image[13][25] + signed_kernel[1][3] ~^ image[13][26] + signed_kernel[1][4] ~^ image[13][27] + signed_kernel[2][0] ~^ image[14][23] + signed_kernel[2][1] ~^ image[14][24] + signed_kernel[2][2] ~^ image[14][25] + signed_kernel[2][3] ~^ image[14][26] + signed_kernel[2][4] ~^ image[14][27] + signed_kernel[3][0] ~^ image[15][23] + signed_kernel[3][1] ~^ image[15][24] + signed_kernel[3][2] ~^ image[15][25] + signed_kernel[3][3] ~^ image[15][26] + signed_kernel[3][4] ~^ image[15][27] + signed_kernel[4][0] ~^ image[16][23] + signed_kernel[4][1] ~^ image[16][24] + signed_kernel[4][2] ~^ image[16][25] + signed_kernel[4][3] ~^ image[16][26] + signed_kernel[4][4] ~^ image[16][27];
assign xor_sum[13][0] = signed_kernel[0][0] ~^ image[13][0] + signed_kernel[0][1] ~^ image[13][1] + signed_kernel[0][2] ~^ image[13][2] + signed_kernel[0][3] ~^ image[13][3] + signed_kernel[0][4] ~^ image[13][4] + signed_kernel[1][0] ~^ image[14][0] + signed_kernel[1][1] ~^ image[14][1] + signed_kernel[1][2] ~^ image[14][2] + signed_kernel[1][3] ~^ image[14][3] + signed_kernel[1][4] ~^ image[14][4] + signed_kernel[2][0] ~^ image[15][0] + signed_kernel[2][1] ~^ image[15][1] + signed_kernel[2][2] ~^ image[15][2] + signed_kernel[2][3] ~^ image[15][3] + signed_kernel[2][4] ~^ image[15][4] + signed_kernel[3][0] ~^ image[16][0] + signed_kernel[3][1] ~^ image[16][1] + signed_kernel[3][2] ~^ image[16][2] + signed_kernel[3][3] ~^ image[16][3] + signed_kernel[3][4] ~^ image[16][4] + signed_kernel[4][0] ~^ image[17][0] + signed_kernel[4][1] ~^ image[17][1] + signed_kernel[4][2] ~^ image[17][2] + signed_kernel[4][3] ~^ image[17][3] + signed_kernel[4][4] ~^ image[17][4];
assign xor_sum[13][1] = signed_kernel[0][0] ~^ image[13][1] + signed_kernel[0][1] ~^ image[13][2] + signed_kernel[0][2] ~^ image[13][3] + signed_kernel[0][3] ~^ image[13][4] + signed_kernel[0][4] ~^ image[13][5] + signed_kernel[1][0] ~^ image[14][1] + signed_kernel[1][1] ~^ image[14][2] + signed_kernel[1][2] ~^ image[14][3] + signed_kernel[1][3] ~^ image[14][4] + signed_kernel[1][4] ~^ image[14][5] + signed_kernel[2][0] ~^ image[15][1] + signed_kernel[2][1] ~^ image[15][2] + signed_kernel[2][2] ~^ image[15][3] + signed_kernel[2][3] ~^ image[15][4] + signed_kernel[2][4] ~^ image[15][5] + signed_kernel[3][0] ~^ image[16][1] + signed_kernel[3][1] ~^ image[16][2] + signed_kernel[3][2] ~^ image[16][3] + signed_kernel[3][3] ~^ image[16][4] + signed_kernel[3][4] ~^ image[16][5] + signed_kernel[4][0] ~^ image[17][1] + signed_kernel[4][1] ~^ image[17][2] + signed_kernel[4][2] ~^ image[17][3] + signed_kernel[4][3] ~^ image[17][4] + signed_kernel[4][4] ~^ image[17][5];
assign xor_sum[13][2] = signed_kernel[0][0] ~^ image[13][2] + signed_kernel[0][1] ~^ image[13][3] + signed_kernel[0][2] ~^ image[13][4] + signed_kernel[0][3] ~^ image[13][5] + signed_kernel[0][4] ~^ image[13][6] + signed_kernel[1][0] ~^ image[14][2] + signed_kernel[1][1] ~^ image[14][3] + signed_kernel[1][2] ~^ image[14][4] + signed_kernel[1][3] ~^ image[14][5] + signed_kernel[1][4] ~^ image[14][6] + signed_kernel[2][0] ~^ image[15][2] + signed_kernel[2][1] ~^ image[15][3] + signed_kernel[2][2] ~^ image[15][4] + signed_kernel[2][3] ~^ image[15][5] + signed_kernel[2][4] ~^ image[15][6] + signed_kernel[3][0] ~^ image[16][2] + signed_kernel[3][1] ~^ image[16][3] + signed_kernel[3][2] ~^ image[16][4] + signed_kernel[3][3] ~^ image[16][5] + signed_kernel[3][4] ~^ image[16][6] + signed_kernel[4][0] ~^ image[17][2] + signed_kernel[4][1] ~^ image[17][3] + signed_kernel[4][2] ~^ image[17][4] + signed_kernel[4][3] ~^ image[17][5] + signed_kernel[4][4] ~^ image[17][6];
assign xor_sum[13][3] = signed_kernel[0][0] ~^ image[13][3] + signed_kernel[0][1] ~^ image[13][4] + signed_kernel[0][2] ~^ image[13][5] + signed_kernel[0][3] ~^ image[13][6] + signed_kernel[0][4] ~^ image[13][7] + signed_kernel[1][0] ~^ image[14][3] + signed_kernel[1][1] ~^ image[14][4] + signed_kernel[1][2] ~^ image[14][5] + signed_kernel[1][3] ~^ image[14][6] + signed_kernel[1][4] ~^ image[14][7] + signed_kernel[2][0] ~^ image[15][3] + signed_kernel[2][1] ~^ image[15][4] + signed_kernel[2][2] ~^ image[15][5] + signed_kernel[2][3] ~^ image[15][6] + signed_kernel[2][4] ~^ image[15][7] + signed_kernel[3][0] ~^ image[16][3] + signed_kernel[3][1] ~^ image[16][4] + signed_kernel[3][2] ~^ image[16][5] + signed_kernel[3][3] ~^ image[16][6] + signed_kernel[3][4] ~^ image[16][7] + signed_kernel[4][0] ~^ image[17][3] + signed_kernel[4][1] ~^ image[17][4] + signed_kernel[4][2] ~^ image[17][5] + signed_kernel[4][3] ~^ image[17][6] + signed_kernel[4][4] ~^ image[17][7];
assign xor_sum[13][4] = signed_kernel[0][0] ~^ image[13][4] + signed_kernel[0][1] ~^ image[13][5] + signed_kernel[0][2] ~^ image[13][6] + signed_kernel[0][3] ~^ image[13][7] + signed_kernel[0][4] ~^ image[13][8] + signed_kernel[1][0] ~^ image[14][4] + signed_kernel[1][1] ~^ image[14][5] + signed_kernel[1][2] ~^ image[14][6] + signed_kernel[1][3] ~^ image[14][7] + signed_kernel[1][4] ~^ image[14][8] + signed_kernel[2][0] ~^ image[15][4] + signed_kernel[2][1] ~^ image[15][5] + signed_kernel[2][2] ~^ image[15][6] + signed_kernel[2][3] ~^ image[15][7] + signed_kernel[2][4] ~^ image[15][8] + signed_kernel[3][0] ~^ image[16][4] + signed_kernel[3][1] ~^ image[16][5] + signed_kernel[3][2] ~^ image[16][6] + signed_kernel[3][3] ~^ image[16][7] + signed_kernel[3][4] ~^ image[16][8] + signed_kernel[4][0] ~^ image[17][4] + signed_kernel[4][1] ~^ image[17][5] + signed_kernel[4][2] ~^ image[17][6] + signed_kernel[4][3] ~^ image[17][7] + signed_kernel[4][4] ~^ image[17][8];
assign xor_sum[13][5] = signed_kernel[0][0] ~^ image[13][5] + signed_kernel[0][1] ~^ image[13][6] + signed_kernel[0][2] ~^ image[13][7] + signed_kernel[0][3] ~^ image[13][8] + signed_kernel[0][4] ~^ image[13][9] + signed_kernel[1][0] ~^ image[14][5] + signed_kernel[1][1] ~^ image[14][6] + signed_kernel[1][2] ~^ image[14][7] + signed_kernel[1][3] ~^ image[14][8] + signed_kernel[1][4] ~^ image[14][9] + signed_kernel[2][0] ~^ image[15][5] + signed_kernel[2][1] ~^ image[15][6] + signed_kernel[2][2] ~^ image[15][7] + signed_kernel[2][3] ~^ image[15][8] + signed_kernel[2][4] ~^ image[15][9] + signed_kernel[3][0] ~^ image[16][5] + signed_kernel[3][1] ~^ image[16][6] + signed_kernel[3][2] ~^ image[16][7] + signed_kernel[3][3] ~^ image[16][8] + signed_kernel[3][4] ~^ image[16][9] + signed_kernel[4][0] ~^ image[17][5] + signed_kernel[4][1] ~^ image[17][6] + signed_kernel[4][2] ~^ image[17][7] + signed_kernel[4][3] ~^ image[17][8] + signed_kernel[4][4] ~^ image[17][9];
assign xor_sum[13][6] = signed_kernel[0][0] ~^ image[13][6] + signed_kernel[0][1] ~^ image[13][7] + signed_kernel[0][2] ~^ image[13][8] + signed_kernel[0][3] ~^ image[13][9] + signed_kernel[0][4] ~^ image[13][10] + signed_kernel[1][0] ~^ image[14][6] + signed_kernel[1][1] ~^ image[14][7] + signed_kernel[1][2] ~^ image[14][8] + signed_kernel[1][3] ~^ image[14][9] + signed_kernel[1][4] ~^ image[14][10] + signed_kernel[2][0] ~^ image[15][6] + signed_kernel[2][1] ~^ image[15][7] + signed_kernel[2][2] ~^ image[15][8] + signed_kernel[2][3] ~^ image[15][9] + signed_kernel[2][4] ~^ image[15][10] + signed_kernel[3][0] ~^ image[16][6] + signed_kernel[3][1] ~^ image[16][7] + signed_kernel[3][2] ~^ image[16][8] + signed_kernel[3][3] ~^ image[16][9] + signed_kernel[3][4] ~^ image[16][10] + signed_kernel[4][0] ~^ image[17][6] + signed_kernel[4][1] ~^ image[17][7] + signed_kernel[4][2] ~^ image[17][8] + signed_kernel[4][3] ~^ image[17][9] + signed_kernel[4][4] ~^ image[17][10];
assign xor_sum[13][7] = signed_kernel[0][0] ~^ image[13][7] + signed_kernel[0][1] ~^ image[13][8] + signed_kernel[0][2] ~^ image[13][9] + signed_kernel[0][3] ~^ image[13][10] + signed_kernel[0][4] ~^ image[13][11] + signed_kernel[1][0] ~^ image[14][7] + signed_kernel[1][1] ~^ image[14][8] + signed_kernel[1][2] ~^ image[14][9] + signed_kernel[1][3] ~^ image[14][10] + signed_kernel[1][4] ~^ image[14][11] + signed_kernel[2][0] ~^ image[15][7] + signed_kernel[2][1] ~^ image[15][8] + signed_kernel[2][2] ~^ image[15][9] + signed_kernel[2][3] ~^ image[15][10] + signed_kernel[2][4] ~^ image[15][11] + signed_kernel[3][0] ~^ image[16][7] + signed_kernel[3][1] ~^ image[16][8] + signed_kernel[3][2] ~^ image[16][9] + signed_kernel[3][3] ~^ image[16][10] + signed_kernel[3][4] ~^ image[16][11] + signed_kernel[4][0] ~^ image[17][7] + signed_kernel[4][1] ~^ image[17][8] + signed_kernel[4][2] ~^ image[17][9] + signed_kernel[4][3] ~^ image[17][10] + signed_kernel[4][4] ~^ image[17][11];
assign xor_sum[13][8] = signed_kernel[0][0] ~^ image[13][8] + signed_kernel[0][1] ~^ image[13][9] + signed_kernel[0][2] ~^ image[13][10] + signed_kernel[0][3] ~^ image[13][11] + signed_kernel[0][4] ~^ image[13][12] + signed_kernel[1][0] ~^ image[14][8] + signed_kernel[1][1] ~^ image[14][9] + signed_kernel[1][2] ~^ image[14][10] + signed_kernel[1][3] ~^ image[14][11] + signed_kernel[1][4] ~^ image[14][12] + signed_kernel[2][0] ~^ image[15][8] + signed_kernel[2][1] ~^ image[15][9] + signed_kernel[2][2] ~^ image[15][10] + signed_kernel[2][3] ~^ image[15][11] + signed_kernel[2][4] ~^ image[15][12] + signed_kernel[3][0] ~^ image[16][8] + signed_kernel[3][1] ~^ image[16][9] + signed_kernel[3][2] ~^ image[16][10] + signed_kernel[3][3] ~^ image[16][11] + signed_kernel[3][4] ~^ image[16][12] + signed_kernel[4][0] ~^ image[17][8] + signed_kernel[4][1] ~^ image[17][9] + signed_kernel[4][2] ~^ image[17][10] + signed_kernel[4][3] ~^ image[17][11] + signed_kernel[4][4] ~^ image[17][12];
assign xor_sum[13][9] = signed_kernel[0][0] ~^ image[13][9] + signed_kernel[0][1] ~^ image[13][10] + signed_kernel[0][2] ~^ image[13][11] + signed_kernel[0][3] ~^ image[13][12] + signed_kernel[0][4] ~^ image[13][13] + signed_kernel[1][0] ~^ image[14][9] + signed_kernel[1][1] ~^ image[14][10] + signed_kernel[1][2] ~^ image[14][11] + signed_kernel[1][3] ~^ image[14][12] + signed_kernel[1][4] ~^ image[14][13] + signed_kernel[2][0] ~^ image[15][9] + signed_kernel[2][1] ~^ image[15][10] + signed_kernel[2][2] ~^ image[15][11] + signed_kernel[2][3] ~^ image[15][12] + signed_kernel[2][4] ~^ image[15][13] + signed_kernel[3][0] ~^ image[16][9] + signed_kernel[3][1] ~^ image[16][10] + signed_kernel[3][2] ~^ image[16][11] + signed_kernel[3][3] ~^ image[16][12] + signed_kernel[3][4] ~^ image[16][13] + signed_kernel[4][0] ~^ image[17][9] + signed_kernel[4][1] ~^ image[17][10] + signed_kernel[4][2] ~^ image[17][11] + signed_kernel[4][3] ~^ image[17][12] + signed_kernel[4][4] ~^ image[17][13];
assign xor_sum[13][10] = signed_kernel[0][0] ~^ image[13][10] + signed_kernel[0][1] ~^ image[13][11] + signed_kernel[0][2] ~^ image[13][12] + signed_kernel[0][3] ~^ image[13][13] + signed_kernel[0][4] ~^ image[13][14] + signed_kernel[1][0] ~^ image[14][10] + signed_kernel[1][1] ~^ image[14][11] + signed_kernel[1][2] ~^ image[14][12] + signed_kernel[1][3] ~^ image[14][13] + signed_kernel[1][4] ~^ image[14][14] + signed_kernel[2][0] ~^ image[15][10] + signed_kernel[2][1] ~^ image[15][11] + signed_kernel[2][2] ~^ image[15][12] + signed_kernel[2][3] ~^ image[15][13] + signed_kernel[2][4] ~^ image[15][14] + signed_kernel[3][0] ~^ image[16][10] + signed_kernel[3][1] ~^ image[16][11] + signed_kernel[3][2] ~^ image[16][12] + signed_kernel[3][3] ~^ image[16][13] + signed_kernel[3][4] ~^ image[16][14] + signed_kernel[4][0] ~^ image[17][10] + signed_kernel[4][1] ~^ image[17][11] + signed_kernel[4][2] ~^ image[17][12] + signed_kernel[4][3] ~^ image[17][13] + signed_kernel[4][4] ~^ image[17][14];
assign xor_sum[13][11] = signed_kernel[0][0] ~^ image[13][11] + signed_kernel[0][1] ~^ image[13][12] + signed_kernel[0][2] ~^ image[13][13] + signed_kernel[0][3] ~^ image[13][14] + signed_kernel[0][4] ~^ image[13][15] + signed_kernel[1][0] ~^ image[14][11] + signed_kernel[1][1] ~^ image[14][12] + signed_kernel[1][2] ~^ image[14][13] + signed_kernel[1][3] ~^ image[14][14] + signed_kernel[1][4] ~^ image[14][15] + signed_kernel[2][0] ~^ image[15][11] + signed_kernel[2][1] ~^ image[15][12] + signed_kernel[2][2] ~^ image[15][13] + signed_kernel[2][3] ~^ image[15][14] + signed_kernel[2][4] ~^ image[15][15] + signed_kernel[3][0] ~^ image[16][11] + signed_kernel[3][1] ~^ image[16][12] + signed_kernel[3][2] ~^ image[16][13] + signed_kernel[3][3] ~^ image[16][14] + signed_kernel[3][4] ~^ image[16][15] + signed_kernel[4][0] ~^ image[17][11] + signed_kernel[4][1] ~^ image[17][12] + signed_kernel[4][2] ~^ image[17][13] + signed_kernel[4][3] ~^ image[17][14] + signed_kernel[4][4] ~^ image[17][15];
assign xor_sum[13][12] = signed_kernel[0][0] ~^ image[13][12] + signed_kernel[0][1] ~^ image[13][13] + signed_kernel[0][2] ~^ image[13][14] + signed_kernel[0][3] ~^ image[13][15] + signed_kernel[0][4] ~^ image[13][16] + signed_kernel[1][0] ~^ image[14][12] + signed_kernel[1][1] ~^ image[14][13] + signed_kernel[1][2] ~^ image[14][14] + signed_kernel[1][3] ~^ image[14][15] + signed_kernel[1][4] ~^ image[14][16] + signed_kernel[2][0] ~^ image[15][12] + signed_kernel[2][1] ~^ image[15][13] + signed_kernel[2][2] ~^ image[15][14] + signed_kernel[2][3] ~^ image[15][15] + signed_kernel[2][4] ~^ image[15][16] + signed_kernel[3][0] ~^ image[16][12] + signed_kernel[3][1] ~^ image[16][13] + signed_kernel[3][2] ~^ image[16][14] + signed_kernel[3][3] ~^ image[16][15] + signed_kernel[3][4] ~^ image[16][16] + signed_kernel[4][0] ~^ image[17][12] + signed_kernel[4][1] ~^ image[17][13] + signed_kernel[4][2] ~^ image[17][14] + signed_kernel[4][3] ~^ image[17][15] + signed_kernel[4][4] ~^ image[17][16];
assign xor_sum[13][13] = signed_kernel[0][0] ~^ image[13][13] + signed_kernel[0][1] ~^ image[13][14] + signed_kernel[0][2] ~^ image[13][15] + signed_kernel[0][3] ~^ image[13][16] + signed_kernel[0][4] ~^ image[13][17] + signed_kernel[1][0] ~^ image[14][13] + signed_kernel[1][1] ~^ image[14][14] + signed_kernel[1][2] ~^ image[14][15] + signed_kernel[1][3] ~^ image[14][16] + signed_kernel[1][4] ~^ image[14][17] + signed_kernel[2][0] ~^ image[15][13] + signed_kernel[2][1] ~^ image[15][14] + signed_kernel[2][2] ~^ image[15][15] + signed_kernel[2][3] ~^ image[15][16] + signed_kernel[2][4] ~^ image[15][17] + signed_kernel[3][0] ~^ image[16][13] + signed_kernel[3][1] ~^ image[16][14] + signed_kernel[3][2] ~^ image[16][15] + signed_kernel[3][3] ~^ image[16][16] + signed_kernel[3][4] ~^ image[16][17] + signed_kernel[4][0] ~^ image[17][13] + signed_kernel[4][1] ~^ image[17][14] + signed_kernel[4][2] ~^ image[17][15] + signed_kernel[4][3] ~^ image[17][16] + signed_kernel[4][4] ~^ image[17][17];
assign xor_sum[13][14] = signed_kernel[0][0] ~^ image[13][14] + signed_kernel[0][1] ~^ image[13][15] + signed_kernel[0][2] ~^ image[13][16] + signed_kernel[0][3] ~^ image[13][17] + signed_kernel[0][4] ~^ image[13][18] + signed_kernel[1][0] ~^ image[14][14] + signed_kernel[1][1] ~^ image[14][15] + signed_kernel[1][2] ~^ image[14][16] + signed_kernel[1][3] ~^ image[14][17] + signed_kernel[1][4] ~^ image[14][18] + signed_kernel[2][0] ~^ image[15][14] + signed_kernel[2][1] ~^ image[15][15] + signed_kernel[2][2] ~^ image[15][16] + signed_kernel[2][3] ~^ image[15][17] + signed_kernel[2][4] ~^ image[15][18] + signed_kernel[3][0] ~^ image[16][14] + signed_kernel[3][1] ~^ image[16][15] + signed_kernel[3][2] ~^ image[16][16] + signed_kernel[3][3] ~^ image[16][17] + signed_kernel[3][4] ~^ image[16][18] + signed_kernel[4][0] ~^ image[17][14] + signed_kernel[4][1] ~^ image[17][15] + signed_kernel[4][2] ~^ image[17][16] + signed_kernel[4][3] ~^ image[17][17] + signed_kernel[4][4] ~^ image[17][18];
assign xor_sum[13][15] = signed_kernel[0][0] ~^ image[13][15] + signed_kernel[0][1] ~^ image[13][16] + signed_kernel[0][2] ~^ image[13][17] + signed_kernel[0][3] ~^ image[13][18] + signed_kernel[0][4] ~^ image[13][19] + signed_kernel[1][0] ~^ image[14][15] + signed_kernel[1][1] ~^ image[14][16] + signed_kernel[1][2] ~^ image[14][17] + signed_kernel[1][3] ~^ image[14][18] + signed_kernel[1][4] ~^ image[14][19] + signed_kernel[2][0] ~^ image[15][15] + signed_kernel[2][1] ~^ image[15][16] + signed_kernel[2][2] ~^ image[15][17] + signed_kernel[2][3] ~^ image[15][18] + signed_kernel[2][4] ~^ image[15][19] + signed_kernel[3][0] ~^ image[16][15] + signed_kernel[3][1] ~^ image[16][16] + signed_kernel[3][2] ~^ image[16][17] + signed_kernel[3][3] ~^ image[16][18] + signed_kernel[3][4] ~^ image[16][19] + signed_kernel[4][0] ~^ image[17][15] + signed_kernel[4][1] ~^ image[17][16] + signed_kernel[4][2] ~^ image[17][17] + signed_kernel[4][3] ~^ image[17][18] + signed_kernel[4][4] ~^ image[17][19];
assign xor_sum[13][16] = signed_kernel[0][0] ~^ image[13][16] + signed_kernel[0][1] ~^ image[13][17] + signed_kernel[0][2] ~^ image[13][18] + signed_kernel[0][3] ~^ image[13][19] + signed_kernel[0][4] ~^ image[13][20] + signed_kernel[1][0] ~^ image[14][16] + signed_kernel[1][1] ~^ image[14][17] + signed_kernel[1][2] ~^ image[14][18] + signed_kernel[1][3] ~^ image[14][19] + signed_kernel[1][4] ~^ image[14][20] + signed_kernel[2][0] ~^ image[15][16] + signed_kernel[2][1] ~^ image[15][17] + signed_kernel[2][2] ~^ image[15][18] + signed_kernel[2][3] ~^ image[15][19] + signed_kernel[2][4] ~^ image[15][20] + signed_kernel[3][0] ~^ image[16][16] + signed_kernel[3][1] ~^ image[16][17] + signed_kernel[3][2] ~^ image[16][18] + signed_kernel[3][3] ~^ image[16][19] + signed_kernel[3][4] ~^ image[16][20] + signed_kernel[4][0] ~^ image[17][16] + signed_kernel[4][1] ~^ image[17][17] + signed_kernel[4][2] ~^ image[17][18] + signed_kernel[4][3] ~^ image[17][19] + signed_kernel[4][4] ~^ image[17][20];
assign xor_sum[13][17] = signed_kernel[0][0] ~^ image[13][17] + signed_kernel[0][1] ~^ image[13][18] + signed_kernel[0][2] ~^ image[13][19] + signed_kernel[0][3] ~^ image[13][20] + signed_kernel[0][4] ~^ image[13][21] + signed_kernel[1][0] ~^ image[14][17] + signed_kernel[1][1] ~^ image[14][18] + signed_kernel[1][2] ~^ image[14][19] + signed_kernel[1][3] ~^ image[14][20] + signed_kernel[1][4] ~^ image[14][21] + signed_kernel[2][0] ~^ image[15][17] + signed_kernel[2][1] ~^ image[15][18] + signed_kernel[2][2] ~^ image[15][19] + signed_kernel[2][3] ~^ image[15][20] + signed_kernel[2][4] ~^ image[15][21] + signed_kernel[3][0] ~^ image[16][17] + signed_kernel[3][1] ~^ image[16][18] + signed_kernel[3][2] ~^ image[16][19] + signed_kernel[3][3] ~^ image[16][20] + signed_kernel[3][4] ~^ image[16][21] + signed_kernel[4][0] ~^ image[17][17] + signed_kernel[4][1] ~^ image[17][18] + signed_kernel[4][2] ~^ image[17][19] + signed_kernel[4][3] ~^ image[17][20] + signed_kernel[4][4] ~^ image[17][21];
assign xor_sum[13][18] = signed_kernel[0][0] ~^ image[13][18] + signed_kernel[0][1] ~^ image[13][19] + signed_kernel[0][2] ~^ image[13][20] + signed_kernel[0][3] ~^ image[13][21] + signed_kernel[0][4] ~^ image[13][22] + signed_kernel[1][0] ~^ image[14][18] + signed_kernel[1][1] ~^ image[14][19] + signed_kernel[1][2] ~^ image[14][20] + signed_kernel[1][3] ~^ image[14][21] + signed_kernel[1][4] ~^ image[14][22] + signed_kernel[2][0] ~^ image[15][18] + signed_kernel[2][1] ~^ image[15][19] + signed_kernel[2][2] ~^ image[15][20] + signed_kernel[2][3] ~^ image[15][21] + signed_kernel[2][4] ~^ image[15][22] + signed_kernel[3][0] ~^ image[16][18] + signed_kernel[3][1] ~^ image[16][19] + signed_kernel[3][2] ~^ image[16][20] + signed_kernel[3][3] ~^ image[16][21] + signed_kernel[3][4] ~^ image[16][22] + signed_kernel[4][0] ~^ image[17][18] + signed_kernel[4][1] ~^ image[17][19] + signed_kernel[4][2] ~^ image[17][20] + signed_kernel[4][3] ~^ image[17][21] + signed_kernel[4][4] ~^ image[17][22];
assign xor_sum[13][19] = signed_kernel[0][0] ~^ image[13][19] + signed_kernel[0][1] ~^ image[13][20] + signed_kernel[0][2] ~^ image[13][21] + signed_kernel[0][3] ~^ image[13][22] + signed_kernel[0][4] ~^ image[13][23] + signed_kernel[1][0] ~^ image[14][19] + signed_kernel[1][1] ~^ image[14][20] + signed_kernel[1][2] ~^ image[14][21] + signed_kernel[1][3] ~^ image[14][22] + signed_kernel[1][4] ~^ image[14][23] + signed_kernel[2][0] ~^ image[15][19] + signed_kernel[2][1] ~^ image[15][20] + signed_kernel[2][2] ~^ image[15][21] + signed_kernel[2][3] ~^ image[15][22] + signed_kernel[2][4] ~^ image[15][23] + signed_kernel[3][0] ~^ image[16][19] + signed_kernel[3][1] ~^ image[16][20] + signed_kernel[3][2] ~^ image[16][21] + signed_kernel[3][3] ~^ image[16][22] + signed_kernel[3][4] ~^ image[16][23] + signed_kernel[4][0] ~^ image[17][19] + signed_kernel[4][1] ~^ image[17][20] + signed_kernel[4][2] ~^ image[17][21] + signed_kernel[4][3] ~^ image[17][22] + signed_kernel[4][4] ~^ image[17][23];
assign xor_sum[13][20] = signed_kernel[0][0] ~^ image[13][20] + signed_kernel[0][1] ~^ image[13][21] + signed_kernel[0][2] ~^ image[13][22] + signed_kernel[0][3] ~^ image[13][23] + signed_kernel[0][4] ~^ image[13][24] + signed_kernel[1][0] ~^ image[14][20] + signed_kernel[1][1] ~^ image[14][21] + signed_kernel[1][2] ~^ image[14][22] + signed_kernel[1][3] ~^ image[14][23] + signed_kernel[1][4] ~^ image[14][24] + signed_kernel[2][0] ~^ image[15][20] + signed_kernel[2][1] ~^ image[15][21] + signed_kernel[2][2] ~^ image[15][22] + signed_kernel[2][3] ~^ image[15][23] + signed_kernel[2][4] ~^ image[15][24] + signed_kernel[3][0] ~^ image[16][20] + signed_kernel[3][1] ~^ image[16][21] + signed_kernel[3][2] ~^ image[16][22] + signed_kernel[3][3] ~^ image[16][23] + signed_kernel[3][4] ~^ image[16][24] + signed_kernel[4][0] ~^ image[17][20] + signed_kernel[4][1] ~^ image[17][21] + signed_kernel[4][2] ~^ image[17][22] + signed_kernel[4][3] ~^ image[17][23] + signed_kernel[4][4] ~^ image[17][24];
assign xor_sum[13][21] = signed_kernel[0][0] ~^ image[13][21] + signed_kernel[0][1] ~^ image[13][22] + signed_kernel[0][2] ~^ image[13][23] + signed_kernel[0][3] ~^ image[13][24] + signed_kernel[0][4] ~^ image[13][25] + signed_kernel[1][0] ~^ image[14][21] + signed_kernel[1][1] ~^ image[14][22] + signed_kernel[1][2] ~^ image[14][23] + signed_kernel[1][3] ~^ image[14][24] + signed_kernel[1][4] ~^ image[14][25] + signed_kernel[2][0] ~^ image[15][21] + signed_kernel[2][1] ~^ image[15][22] + signed_kernel[2][2] ~^ image[15][23] + signed_kernel[2][3] ~^ image[15][24] + signed_kernel[2][4] ~^ image[15][25] + signed_kernel[3][0] ~^ image[16][21] + signed_kernel[3][1] ~^ image[16][22] + signed_kernel[3][2] ~^ image[16][23] + signed_kernel[3][3] ~^ image[16][24] + signed_kernel[3][4] ~^ image[16][25] + signed_kernel[4][0] ~^ image[17][21] + signed_kernel[4][1] ~^ image[17][22] + signed_kernel[4][2] ~^ image[17][23] + signed_kernel[4][3] ~^ image[17][24] + signed_kernel[4][4] ~^ image[17][25];
assign xor_sum[13][22] = signed_kernel[0][0] ~^ image[13][22] + signed_kernel[0][1] ~^ image[13][23] + signed_kernel[0][2] ~^ image[13][24] + signed_kernel[0][3] ~^ image[13][25] + signed_kernel[0][4] ~^ image[13][26] + signed_kernel[1][0] ~^ image[14][22] + signed_kernel[1][1] ~^ image[14][23] + signed_kernel[1][2] ~^ image[14][24] + signed_kernel[1][3] ~^ image[14][25] + signed_kernel[1][4] ~^ image[14][26] + signed_kernel[2][0] ~^ image[15][22] + signed_kernel[2][1] ~^ image[15][23] + signed_kernel[2][2] ~^ image[15][24] + signed_kernel[2][3] ~^ image[15][25] + signed_kernel[2][4] ~^ image[15][26] + signed_kernel[3][0] ~^ image[16][22] + signed_kernel[3][1] ~^ image[16][23] + signed_kernel[3][2] ~^ image[16][24] + signed_kernel[3][3] ~^ image[16][25] + signed_kernel[3][4] ~^ image[16][26] + signed_kernel[4][0] ~^ image[17][22] + signed_kernel[4][1] ~^ image[17][23] + signed_kernel[4][2] ~^ image[17][24] + signed_kernel[4][3] ~^ image[17][25] + signed_kernel[4][4] ~^ image[17][26];
assign xor_sum[13][23] = signed_kernel[0][0] ~^ image[13][23] + signed_kernel[0][1] ~^ image[13][24] + signed_kernel[0][2] ~^ image[13][25] + signed_kernel[0][3] ~^ image[13][26] + signed_kernel[0][4] ~^ image[13][27] + signed_kernel[1][0] ~^ image[14][23] + signed_kernel[1][1] ~^ image[14][24] + signed_kernel[1][2] ~^ image[14][25] + signed_kernel[1][3] ~^ image[14][26] + signed_kernel[1][4] ~^ image[14][27] + signed_kernel[2][0] ~^ image[15][23] + signed_kernel[2][1] ~^ image[15][24] + signed_kernel[2][2] ~^ image[15][25] + signed_kernel[2][3] ~^ image[15][26] + signed_kernel[2][4] ~^ image[15][27] + signed_kernel[3][0] ~^ image[16][23] + signed_kernel[3][1] ~^ image[16][24] + signed_kernel[3][2] ~^ image[16][25] + signed_kernel[3][3] ~^ image[16][26] + signed_kernel[3][4] ~^ image[16][27] + signed_kernel[4][0] ~^ image[17][23] + signed_kernel[4][1] ~^ image[17][24] + signed_kernel[4][2] ~^ image[17][25] + signed_kernel[4][3] ~^ image[17][26] + signed_kernel[4][4] ~^ image[17][27];
assign xor_sum[14][0] = signed_kernel[0][0] ~^ image[14][0] + signed_kernel[0][1] ~^ image[14][1] + signed_kernel[0][2] ~^ image[14][2] + signed_kernel[0][3] ~^ image[14][3] + signed_kernel[0][4] ~^ image[14][4] + signed_kernel[1][0] ~^ image[15][0] + signed_kernel[1][1] ~^ image[15][1] + signed_kernel[1][2] ~^ image[15][2] + signed_kernel[1][3] ~^ image[15][3] + signed_kernel[1][4] ~^ image[15][4] + signed_kernel[2][0] ~^ image[16][0] + signed_kernel[2][1] ~^ image[16][1] + signed_kernel[2][2] ~^ image[16][2] + signed_kernel[2][3] ~^ image[16][3] + signed_kernel[2][4] ~^ image[16][4] + signed_kernel[3][0] ~^ image[17][0] + signed_kernel[3][1] ~^ image[17][1] + signed_kernel[3][2] ~^ image[17][2] + signed_kernel[3][3] ~^ image[17][3] + signed_kernel[3][4] ~^ image[17][4] + signed_kernel[4][0] ~^ image[18][0] + signed_kernel[4][1] ~^ image[18][1] + signed_kernel[4][2] ~^ image[18][2] + signed_kernel[4][3] ~^ image[18][3] + signed_kernel[4][4] ~^ image[18][4];
assign xor_sum[14][1] = signed_kernel[0][0] ~^ image[14][1] + signed_kernel[0][1] ~^ image[14][2] + signed_kernel[0][2] ~^ image[14][3] + signed_kernel[0][3] ~^ image[14][4] + signed_kernel[0][4] ~^ image[14][5] + signed_kernel[1][0] ~^ image[15][1] + signed_kernel[1][1] ~^ image[15][2] + signed_kernel[1][2] ~^ image[15][3] + signed_kernel[1][3] ~^ image[15][4] + signed_kernel[1][4] ~^ image[15][5] + signed_kernel[2][0] ~^ image[16][1] + signed_kernel[2][1] ~^ image[16][2] + signed_kernel[2][2] ~^ image[16][3] + signed_kernel[2][3] ~^ image[16][4] + signed_kernel[2][4] ~^ image[16][5] + signed_kernel[3][0] ~^ image[17][1] + signed_kernel[3][1] ~^ image[17][2] + signed_kernel[3][2] ~^ image[17][3] + signed_kernel[3][3] ~^ image[17][4] + signed_kernel[3][4] ~^ image[17][5] + signed_kernel[4][0] ~^ image[18][1] + signed_kernel[4][1] ~^ image[18][2] + signed_kernel[4][2] ~^ image[18][3] + signed_kernel[4][3] ~^ image[18][4] + signed_kernel[4][4] ~^ image[18][5];
assign xor_sum[14][2] = signed_kernel[0][0] ~^ image[14][2] + signed_kernel[0][1] ~^ image[14][3] + signed_kernel[0][2] ~^ image[14][4] + signed_kernel[0][3] ~^ image[14][5] + signed_kernel[0][4] ~^ image[14][6] + signed_kernel[1][0] ~^ image[15][2] + signed_kernel[1][1] ~^ image[15][3] + signed_kernel[1][2] ~^ image[15][4] + signed_kernel[1][3] ~^ image[15][5] + signed_kernel[1][4] ~^ image[15][6] + signed_kernel[2][0] ~^ image[16][2] + signed_kernel[2][1] ~^ image[16][3] + signed_kernel[2][2] ~^ image[16][4] + signed_kernel[2][3] ~^ image[16][5] + signed_kernel[2][4] ~^ image[16][6] + signed_kernel[3][0] ~^ image[17][2] + signed_kernel[3][1] ~^ image[17][3] + signed_kernel[3][2] ~^ image[17][4] + signed_kernel[3][3] ~^ image[17][5] + signed_kernel[3][4] ~^ image[17][6] + signed_kernel[4][0] ~^ image[18][2] + signed_kernel[4][1] ~^ image[18][3] + signed_kernel[4][2] ~^ image[18][4] + signed_kernel[4][3] ~^ image[18][5] + signed_kernel[4][4] ~^ image[18][6];
assign xor_sum[14][3] = signed_kernel[0][0] ~^ image[14][3] + signed_kernel[0][1] ~^ image[14][4] + signed_kernel[0][2] ~^ image[14][5] + signed_kernel[0][3] ~^ image[14][6] + signed_kernel[0][4] ~^ image[14][7] + signed_kernel[1][0] ~^ image[15][3] + signed_kernel[1][1] ~^ image[15][4] + signed_kernel[1][2] ~^ image[15][5] + signed_kernel[1][3] ~^ image[15][6] + signed_kernel[1][4] ~^ image[15][7] + signed_kernel[2][0] ~^ image[16][3] + signed_kernel[2][1] ~^ image[16][4] + signed_kernel[2][2] ~^ image[16][5] + signed_kernel[2][3] ~^ image[16][6] + signed_kernel[2][4] ~^ image[16][7] + signed_kernel[3][0] ~^ image[17][3] + signed_kernel[3][1] ~^ image[17][4] + signed_kernel[3][2] ~^ image[17][5] + signed_kernel[3][3] ~^ image[17][6] + signed_kernel[3][4] ~^ image[17][7] + signed_kernel[4][0] ~^ image[18][3] + signed_kernel[4][1] ~^ image[18][4] + signed_kernel[4][2] ~^ image[18][5] + signed_kernel[4][3] ~^ image[18][6] + signed_kernel[4][4] ~^ image[18][7];
assign xor_sum[14][4] = signed_kernel[0][0] ~^ image[14][4] + signed_kernel[0][1] ~^ image[14][5] + signed_kernel[0][2] ~^ image[14][6] + signed_kernel[0][3] ~^ image[14][7] + signed_kernel[0][4] ~^ image[14][8] + signed_kernel[1][0] ~^ image[15][4] + signed_kernel[1][1] ~^ image[15][5] + signed_kernel[1][2] ~^ image[15][6] + signed_kernel[1][3] ~^ image[15][7] + signed_kernel[1][4] ~^ image[15][8] + signed_kernel[2][0] ~^ image[16][4] + signed_kernel[2][1] ~^ image[16][5] + signed_kernel[2][2] ~^ image[16][6] + signed_kernel[2][3] ~^ image[16][7] + signed_kernel[2][4] ~^ image[16][8] + signed_kernel[3][0] ~^ image[17][4] + signed_kernel[3][1] ~^ image[17][5] + signed_kernel[3][2] ~^ image[17][6] + signed_kernel[3][3] ~^ image[17][7] + signed_kernel[3][4] ~^ image[17][8] + signed_kernel[4][0] ~^ image[18][4] + signed_kernel[4][1] ~^ image[18][5] + signed_kernel[4][2] ~^ image[18][6] + signed_kernel[4][3] ~^ image[18][7] + signed_kernel[4][4] ~^ image[18][8];
assign xor_sum[14][5] = signed_kernel[0][0] ~^ image[14][5] + signed_kernel[0][1] ~^ image[14][6] + signed_kernel[0][2] ~^ image[14][7] + signed_kernel[0][3] ~^ image[14][8] + signed_kernel[0][4] ~^ image[14][9] + signed_kernel[1][0] ~^ image[15][5] + signed_kernel[1][1] ~^ image[15][6] + signed_kernel[1][2] ~^ image[15][7] + signed_kernel[1][3] ~^ image[15][8] + signed_kernel[1][4] ~^ image[15][9] + signed_kernel[2][0] ~^ image[16][5] + signed_kernel[2][1] ~^ image[16][6] + signed_kernel[2][2] ~^ image[16][7] + signed_kernel[2][3] ~^ image[16][8] + signed_kernel[2][4] ~^ image[16][9] + signed_kernel[3][0] ~^ image[17][5] + signed_kernel[3][1] ~^ image[17][6] + signed_kernel[3][2] ~^ image[17][7] + signed_kernel[3][3] ~^ image[17][8] + signed_kernel[3][4] ~^ image[17][9] + signed_kernel[4][0] ~^ image[18][5] + signed_kernel[4][1] ~^ image[18][6] + signed_kernel[4][2] ~^ image[18][7] + signed_kernel[4][3] ~^ image[18][8] + signed_kernel[4][4] ~^ image[18][9];
assign xor_sum[14][6] = signed_kernel[0][0] ~^ image[14][6] + signed_kernel[0][1] ~^ image[14][7] + signed_kernel[0][2] ~^ image[14][8] + signed_kernel[0][3] ~^ image[14][9] + signed_kernel[0][4] ~^ image[14][10] + signed_kernel[1][0] ~^ image[15][6] + signed_kernel[1][1] ~^ image[15][7] + signed_kernel[1][2] ~^ image[15][8] + signed_kernel[1][3] ~^ image[15][9] + signed_kernel[1][4] ~^ image[15][10] + signed_kernel[2][0] ~^ image[16][6] + signed_kernel[2][1] ~^ image[16][7] + signed_kernel[2][2] ~^ image[16][8] + signed_kernel[2][3] ~^ image[16][9] + signed_kernel[2][4] ~^ image[16][10] + signed_kernel[3][0] ~^ image[17][6] + signed_kernel[3][1] ~^ image[17][7] + signed_kernel[3][2] ~^ image[17][8] + signed_kernel[3][3] ~^ image[17][9] + signed_kernel[3][4] ~^ image[17][10] + signed_kernel[4][0] ~^ image[18][6] + signed_kernel[4][1] ~^ image[18][7] + signed_kernel[4][2] ~^ image[18][8] + signed_kernel[4][3] ~^ image[18][9] + signed_kernel[4][4] ~^ image[18][10];
assign xor_sum[14][7] = signed_kernel[0][0] ~^ image[14][7] + signed_kernel[0][1] ~^ image[14][8] + signed_kernel[0][2] ~^ image[14][9] + signed_kernel[0][3] ~^ image[14][10] + signed_kernel[0][4] ~^ image[14][11] + signed_kernel[1][0] ~^ image[15][7] + signed_kernel[1][1] ~^ image[15][8] + signed_kernel[1][2] ~^ image[15][9] + signed_kernel[1][3] ~^ image[15][10] + signed_kernel[1][4] ~^ image[15][11] + signed_kernel[2][0] ~^ image[16][7] + signed_kernel[2][1] ~^ image[16][8] + signed_kernel[2][2] ~^ image[16][9] + signed_kernel[2][3] ~^ image[16][10] + signed_kernel[2][4] ~^ image[16][11] + signed_kernel[3][0] ~^ image[17][7] + signed_kernel[3][1] ~^ image[17][8] + signed_kernel[3][2] ~^ image[17][9] + signed_kernel[3][3] ~^ image[17][10] + signed_kernel[3][4] ~^ image[17][11] + signed_kernel[4][0] ~^ image[18][7] + signed_kernel[4][1] ~^ image[18][8] + signed_kernel[4][2] ~^ image[18][9] + signed_kernel[4][3] ~^ image[18][10] + signed_kernel[4][4] ~^ image[18][11];
assign xor_sum[14][8] = signed_kernel[0][0] ~^ image[14][8] + signed_kernel[0][1] ~^ image[14][9] + signed_kernel[0][2] ~^ image[14][10] + signed_kernel[0][3] ~^ image[14][11] + signed_kernel[0][4] ~^ image[14][12] + signed_kernel[1][0] ~^ image[15][8] + signed_kernel[1][1] ~^ image[15][9] + signed_kernel[1][2] ~^ image[15][10] + signed_kernel[1][3] ~^ image[15][11] + signed_kernel[1][4] ~^ image[15][12] + signed_kernel[2][0] ~^ image[16][8] + signed_kernel[2][1] ~^ image[16][9] + signed_kernel[2][2] ~^ image[16][10] + signed_kernel[2][3] ~^ image[16][11] + signed_kernel[2][4] ~^ image[16][12] + signed_kernel[3][0] ~^ image[17][8] + signed_kernel[3][1] ~^ image[17][9] + signed_kernel[3][2] ~^ image[17][10] + signed_kernel[3][3] ~^ image[17][11] + signed_kernel[3][4] ~^ image[17][12] + signed_kernel[4][0] ~^ image[18][8] + signed_kernel[4][1] ~^ image[18][9] + signed_kernel[4][2] ~^ image[18][10] + signed_kernel[4][3] ~^ image[18][11] + signed_kernel[4][4] ~^ image[18][12];
assign xor_sum[14][9] = signed_kernel[0][0] ~^ image[14][9] + signed_kernel[0][1] ~^ image[14][10] + signed_kernel[0][2] ~^ image[14][11] + signed_kernel[0][3] ~^ image[14][12] + signed_kernel[0][4] ~^ image[14][13] + signed_kernel[1][0] ~^ image[15][9] + signed_kernel[1][1] ~^ image[15][10] + signed_kernel[1][2] ~^ image[15][11] + signed_kernel[1][3] ~^ image[15][12] + signed_kernel[1][4] ~^ image[15][13] + signed_kernel[2][0] ~^ image[16][9] + signed_kernel[2][1] ~^ image[16][10] + signed_kernel[2][2] ~^ image[16][11] + signed_kernel[2][3] ~^ image[16][12] + signed_kernel[2][4] ~^ image[16][13] + signed_kernel[3][0] ~^ image[17][9] + signed_kernel[3][1] ~^ image[17][10] + signed_kernel[3][2] ~^ image[17][11] + signed_kernel[3][3] ~^ image[17][12] + signed_kernel[3][4] ~^ image[17][13] + signed_kernel[4][0] ~^ image[18][9] + signed_kernel[4][1] ~^ image[18][10] + signed_kernel[4][2] ~^ image[18][11] + signed_kernel[4][3] ~^ image[18][12] + signed_kernel[4][4] ~^ image[18][13];
assign xor_sum[14][10] = signed_kernel[0][0] ~^ image[14][10] + signed_kernel[0][1] ~^ image[14][11] + signed_kernel[0][2] ~^ image[14][12] + signed_kernel[0][3] ~^ image[14][13] + signed_kernel[0][4] ~^ image[14][14] + signed_kernel[1][0] ~^ image[15][10] + signed_kernel[1][1] ~^ image[15][11] + signed_kernel[1][2] ~^ image[15][12] + signed_kernel[1][3] ~^ image[15][13] + signed_kernel[1][4] ~^ image[15][14] + signed_kernel[2][0] ~^ image[16][10] + signed_kernel[2][1] ~^ image[16][11] + signed_kernel[2][2] ~^ image[16][12] + signed_kernel[2][3] ~^ image[16][13] + signed_kernel[2][4] ~^ image[16][14] + signed_kernel[3][0] ~^ image[17][10] + signed_kernel[3][1] ~^ image[17][11] + signed_kernel[3][2] ~^ image[17][12] + signed_kernel[3][3] ~^ image[17][13] + signed_kernel[3][4] ~^ image[17][14] + signed_kernel[4][0] ~^ image[18][10] + signed_kernel[4][1] ~^ image[18][11] + signed_kernel[4][2] ~^ image[18][12] + signed_kernel[4][3] ~^ image[18][13] + signed_kernel[4][4] ~^ image[18][14];
assign xor_sum[14][11] = signed_kernel[0][0] ~^ image[14][11] + signed_kernel[0][1] ~^ image[14][12] + signed_kernel[0][2] ~^ image[14][13] + signed_kernel[0][3] ~^ image[14][14] + signed_kernel[0][4] ~^ image[14][15] + signed_kernel[1][0] ~^ image[15][11] + signed_kernel[1][1] ~^ image[15][12] + signed_kernel[1][2] ~^ image[15][13] + signed_kernel[1][3] ~^ image[15][14] + signed_kernel[1][4] ~^ image[15][15] + signed_kernel[2][0] ~^ image[16][11] + signed_kernel[2][1] ~^ image[16][12] + signed_kernel[2][2] ~^ image[16][13] + signed_kernel[2][3] ~^ image[16][14] + signed_kernel[2][4] ~^ image[16][15] + signed_kernel[3][0] ~^ image[17][11] + signed_kernel[3][1] ~^ image[17][12] + signed_kernel[3][2] ~^ image[17][13] + signed_kernel[3][3] ~^ image[17][14] + signed_kernel[3][4] ~^ image[17][15] + signed_kernel[4][0] ~^ image[18][11] + signed_kernel[4][1] ~^ image[18][12] + signed_kernel[4][2] ~^ image[18][13] + signed_kernel[4][3] ~^ image[18][14] + signed_kernel[4][4] ~^ image[18][15];
assign xor_sum[14][12] = signed_kernel[0][0] ~^ image[14][12] + signed_kernel[0][1] ~^ image[14][13] + signed_kernel[0][2] ~^ image[14][14] + signed_kernel[0][3] ~^ image[14][15] + signed_kernel[0][4] ~^ image[14][16] + signed_kernel[1][0] ~^ image[15][12] + signed_kernel[1][1] ~^ image[15][13] + signed_kernel[1][2] ~^ image[15][14] + signed_kernel[1][3] ~^ image[15][15] + signed_kernel[1][4] ~^ image[15][16] + signed_kernel[2][0] ~^ image[16][12] + signed_kernel[2][1] ~^ image[16][13] + signed_kernel[2][2] ~^ image[16][14] + signed_kernel[2][3] ~^ image[16][15] + signed_kernel[2][4] ~^ image[16][16] + signed_kernel[3][0] ~^ image[17][12] + signed_kernel[3][1] ~^ image[17][13] + signed_kernel[3][2] ~^ image[17][14] + signed_kernel[3][3] ~^ image[17][15] + signed_kernel[3][4] ~^ image[17][16] + signed_kernel[4][0] ~^ image[18][12] + signed_kernel[4][1] ~^ image[18][13] + signed_kernel[4][2] ~^ image[18][14] + signed_kernel[4][3] ~^ image[18][15] + signed_kernel[4][4] ~^ image[18][16];
assign xor_sum[14][13] = signed_kernel[0][0] ~^ image[14][13] + signed_kernel[0][1] ~^ image[14][14] + signed_kernel[0][2] ~^ image[14][15] + signed_kernel[0][3] ~^ image[14][16] + signed_kernel[0][4] ~^ image[14][17] + signed_kernel[1][0] ~^ image[15][13] + signed_kernel[1][1] ~^ image[15][14] + signed_kernel[1][2] ~^ image[15][15] + signed_kernel[1][3] ~^ image[15][16] + signed_kernel[1][4] ~^ image[15][17] + signed_kernel[2][0] ~^ image[16][13] + signed_kernel[2][1] ~^ image[16][14] + signed_kernel[2][2] ~^ image[16][15] + signed_kernel[2][3] ~^ image[16][16] + signed_kernel[2][4] ~^ image[16][17] + signed_kernel[3][0] ~^ image[17][13] + signed_kernel[3][1] ~^ image[17][14] + signed_kernel[3][2] ~^ image[17][15] + signed_kernel[3][3] ~^ image[17][16] + signed_kernel[3][4] ~^ image[17][17] + signed_kernel[4][0] ~^ image[18][13] + signed_kernel[4][1] ~^ image[18][14] + signed_kernel[4][2] ~^ image[18][15] + signed_kernel[4][3] ~^ image[18][16] + signed_kernel[4][4] ~^ image[18][17];
assign xor_sum[14][14] = signed_kernel[0][0] ~^ image[14][14] + signed_kernel[0][1] ~^ image[14][15] + signed_kernel[0][2] ~^ image[14][16] + signed_kernel[0][3] ~^ image[14][17] + signed_kernel[0][4] ~^ image[14][18] + signed_kernel[1][0] ~^ image[15][14] + signed_kernel[1][1] ~^ image[15][15] + signed_kernel[1][2] ~^ image[15][16] + signed_kernel[1][3] ~^ image[15][17] + signed_kernel[1][4] ~^ image[15][18] + signed_kernel[2][0] ~^ image[16][14] + signed_kernel[2][1] ~^ image[16][15] + signed_kernel[2][2] ~^ image[16][16] + signed_kernel[2][3] ~^ image[16][17] + signed_kernel[2][4] ~^ image[16][18] + signed_kernel[3][0] ~^ image[17][14] + signed_kernel[3][1] ~^ image[17][15] + signed_kernel[3][2] ~^ image[17][16] + signed_kernel[3][3] ~^ image[17][17] + signed_kernel[3][4] ~^ image[17][18] + signed_kernel[4][0] ~^ image[18][14] + signed_kernel[4][1] ~^ image[18][15] + signed_kernel[4][2] ~^ image[18][16] + signed_kernel[4][3] ~^ image[18][17] + signed_kernel[4][4] ~^ image[18][18];
assign xor_sum[14][15] = signed_kernel[0][0] ~^ image[14][15] + signed_kernel[0][1] ~^ image[14][16] + signed_kernel[0][2] ~^ image[14][17] + signed_kernel[0][3] ~^ image[14][18] + signed_kernel[0][4] ~^ image[14][19] + signed_kernel[1][0] ~^ image[15][15] + signed_kernel[1][1] ~^ image[15][16] + signed_kernel[1][2] ~^ image[15][17] + signed_kernel[1][3] ~^ image[15][18] + signed_kernel[1][4] ~^ image[15][19] + signed_kernel[2][0] ~^ image[16][15] + signed_kernel[2][1] ~^ image[16][16] + signed_kernel[2][2] ~^ image[16][17] + signed_kernel[2][3] ~^ image[16][18] + signed_kernel[2][4] ~^ image[16][19] + signed_kernel[3][0] ~^ image[17][15] + signed_kernel[3][1] ~^ image[17][16] + signed_kernel[3][2] ~^ image[17][17] + signed_kernel[3][3] ~^ image[17][18] + signed_kernel[3][4] ~^ image[17][19] + signed_kernel[4][0] ~^ image[18][15] + signed_kernel[4][1] ~^ image[18][16] + signed_kernel[4][2] ~^ image[18][17] + signed_kernel[4][3] ~^ image[18][18] + signed_kernel[4][4] ~^ image[18][19];
assign xor_sum[14][16] = signed_kernel[0][0] ~^ image[14][16] + signed_kernel[0][1] ~^ image[14][17] + signed_kernel[0][2] ~^ image[14][18] + signed_kernel[0][3] ~^ image[14][19] + signed_kernel[0][4] ~^ image[14][20] + signed_kernel[1][0] ~^ image[15][16] + signed_kernel[1][1] ~^ image[15][17] + signed_kernel[1][2] ~^ image[15][18] + signed_kernel[1][3] ~^ image[15][19] + signed_kernel[1][4] ~^ image[15][20] + signed_kernel[2][0] ~^ image[16][16] + signed_kernel[2][1] ~^ image[16][17] + signed_kernel[2][2] ~^ image[16][18] + signed_kernel[2][3] ~^ image[16][19] + signed_kernel[2][4] ~^ image[16][20] + signed_kernel[3][0] ~^ image[17][16] + signed_kernel[3][1] ~^ image[17][17] + signed_kernel[3][2] ~^ image[17][18] + signed_kernel[3][3] ~^ image[17][19] + signed_kernel[3][4] ~^ image[17][20] + signed_kernel[4][0] ~^ image[18][16] + signed_kernel[4][1] ~^ image[18][17] + signed_kernel[4][2] ~^ image[18][18] + signed_kernel[4][3] ~^ image[18][19] + signed_kernel[4][4] ~^ image[18][20];
assign xor_sum[14][17] = signed_kernel[0][0] ~^ image[14][17] + signed_kernel[0][1] ~^ image[14][18] + signed_kernel[0][2] ~^ image[14][19] + signed_kernel[0][3] ~^ image[14][20] + signed_kernel[0][4] ~^ image[14][21] + signed_kernel[1][0] ~^ image[15][17] + signed_kernel[1][1] ~^ image[15][18] + signed_kernel[1][2] ~^ image[15][19] + signed_kernel[1][3] ~^ image[15][20] + signed_kernel[1][4] ~^ image[15][21] + signed_kernel[2][0] ~^ image[16][17] + signed_kernel[2][1] ~^ image[16][18] + signed_kernel[2][2] ~^ image[16][19] + signed_kernel[2][3] ~^ image[16][20] + signed_kernel[2][4] ~^ image[16][21] + signed_kernel[3][0] ~^ image[17][17] + signed_kernel[3][1] ~^ image[17][18] + signed_kernel[3][2] ~^ image[17][19] + signed_kernel[3][3] ~^ image[17][20] + signed_kernel[3][4] ~^ image[17][21] + signed_kernel[4][0] ~^ image[18][17] + signed_kernel[4][1] ~^ image[18][18] + signed_kernel[4][2] ~^ image[18][19] + signed_kernel[4][3] ~^ image[18][20] + signed_kernel[4][4] ~^ image[18][21];
assign xor_sum[14][18] = signed_kernel[0][0] ~^ image[14][18] + signed_kernel[0][1] ~^ image[14][19] + signed_kernel[0][2] ~^ image[14][20] + signed_kernel[0][3] ~^ image[14][21] + signed_kernel[0][4] ~^ image[14][22] + signed_kernel[1][0] ~^ image[15][18] + signed_kernel[1][1] ~^ image[15][19] + signed_kernel[1][2] ~^ image[15][20] + signed_kernel[1][3] ~^ image[15][21] + signed_kernel[1][4] ~^ image[15][22] + signed_kernel[2][0] ~^ image[16][18] + signed_kernel[2][1] ~^ image[16][19] + signed_kernel[2][2] ~^ image[16][20] + signed_kernel[2][3] ~^ image[16][21] + signed_kernel[2][4] ~^ image[16][22] + signed_kernel[3][0] ~^ image[17][18] + signed_kernel[3][1] ~^ image[17][19] + signed_kernel[3][2] ~^ image[17][20] + signed_kernel[3][3] ~^ image[17][21] + signed_kernel[3][4] ~^ image[17][22] + signed_kernel[4][0] ~^ image[18][18] + signed_kernel[4][1] ~^ image[18][19] + signed_kernel[4][2] ~^ image[18][20] + signed_kernel[4][3] ~^ image[18][21] + signed_kernel[4][4] ~^ image[18][22];
assign xor_sum[14][19] = signed_kernel[0][0] ~^ image[14][19] + signed_kernel[0][1] ~^ image[14][20] + signed_kernel[0][2] ~^ image[14][21] + signed_kernel[0][3] ~^ image[14][22] + signed_kernel[0][4] ~^ image[14][23] + signed_kernel[1][0] ~^ image[15][19] + signed_kernel[1][1] ~^ image[15][20] + signed_kernel[1][2] ~^ image[15][21] + signed_kernel[1][3] ~^ image[15][22] + signed_kernel[1][4] ~^ image[15][23] + signed_kernel[2][0] ~^ image[16][19] + signed_kernel[2][1] ~^ image[16][20] + signed_kernel[2][2] ~^ image[16][21] + signed_kernel[2][3] ~^ image[16][22] + signed_kernel[2][4] ~^ image[16][23] + signed_kernel[3][0] ~^ image[17][19] + signed_kernel[3][1] ~^ image[17][20] + signed_kernel[3][2] ~^ image[17][21] + signed_kernel[3][3] ~^ image[17][22] + signed_kernel[3][4] ~^ image[17][23] + signed_kernel[4][0] ~^ image[18][19] + signed_kernel[4][1] ~^ image[18][20] + signed_kernel[4][2] ~^ image[18][21] + signed_kernel[4][3] ~^ image[18][22] + signed_kernel[4][4] ~^ image[18][23];
assign xor_sum[14][20] = signed_kernel[0][0] ~^ image[14][20] + signed_kernel[0][1] ~^ image[14][21] + signed_kernel[0][2] ~^ image[14][22] + signed_kernel[0][3] ~^ image[14][23] + signed_kernel[0][4] ~^ image[14][24] + signed_kernel[1][0] ~^ image[15][20] + signed_kernel[1][1] ~^ image[15][21] + signed_kernel[1][2] ~^ image[15][22] + signed_kernel[1][3] ~^ image[15][23] + signed_kernel[1][4] ~^ image[15][24] + signed_kernel[2][0] ~^ image[16][20] + signed_kernel[2][1] ~^ image[16][21] + signed_kernel[2][2] ~^ image[16][22] + signed_kernel[2][3] ~^ image[16][23] + signed_kernel[2][4] ~^ image[16][24] + signed_kernel[3][0] ~^ image[17][20] + signed_kernel[3][1] ~^ image[17][21] + signed_kernel[3][2] ~^ image[17][22] + signed_kernel[3][3] ~^ image[17][23] + signed_kernel[3][4] ~^ image[17][24] + signed_kernel[4][0] ~^ image[18][20] + signed_kernel[4][1] ~^ image[18][21] + signed_kernel[4][2] ~^ image[18][22] + signed_kernel[4][3] ~^ image[18][23] + signed_kernel[4][4] ~^ image[18][24];
assign xor_sum[14][21] = signed_kernel[0][0] ~^ image[14][21] + signed_kernel[0][1] ~^ image[14][22] + signed_kernel[0][2] ~^ image[14][23] + signed_kernel[0][3] ~^ image[14][24] + signed_kernel[0][4] ~^ image[14][25] + signed_kernel[1][0] ~^ image[15][21] + signed_kernel[1][1] ~^ image[15][22] + signed_kernel[1][2] ~^ image[15][23] + signed_kernel[1][3] ~^ image[15][24] + signed_kernel[1][4] ~^ image[15][25] + signed_kernel[2][0] ~^ image[16][21] + signed_kernel[2][1] ~^ image[16][22] + signed_kernel[2][2] ~^ image[16][23] + signed_kernel[2][3] ~^ image[16][24] + signed_kernel[2][4] ~^ image[16][25] + signed_kernel[3][0] ~^ image[17][21] + signed_kernel[3][1] ~^ image[17][22] + signed_kernel[3][2] ~^ image[17][23] + signed_kernel[3][3] ~^ image[17][24] + signed_kernel[3][4] ~^ image[17][25] + signed_kernel[4][0] ~^ image[18][21] + signed_kernel[4][1] ~^ image[18][22] + signed_kernel[4][2] ~^ image[18][23] + signed_kernel[4][3] ~^ image[18][24] + signed_kernel[4][4] ~^ image[18][25];
assign xor_sum[14][22] = signed_kernel[0][0] ~^ image[14][22] + signed_kernel[0][1] ~^ image[14][23] + signed_kernel[0][2] ~^ image[14][24] + signed_kernel[0][3] ~^ image[14][25] + signed_kernel[0][4] ~^ image[14][26] + signed_kernel[1][0] ~^ image[15][22] + signed_kernel[1][1] ~^ image[15][23] + signed_kernel[1][2] ~^ image[15][24] + signed_kernel[1][3] ~^ image[15][25] + signed_kernel[1][4] ~^ image[15][26] + signed_kernel[2][0] ~^ image[16][22] + signed_kernel[2][1] ~^ image[16][23] + signed_kernel[2][2] ~^ image[16][24] + signed_kernel[2][3] ~^ image[16][25] + signed_kernel[2][4] ~^ image[16][26] + signed_kernel[3][0] ~^ image[17][22] + signed_kernel[3][1] ~^ image[17][23] + signed_kernel[3][2] ~^ image[17][24] + signed_kernel[3][3] ~^ image[17][25] + signed_kernel[3][4] ~^ image[17][26] + signed_kernel[4][0] ~^ image[18][22] + signed_kernel[4][1] ~^ image[18][23] + signed_kernel[4][2] ~^ image[18][24] + signed_kernel[4][3] ~^ image[18][25] + signed_kernel[4][4] ~^ image[18][26];
assign xor_sum[14][23] = signed_kernel[0][0] ~^ image[14][23] + signed_kernel[0][1] ~^ image[14][24] + signed_kernel[0][2] ~^ image[14][25] + signed_kernel[0][3] ~^ image[14][26] + signed_kernel[0][4] ~^ image[14][27] + signed_kernel[1][0] ~^ image[15][23] + signed_kernel[1][1] ~^ image[15][24] + signed_kernel[1][2] ~^ image[15][25] + signed_kernel[1][3] ~^ image[15][26] + signed_kernel[1][4] ~^ image[15][27] + signed_kernel[2][0] ~^ image[16][23] + signed_kernel[2][1] ~^ image[16][24] + signed_kernel[2][2] ~^ image[16][25] + signed_kernel[2][3] ~^ image[16][26] + signed_kernel[2][4] ~^ image[16][27] + signed_kernel[3][0] ~^ image[17][23] + signed_kernel[3][1] ~^ image[17][24] + signed_kernel[3][2] ~^ image[17][25] + signed_kernel[3][3] ~^ image[17][26] + signed_kernel[3][4] ~^ image[17][27] + signed_kernel[4][0] ~^ image[18][23] + signed_kernel[4][1] ~^ image[18][24] + signed_kernel[4][2] ~^ image[18][25] + signed_kernel[4][3] ~^ image[18][26] + signed_kernel[4][4] ~^ image[18][27];
assign xor_sum[15][0] = signed_kernel[0][0] ~^ image[15][0] + signed_kernel[0][1] ~^ image[15][1] + signed_kernel[0][2] ~^ image[15][2] + signed_kernel[0][3] ~^ image[15][3] + signed_kernel[0][4] ~^ image[15][4] + signed_kernel[1][0] ~^ image[16][0] + signed_kernel[1][1] ~^ image[16][1] + signed_kernel[1][2] ~^ image[16][2] + signed_kernel[1][3] ~^ image[16][3] + signed_kernel[1][4] ~^ image[16][4] + signed_kernel[2][0] ~^ image[17][0] + signed_kernel[2][1] ~^ image[17][1] + signed_kernel[2][2] ~^ image[17][2] + signed_kernel[2][3] ~^ image[17][3] + signed_kernel[2][4] ~^ image[17][4] + signed_kernel[3][0] ~^ image[18][0] + signed_kernel[3][1] ~^ image[18][1] + signed_kernel[3][2] ~^ image[18][2] + signed_kernel[3][3] ~^ image[18][3] + signed_kernel[3][4] ~^ image[18][4] + signed_kernel[4][0] ~^ image[19][0] + signed_kernel[4][1] ~^ image[19][1] + signed_kernel[4][2] ~^ image[19][2] + signed_kernel[4][3] ~^ image[19][3] + signed_kernel[4][4] ~^ image[19][4];
assign xor_sum[15][1] = signed_kernel[0][0] ~^ image[15][1] + signed_kernel[0][1] ~^ image[15][2] + signed_kernel[0][2] ~^ image[15][3] + signed_kernel[0][3] ~^ image[15][4] + signed_kernel[0][4] ~^ image[15][5] + signed_kernel[1][0] ~^ image[16][1] + signed_kernel[1][1] ~^ image[16][2] + signed_kernel[1][2] ~^ image[16][3] + signed_kernel[1][3] ~^ image[16][4] + signed_kernel[1][4] ~^ image[16][5] + signed_kernel[2][0] ~^ image[17][1] + signed_kernel[2][1] ~^ image[17][2] + signed_kernel[2][2] ~^ image[17][3] + signed_kernel[2][3] ~^ image[17][4] + signed_kernel[2][4] ~^ image[17][5] + signed_kernel[3][0] ~^ image[18][1] + signed_kernel[3][1] ~^ image[18][2] + signed_kernel[3][2] ~^ image[18][3] + signed_kernel[3][3] ~^ image[18][4] + signed_kernel[3][4] ~^ image[18][5] + signed_kernel[4][0] ~^ image[19][1] + signed_kernel[4][1] ~^ image[19][2] + signed_kernel[4][2] ~^ image[19][3] + signed_kernel[4][3] ~^ image[19][4] + signed_kernel[4][4] ~^ image[19][5];
assign xor_sum[15][2] = signed_kernel[0][0] ~^ image[15][2] + signed_kernel[0][1] ~^ image[15][3] + signed_kernel[0][2] ~^ image[15][4] + signed_kernel[0][3] ~^ image[15][5] + signed_kernel[0][4] ~^ image[15][6] + signed_kernel[1][0] ~^ image[16][2] + signed_kernel[1][1] ~^ image[16][3] + signed_kernel[1][2] ~^ image[16][4] + signed_kernel[1][3] ~^ image[16][5] + signed_kernel[1][4] ~^ image[16][6] + signed_kernel[2][0] ~^ image[17][2] + signed_kernel[2][1] ~^ image[17][3] + signed_kernel[2][2] ~^ image[17][4] + signed_kernel[2][3] ~^ image[17][5] + signed_kernel[2][4] ~^ image[17][6] + signed_kernel[3][0] ~^ image[18][2] + signed_kernel[3][1] ~^ image[18][3] + signed_kernel[3][2] ~^ image[18][4] + signed_kernel[3][3] ~^ image[18][5] + signed_kernel[3][4] ~^ image[18][6] + signed_kernel[4][0] ~^ image[19][2] + signed_kernel[4][1] ~^ image[19][3] + signed_kernel[4][2] ~^ image[19][4] + signed_kernel[4][3] ~^ image[19][5] + signed_kernel[4][4] ~^ image[19][6];
assign xor_sum[15][3] = signed_kernel[0][0] ~^ image[15][3] + signed_kernel[0][1] ~^ image[15][4] + signed_kernel[0][2] ~^ image[15][5] + signed_kernel[0][3] ~^ image[15][6] + signed_kernel[0][4] ~^ image[15][7] + signed_kernel[1][0] ~^ image[16][3] + signed_kernel[1][1] ~^ image[16][4] + signed_kernel[1][2] ~^ image[16][5] + signed_kernel[1][3] ~^ image[16][6] + signed_kernel[1][4] ~^ image[16][7] + signed_kernel[2][0] ~^ image[17][3] + signed_kernel[2][1] ~^ image[17][4] + signed_kernel[2][2] ~^ image[17][5] + signed_kernel[2][3] ~^ image[17][6] + signed_kernel[2][4] ~^ image[17][7] + signed_kernel[3][0] ~^ image[18][3] + signed_kernel[3][1] ~^ image[18][4] + signed_kernel[3][2] ~^ image[18][5] + signed_kernel[3][3] ~^ image[18][6] + signed_kernel[3][4] ~^ image[18][7] + signed_kernel[4][0] ~^ image[19][3] + signed_kernel[4][1] ~^ image[19][4] + signed_kernel[4][2] ~^ image[19][5] + signed_kernel[4][3] ~^ image[19][6] + signed_kernel[4][4] ~^ image[19][7];
assign xor_sum[15][4] = signed_kernel[0][0] ~^ image[15][4] + signed_kernel[0][1] ~^ image[15][5] + signed_kernel[0][2] ~^ image[15][6] + signed_kernel[0][3] ~^ image[15][7] + signed_kernel[0][4] ~^ image[15][8] + signed_kernel[1][0] ~^ image[16][4] + signed_kernel[1][1] ~^ image[16][5] + signed_kernel[1][2] ~^ image[16][6] + signed_kernel[1][3] ~^ image[16][7] + signed_kernel[1][4] ~^ image[16][8] + signed_kernel[2][0] ~^ image[17][4] + signed_kernel[2][1] ~^ image[17][5] + signed_kernel[2][2] ~^ image[17][6] + signed_kernel[2][3] ~^ image[17][7] + signed_kernel[2][4] ~^ image[17][8] + signed_kernel[3][0] ~^ image[18][4] + signed_kernel[3][1] ~^ image[18][5] + signed_kernel[3][2] ~^ image[18][6] + signed_kernel[3][3] ~^ image[18][7] + signed_kernel[3][4] ~^ image[18][8] + signed_kernel[4][0] ~^ image[19][4] + signed_kernel[4][1] ~^ image[19][5] + signed_kernel[4][2] ~^ image[19][6] + signed_kernel[4][3] ~^ image[19][7] + signed_kernel[4][4] ~^ image[19][8];
assign xor_sum[15][5] = signed_kernel[0][0] ~^ image[15][5] + signed_kernel[0][1] ~^ image[15][6] + signed_kernel[0][2] ~^ image[15][7] + signed_kernel[0][3] ~^ image[15][8] + signed_kernel[0][4] ~^ image[15][9] + signed_kernel[1][0] ~^ image[16][5] + signed_kernel[1][1] ~^ image[16][6] + signed_kernel[1][2] ~^ image[16][7] + signed_kernel[1][3] ~^ image[16][8] + signed_kernel[1][4] ~^ image[16][9] + signed_kernel[2][0] ~^ image[17][5] + signed_kernel[2][1] ~^ image[17][6] + signed_kernel[2][2] ~^ image[17][7] + signed_kernel[2][3] ~^ image[17][8] + signed_kernel[2][4] ~^ image[17][9] + signed_kernel[3][0] ~^ image[18][5] + signed_kernel[3][1] ~^ image[18][6] + signed_kernel[3][2] ~^ image[18][7] + signed_kernel[3][3] ~^ image[18][8] + signed_kernel[3][4] ~^ image[18][9] + signed_kernel[4][0] ~^ image[19][5] + signed_kernel[4][1] ~^ image[19][6] + signed_kernel[4][2] ~^ image[19][7] + signed_kernel[4][3] ~^ image[19][8] + signed_kernel[4][4] ~^ image[19][9];
assign xor_sum[15][6] = signed_kernel[0][0] ~^ image[15][6] + signed_kernel[0][1] ~^ image[15][7] + signed_kernel[0][2] ~^ image[15][8] + signed_kernel[0][3] ~^ image[15][9] + signed_kernel[0][4] ~^ image[15][10] + signed_kernel[1][0] ~^ image[16][6] + signed_kernel[1][1] ~^ image[16][7] + signed_kernel[1][2] ~^ image[16][8] + signed_kernel[1][3] ~^ image[16][9] + signed_kernel[1][4] ~^ image[16][10] + signed_kernel[2][0] ~^ image[17][6] + signed_kernel[2][1] ~^ image[17][7] + signed_kernel[2][2] ~^ image[17][8] + signed_kernel[2][3] ~^ image[17][9] + signed_kernel[2][4] ~^ image[17][10] + signed_kernel[3][0] ~^ image[18][6] + signed_kernel[3][1] ~^ image[18][7] + signed_kernel[3][2] ~^ image[18][8] + signed_kernel[3][3] ~^ image[18][9] + signed_kernel[3][4] ~^ image[18][10] + signed_kernel[4][0] ~^ image[19][6] + signed_kernel[4][1] ~^ image[19][7] + signed_kernel[4][2] ~^ image[19][8] + signed_kernel[4][3] ~^ image[19][9] + signed_kernel[4][4] ~^ image[19][10];
assign xor_sum[15][7] = signed_kernel[0][0] ~^ image[15][7] + signed_kernel[0][1] ~^ image[15][8] + signed_kernel[0][2] ~^ image[15][9] + signed_kernel[0][3] ~^ image[15][10] + signed_kernel[0][4] ~^ image[15][11] + signed_kernel[1][0] ~^ image[16][7] + signed_kernel[1][1] ~^ image[16][8] + signed_kernel[1][2] ~^ image[16][9] + signed_kernel[1][3] ~^ image[16][10] + signed_kernel[1][4] ~^ image[16][11] + signed_kernel[2][0] ~^ image[17][7] + signed_kernel[2][1] ~^ image[17][8] + signed_kernel[2][2] ~^ image[17][9] + signed_kernel[2][3] ~^ image[17][10] + signed_kernel[2][4] ~^ image[17][11] + signed_kernel[3][0] ~^ image[18][7] + signed_kernel[3][1] ~^ image[18][8] + signed_kernel[3][2] ~^ image[18][9] + signed_kernel[3][3] ~^ image[18][10] + signed_kernel[3][4] ~^ image[18][11] + signed_kernel[4][0] ~^ image[19][7] + signed_kernel[4][1] ~^ image[19][8] + signed_kernel[4][2] ~^ image[19][9] + signed_kernel[4][3] ~^ image[19][10] + signed_kernel[4][4] ~^ image[19][11];
assign xor_sum[15][8] = signed_kernel[0][0] ~^ image[15][8] + signed_kernel[0][1] ~^ image[15][9] + signed_kernel[0][2] ~^ image[15][10] + signed_kernel[0][3] ~^ image[15][11] + signed_kernel[0][4] ~^ image[15][12] + signed_kernel[1][0] ~^ image[16][8] + signed_kernel[1][1] ~^ image[16][9] + signed_kernel[1][2] ~^ image[16][10] + signed_kernel[1][3] ~^ image[16][11] + signed_kernel[1][4] ~^ image[16][12] + signed_kernel[2][0] ~^ image[17][8] + signed_kernel[2][1] ~^ image[17][9] + signed_kernel[2][2] ~^ image[17][10] + signed_kernel[2][3] ~^ image[17][11] + signed_kernel[2][4] ~^ image[17][12] + signed_kernel[3][0] ~^ image[18][8] + signed_kernel[3][1] ~^ image[18][9] + signed_kernel[3][2] ~^ image[18][10] + signed_kernel[3][3] ~^ image[18][11] + signed_kernel[3][4] ~^ image[18][12] + signed_kernel[4][0] ~^ image[19][8] + signed_kernel[4][1] ~^ image[19][9] + signed_kernel[4][2] ~^ image[19][10] + signed_kernel[4][3] ~^ image[19][11] + signed_kernel[4][4] ~^ image[19][12];
assign xor_sum[15][9] = signed_kernel[0][0] ~^ image[15][9] + signed_kernel[0][1] ~^ image[15][10] + signed_kernel[0][2] ~^ image[15][11] + signed_kernel[0][3] ~^ image[15][12] + signed_kernel[0][4] ~^ image[15][13] + signed_kernel[1][0] ~^ image[16][9] + signed_kernel[1][1] ~^ image[16][10] + signed_kernel[1][2] ~^ image[16][11] + signed_kernel[1][3] ~^ image[16][12] + signed_kernel[1][4] ~^ image[16][13] + signed_kernel[2][0] ~^ image[17][9] + signed_kernel[2][1] ~^ image[17][10] + signed_kernel[2][2] ~^ image[17][11] + signed_kernel[2][3] ~^ image[17][12] + signed_kernel[2][4] ~^ image[17][13] + signed_kernel[3][0] ~^ image[18][9] + signed_kernel[3][1] ~^ image[18][10] + signed_kernel[3][2] ~^ image[18][11] + signed_kernel[3][3] ~^ image[18][12] + signed_kernel[3][4] ~^ image[18][13] + signed_kernel[4][0] ~^ image[19][9] + signed_kernel[4][1] ~^ image[19][10] + signed_kernel[4][2] ~^ image[19][11] + signed_kernel[4][3] ~^ image[19][12] + signed_kernel[4][4] ~^ image[19][13];
assign xor_sum[15][10] = signed_kernel[0][0] ~^ image[15][10] + signed_kernel[0][1] ~^ image[15][11] + signed_kernel[0][2] ~^ image[15][12] + signed_kernel[0][3] ~^ image[15][13] + signed_kernel[0][4] ~^ image[15][14] + signed_kernel[1][0] ~^ image[16][10] + signed_kernel[1][1] ~^ image[16][11] + signed_kernel[1][2] ~^ image[16][12] + signed_kernel[1][3] ~^ image[16][13] + signed_kernel[1][4] ~^ image[16][14] + signed_kernel[2][0] ~^ image[17][10] + signed_kernel[2][1] ~^ image[17][11] + signed_kernel[2][2] ~^ image[17][12] + signed_kernel[2][3] ~^ image[17][13] + signed_kernel[2][4] ~^ image[17][14] + signed_kernel[3][0] ~^ image[18][10] + signed_kernel[3][1] ~^ image[18][11] + signed_kernel[3][2] ~^ image[18][12] + signed_kernel[3][3] ~^ image[18][13] + signed_kernel[3][4] ~^ image[18][14] + signed_kernel[4][0] ~^ image[19][10] + signed_kernel[4][1] ~^ image[19][11] + signed_kernel[4][2] ~^ image[19][12] + signed_kernel[4][3] ~^ image[19][13] + signed_kernel[4][4] ~^ image[19][14];
assign xor_sum[15][11] = signed_kernel[0][0] ~^ image[15][11] + signed_kernel[0][1] ~^ image[15][12] + signed_kernel[0][2] ~^ image[15][13] + signed_kernel[0][3] ~^ image[15][14] + signed_kernel[0][4] ~^ image[15][15] + signed_kernel[1][0] ~^ image[16][11] + signed_kernel[1][1] ~^ image[16][12] + signed_kernel[1][2] ~^ image[16][13] + signed_kernel[1][3] ~^ image[16][14] + signed_kernel[1][4] ~^ image[16][15] + signed_kernel[2][0] ~^ image[17][11] + signed_kernel[2][1] ~^ image[17][12] + signed_kernel[2][2] ~^ image[17][13] + signed_kernel[2][3] ~^ image[17][14] + signed_kernel[2][4] ~^ image[17][15] + signed_kernel[3][0] ~^ image[18][11] + signed_kernel[3][1] ~^ image[18][12] + signed_kernel[3][2] ~^ image[18][13] + signed_kernel[3][3] ~^ image[18][14] + signed_kernel[3][4] ~^ image[18][15] + signed_kernel[4][0] ~^ image[19][11] + signed_kernel[4][1] ~^ image[19][12] + signed_kernel[4][2] ~^ image[19][13] + signed_kernel[4][3] ~^ image[19][14] + signed_kernel[4][4] ~^ image[19][15];
assign xor_sum[15][12] = signed_kernel[0][0] ~^ image[15][12] + signed_kernel[0][1] ~^ image[15][13] + signed_kernel[0][2] ~^ image[15][14] + signed_kernel[0][3] ~^ image[15][15] + signed_kernel[0][4] ~^ image[15][16] + signed_kernel[1][0] ~^ image[16][12] + signed_kernel[1][1] ~^ image[16][13] + signed_kernel[1][2] ~^ image[16][14] + signed_kernel[1][3] ~^ image[16][15] + signed_kernel[1][4] ~^ image[16][16] + signed_kernel[2][0] ~^ image[17][12] + signed_kernel[2][1] ~^ image[17][13] + signed_kernel[2][2] ~^ image[17][14] + signed_kernel[2][3] ~^ image[17][15] + signed_kernel[2][4] ~^ image[17][16] + signed_kernel[3][0] ~^ image[18][12] + signed_kernel[3][1] ~^ image[18][13] + signed_kernel[3][2] ~^ image[18][14] + signed_kernel[3][3] ~^ image[18][15] + signed_kernel[3][4] ~^ image[18][16] + signed_kernel[4][0] ~^ image[19][12] + signed_kernel[4][1] ~^ image[19][13] + signed_kernel[4][2] ~^ image[19][14] + signed_kernel[4][3] ~^ image[19][15] + signed_kernel[4][4] ~^ image[19][16];
assign xor_sum[15][13] = signed_kernel[0][0] ~^ image[15][13] + signed_kernel[0][1] ~^ image[15][14] + signed_kernel[0][2] ~^ image[15][15] + signed_kernel[0][3] ~^ image[15][16] + signed_kernel[0][4] ~^ image[15][17] + signed_kernel[1][0] ~^ image[16][13] + signed_kernel[1][1] ~^ image[16][14] + signed_kernel[1][2] ~^ image[16][15] + signed_kernel[1][3] ~^ image[16][16] + signed_kernel[1][4] ~^ image[16][17] + signed_kernel[2][0] ~^ image[17][13] + signed_kernel[2][1] ~^ image[17][14] + signed_kernel[2][2] ~^ image[17][15] + signed_kernel[2][3] ~^ image[17][16] + signed_kernel[2][4] ~^ image[17][17] + signed_kernel[3][0] ~^ image[18][13] + signed_kernel[3][1] ~^ image[18][14] + signed_kernel[3][2] ~^ image[18][15] + signed_kernel[3][3] ~^ image[18][16] + signed_kernel[3][4] ~^ image[18][17] + signed_kernel[4][0] ~^ image[19][13] + signed_kernel[4][1] ~^ image[19][14] + signed_kernel[4][2] ~^ image[19][15] + signed_kernel[4][3] ~^ image[19][16] + signed_kernel[4][4] ~^ image[19][17];
assign xor_sum[15][14] = signed_kernel[0][0] ~^ image[15][14] + signed_kernel[0][1] ~^ image[15][15] + signed_kernel[0][2] ~^ image[15][16] + signed_kernel[0][3] ~^ image[15][17] + signed_kernel[0][4] ~^ image[15][18] + signed_kernel[1][0] ~^ image[16][14] + signed_kernel[1][1] ~^ image[16][15] + signed_kernel[1][2] ~^ image[16][16] + signed_kernel[1][3] ~^ image[16][17] + signed_kernel[1][4] ~^ image[16][18] + signed_kernel[2][0] ~^ image[17][14] + signed_kernel[2][1] ~^ image[17][15] + signed_kernel[2][2] ~^ image[17][16] + signed_kernel[2][3] ~^ image[17][17] + signed_kernel[2][4] ~^ image[17][18] + signed_kernel[3][0] ~^ image[18][14] + signed_kernel[3][1] ~^ image[18][15] + signed_kernel[3][2] ~^ image[18][16] + signed_kernel[3][3] ~^ image[18][17] + signed_kernel[3][4] ~^ image[18][18] + signed_kernel[4][0] ~^ image[19][14] + signed_kernel[4][1] ~^ image[19][15] + signed_kernel[4][2] ~^ image[19][16] + signed_kernel[4][3] ~^ image[19][17] + signed_kernel[4][4] ~^ image[19][18];
assign xor_sum[15][15] = signed_kernel[0][0] ~^ image[15][15] + signed_kernel[0][1] ~^ image[15][16] + signed_kernel[0][2] ~^ image[15][17] + signed_kernel[0][3] ~^ image[15][18] + signed_kernel[0][4] ~^ image[15][19] + signed_kernel[1][0] ~^ image[16][15] + signed_kernel[1][1] ~^ image[16][16] + signed_kernel[1][2] ~^ image[16][17] + signed_kernel[1][3] ~^ image[16][18] + signed_kernel[1][4] ~^ image[16][19] + signed_kernel[2][0] ~^ image[17][15] + signed_kernel[2][1] ~^ image[17][16] + signed_kernel[2][2] ~^ image[17][17] + signed_kernel[2][3] ~^ image[17][18] + signed_kernel[2][4] ~^ image[17][19] + signed_kernel[3][0] ~^ image[18][15] + signed_kernel[3][1] ~^ image[18][16] + signed_kernel[3][2] ~^ image[18][17] + signed_kernel[3][3] ~^ image[18][18] + signed_kernel[3][4] ~^ image[18][19] + signed_kernel[4][0] ~^ image[19][15] + signed_kernel[4][1] ~^ image[19][16] + signed_kernel[4][2] ~^ image[19][17] + signed_kernel[4][3] ~^ image[19][18] + signed_kernel[4][4] ~^ image[19][19];
assign xor_sum[15][16] = signed_kernel[0][0] ~^ image[15][16] + signed_kernel[0][1] ~^ image[15][17] + signed_kernel[0][2] ~^ image[15][18] + signed_kernel[0][3] ~^ image[15][19] + signed_kernel[0][4] ~^ image[15][20] + signed_kernel[1][0] ~^ image[16][16] + signed_kernel[1][1] ~^ image[16][17] + signed_kernel[1][2] ~^ image[16][18] + signed_kernel[1][3] ~^ image[16][19] + signed_kernel[1][4] ~^ image[16][20] + signed_kernel[2][0] ~^ image[17][16] + signed_kernel[2][1] ~^ image[17][17] + signed_kernel[2][2] ~^ image[17][18] + signed_kernel[2][3] ~^ image[17][19] + signed_kernel[2][4] ~^ image[17][20] + signed_kernel[3][0] ~^ image[18][16] + signed_kernel[3][1] ~^ image[18][17] + signed_kernel[3][2] ~^ image[18][18] + signed_kernel[3][3] ~^ image[18][19] + signed_kernel[3][4] ~^ image[18][20] + signed_kernel[4][0] ~^ image[19][16] + signed_kernel[4][1] ~^ image[19][17] + signed_kernel[4][2] ~^ image[19][18] + signed_kernel[4][3] ~^ image[19][19] + signed_kernel[4][4] ~^ image[19][20];
assign xor_sum[15][17] = signed_kernel[0][0] ~^ image[15][17] + signed_kernel[0][1] ~^ image[15][18] + signed_kernel[0][2] ~^ image[15][19] + signed_kernel[0][3] ~^ image[15][20] + signed_kernel[0][4] ~^ image[15][21] + signed_kernel[1][0] ~^ image[16][17] + signed_kernel[1][1] ~^ image[16][18] + signed_kernel[1][2] ~^ image[16][19] + signed_kernel[1][3] ~^ image[16][20] + signed_kernel[1][4] ~^ image[16][21] + signed_kernel[2][0] ~^ image[17][17] + signed_kernel[2][1] ~^ image[17][18] + signed_kernel[2][2] ~^ image[17][19] + signed_kernel[2][3] ~^ image[17][20] + signed_kernel[2][4] ~^ image[17][21] + signed_kernel[3][0] ~^ image[18][17] + signed_kernel[3][1] ~^ image[18][18] + signed_kernel[3][2] ~^ image[18][19] + signed_kernel[3][3] ~^ image[18][20] + signed_kernel[3][4] ~^ image[18][21] + signed_kernel[4][0] ~^ image[19][17] + signed_kernel[4][1] ~^ image[19][18] + signed_kernel[4][2] ~^ image[19][19] + signed_kernel[4][3] ~^ image[19][20] + signed_kernel[4][4] ~^ image[19][21];
assign xor_sum[15][18] = signed_kernel[0][0] ~^ image[15][18] + signed_kernel[0][1] ~^ image[15][19] + signed_kernel[0][2] ~^ image[15][20] + signed_kernel[0][3] ~^ image[15][21] + signed_kernel[0][4] ~^ image[15][22] + signed_kernel[1][0] ~^ image[16][18] + signed_kernel[1][1] ~^ image[16][19] + signed_kernel[1][2] ~^ image[16][20] + signed_kernel[1][3] ~^ image[16][21] + signed_kernel[1][4] ~^ image[16][22] + signed_kernel[2][0] ~^ image[17][18] + signed_kernel[2][1] ~^ image[17][19] + signed_kernel[2][2] ~^ image[17][20] + signed_kernel[2][3] ~^ image[17][21] + signed_kernel[2][4] ~^ image[17][22] + signed_kernel[3][0] ~^ image[18][18] + signed_kernel[3][1] ~^ image[18][19] + signed_kernel[3][2] ~^ image[18][20] + signed_kernel[3][3] ~^ image[18][21] + signed_kernel[3][4] ~^ image[18][22] + signed_kernel[4][0] ~^ image[19][18] + signed_kernel[4][1] ~^ image[19][19] + signed_kernel[4][2] ~^ image[19][20] + signed_kernel[4][3] ~^ image[19][21] + signed_kernel[4][4] ~^ image[19][22];
assign xor_sum[15][19] = signed_kernel[0][0] ~^ image[15][19] + signed_kernel[0][1] ~^ image[15][20] + signed_kernel[0][2] ~^ image[15][21] + signed_kernel[0][3] ~^ image[15][22] + signed_kernel[0][4] ~^ image[15][23] + signed_kernel[1][0] ~^ image[16][19] + signed_kernel[1][1] ~^ image[16][20] + signed_kernel[1][2] ~^ image[16][21] + signed_kernel[1][3] ~^ image[16][22] + signed_kernel[1][4] ~^ image[16][23] + signed_kernel[2][0] ~^ image[17][19] + signed_kernel[2][1] ~^ image[17][20] + signed_kernel[2][2] ~^ image[17][21] + signed_kernel[2][3] ~^ image[17][22] + signed_kernel[2][4] ~^ image[17][23] + signed_kernel[3][0] ~^ image[18][19] + signed_kernel[3][1] ~^ image[18][20] + signed_kernel[3][2] ~^ image[18][21] + signed_kernel[3][3] ~^ image[18][22] + signed_kernel[3][4] ~^ image[18][23] + signed_kernel[4][0] ~^ image[19][19] + signed_kernel[4][1] ~^ image[19][20] + signed_kernel[4][2] ~^ image[19][21] + signed_kernel[4][3] ~^ image[19][22] + signed_kernel[4][4] ~^ image[19][23];
assign xor_sum[15][20] = signed_kernel[0][0] ~^ image[15][20] + signed_kernel[0][1] ~^ image[15][21] + signed_kernel[0][2] ~^ image[15][22] + signed_kernel[0][3] ~^ image[15][23] + signed_kernel[0][4] ~^ image[15][24] + signed_kernel[1][0] ~^ image[16][20] + signed_kernel[1][1] ~^ image[16][21] + signed_kernel[1][2] ~^ image[16][22] + signed_kernel[1][3] ~^ image[16][23] + signed_kernel[1][4] ~^ image[16][24] + signed_kernel[2][0] ~^ image[17][20] + signed_kernel[2][1] ~^ image[17][21] + signed_kernel[2][2] ~^ image[17][22] + signed_kernel[2][3] ~^ image[17][23] + signed_kernel[2][4] ~^ image[17][24] + signed_kernel[3][0] ~^ image[18][20] + signed_kernel[3][1] ~^ image[18][21] + signed_kernel[3][2] ~^ image[18][22] + signed_kernel[3][3] ~^ image[18][23] + signed_kernel[3][4] ~^ image[18][24] + signed_kernel[4][0] ~^ image[19][20] + signed_kernel[4][1] ~^ image[19][21] + signed_kernel[4][2] ~^ image[19][22] + signed_kernel[4][3] ~^ image[19][23] + signed_kernel[4][4] ~^ image[19][24];
assign xor_sum[15][21] = signed_kernel[0][0] ~^ image[15][21] + signed_kernel[0][1] ~^ image[15][22] + signed_kernel[0][2] ~^ image[15][23] + signed_kernel[0][3] ~^ image[15][24] + signed_kernel[0][4] ~^ image[15][25] + signed_kernel[1][0] ~^ image[16][21] + signed_kernel[1][1] ~^ image[16][22] + signed_kernel[1][2] ~^ image[16][23] + signed_kernel[1][3] ~^ image[16][24] + signed_kernel[1][4] ~^ image[16][25] + signed_kernel[2][0] ~^ image[17][21] + signed_kernel[2][1] ~^ image[17][22] + signed_kernel[2][2] ~^ image[17][23] + signed_kernel[2][3] ~^ image[17][24] + signed_kernel[2][4] ~^ image[17][25] + signed_kernel[3][0] ~^ image[18][21] + signed_kernel[3][1] ~^ image[18][22] + signed_kernel[3][2] ~^ image[18][23] + signed_kernel[3][3] ~^ image[18][24] + signed_kernel[3][4] ~^ image[18][25] + signed_kernel[4][0] ~^ image[19][21] + signed_kernel[4][1] ~^ image[19][22] + signed_kernel[4][2] ~^ image[19][23] + signed_kernel[4][3] ~^ image[19][24] + signed_kernel[4][4] ~^ image[19][25];
assign xor_sum[15][22] = signed_kernel[0][0] ~^ image[15][22] + signed_kernel[0][1] ~^ image[15][23] + signed_kernel[0][2] ~^ image[15][24] + signed_kernel[0][3] ~^ image[15][25] + signed_kernel[0][4] ~^ image[15][26] + signed_kernel[1][0] ~^ image[16][22] + signed_kernel[1][1] ~^ image[16][23] + signed_kernel[1][2] ~^ image[16][24] + signed_kernel[1][3] ~^ image[16][25] + signed_kernel[1][4] ~^ image[16][26] + signed_kernel[2][0] ~^ image[17][22] + signed_kernel[2][1] ~^ image[17][23] + signed_kernel[2][2] ~^ image[17][24] + signed_kernel[2][3] ~^ image[17][25] + signed_kernel[2][4] ~^ image[17][26] + signed_kernel[3][0] ~^ image[18][22] + signed_kernel[3][1] ~^ image[18][23] + signed_kernel[3][2] ~^ image[18][24] + signed_kernel[3][3] ~^ image[18][25] + signed_kernel[3][4] ~^ image[18][26] + signed_kernel[4][0] ~^ image[19][22] + signed_kernel[4][1] ~^ image[19][23] + signed_kernel[4][2] ~^ image[19][24] + signed_kernel[4][3] ~^ image[19][25] + signed_kernel[4][4] ~^ image[19][26];
assign xor_sum[15][23] = signed_kernel[0][0] ~^ image[15][23] + signed_kernel[0][1] ~^ image[15][24] + signed_kernel[0][2] ~^ image[15][25] + signed_kernel[0][3] ~^ image[15][26] + signed_kernel[0][4] ~^ image[15][27] + signed_kernel[1][0] ~^ image[16][23] + signed_kernel[1][1] ~^ image[16][24] + signed_kernel[1][2] ~^ image[16][25] + signed_kernel[1][3] ~^ image[16][26] + signed_kernel[1][4] ~^ image[16][27] + signed_kernel[2][0] ~^ image[17][23] + signed_kernel[2][1] ~^ image[17][24] + signed_kernel[2][2] ~^ image[17][25] + signed_kernel[2][3] ~^ image[17][26] + signed_kernel[2][4] ~^ image[17][27] + signed_kernel[3][0] ~^ image[18][23] + signed_kernel[3][1] ~^ image[18][24] + signed_kernel[3][2] ~^ image[18][25] + signed_kernel[3][3] ~^ image[18][26] + signed_kernel[3][4] ~^ image[18][27] + signed_kernel[4][0] ~^ image[19][23] + signed_kernel[4][1] ~^ image[19][24] + signed_kernel[4][2] ~^ image[19][25] + signed_kernel[4][3] ~^ image[19][26] + signed_kernel[4][4] ~^ image[19][27];
assign xor_sum[16][0] = signed_kernel[0][0] ~^ image[16][0] + signed_kernel[0][1] ~^ image[16][1] + signed_kernel[0][2] ~^ image[16][2] + signed_kernel[0][3] ~^ image[16][3] + signed_kernel[0][4] ~^ image[16][4] + signed_kernel[1][0] ~^ image[17][0] + signed_kernel[1][1] ~^ image[17][1] + signed_kernel[1][2] ~^ image[17][2] + signed_kernel[1][3] ~^ image[17][3] + signed_kernel[1][4] ~^ image[17][4] + signed_kernel[2][0] ~^ image[18][0] + signed_kernel[2][1] ~^ image[18][1] + signed_kernel[2][2] ~^ image[18][2] + signed_kernel[2][3] ~^ image[18][3] + signed_kernel[2][4] ~^ image[18][4] + signed_kernel[3][0] ~^ image[19][0] + signed_kernel[3][1] ~^ image[19][1] + signed_kernel[3][2] ~^ image[19][2] + signed_kernel[3][3] ~^ image[19][3] + signed_kernel[3][4] ~^ image[19][4] + signed_kernel[4][0] ~^ image[20][0] + signed_kernel[4][1] ~^ image[20][1] + signed_kernel[4][2] ~^ image[20][2] + signed_kernel[4][3] ~^ image[20][3] + signed_kernel[4][4] ~^ image[20][4];
assign xor_sum[16][1] = signed_kernel[0][0] ~^ image[16][1] + signed_kernel[0][1] ~^ image[16][2] + signed_kernel[0][2] ~^ image[16][3] + signed_kernel[0][3] ~^ image[16][4] + signed_kernel[0][4] ~^ image[16][5] + signed_kernel[1][0] ~^ image[17][1] + signed_kernel[1][1] ~^ image[17][2] + signed_kernel[1][2] ~^ image[17][3] + signed_kernel[1][3] ~^ image[17][4] + signed_kernel[1][4] ~^ image[17][5] + signed_kernel[2][0] ~^ image[18][1] + signed_kernel[2][1] ~^ image[18][2] + signed_kernel[2][2] ~^ image[18][3] + signed_kernel[2][3] ~^ image[18][4] + signed_kernel[2][4] ~^ image[18][5] + signed_kernel[3][0] ~^ image[19][1] + signed_kernel[3][1] ~^ image[19][2] + signed_kernel[3][2] ~^ image[19][3] + signed_kernel[3][3] ~^ image[19][4] + signed_kernel[3][4] ~^ image[19][5] + signed_kernel[4][0] ~^ image[20][1] + signed_kernel[4][1] ~^ image[20][2] + signed_kernel[4][2] ~^ image[20][3] + signed_kernel[4][3] ~^ image[20][4] + signed_kernel[4][4] ~^ image[20][5];
assign xor_sum[16][2] = signed_kernel[0][0] ~^ image[16][2] + signed_kernel[0][1] ~^ image[16][3] + signed_kernel[0][2] ~^ image[16][4] + signed_kernel[0][3] ~^ image[16][5] + signed_kernel[0][4] ~^ image[16][6] + signed_kernel[1][0] ~^ image[17][2] + signed_kernel[1][1] ~^ image[17][3] + signed_kernel[1][2] ~^ image[17][4] + signed_kernel[1][3] ~^ image[17][5] + signed_kernel[1][4] ~^ image[17][6] + signed_kernel[2][0] ~^ image[18][2] + signed_kernel[2][1] ~^ image[18][3] + signed_kernel[2][2] ~^ image[18][4] + signed_kernel[2][3] ~^ image[18][5] + signed_kernel[2][4] ~^ image[18][6] + signed_kernel[3][0] ~^ image[19][2] + signed_kernel[3][1] ~^ image[19][3] + signed_kernel[3][2] ~^ image[19][4] + signed_kernel[3][3] ~^ image[19][5] + signed_kernel[3][4] ~^ image[19][6] + signed_kernel[4][0] ~^ image[20][2] + signed_kernel[4][1] ~^ image[20][3] + signed_kernel[4][2] ~^ image[20][4] + signed_kernel[4][3] ~^ image[20][5] + signed_kernel[4][4] ~^ image[20][6];
assign xor_sum[16][3] = signed_kernel[0][0] ~^ image[16][3] + signed_kernel[0][1] ~^ image[16][4] + signed_kernel[0][2] ~^ image[16][5] + signed_kernel[0][3] ~^ image[16][6] + signed_kernel[0][4] ~^ image[16][7] + signed_kernel[1][0] ~^ image[17][3] + signed_kernel[1][1] ~^ image[17][4] + signed_kernel[1][2] ~^ image[17][5] + signed_kernel[1][3] ~^ image[17][6] + signed_kernel[1][4] ~^ image[17][7] + signed_kernel[2][0] ~^ image[18][3] + signed_kernel[2][1] ~^ image[18][4] + signed_kernel[2][2] ~^ image[18][5] + signed_kernel[2][3] ~^ image[18][6] + signed_kernel[2][4] ~^ image[18][7] + signed_kernel[3][0] ~^ image[19][3] + signed_kernel[3][1] ~^ image[19][4] + signed_kernel[3][2] ~^ image[19][5] + signed_kernel[3][3] ~^ image[19][6] + signed_kernel[3][4] ~^ image[19][7] + signed_kernel[4][0] ~^ image[20][3] + signed_kernel[4][1] ~^ image[20][4] + signed_kernel[4][2] ~^ image[20][5] + signed_kernel[4][3] ~^ image[20][6] + signed_kernel[4][4] ~^ image[20][7];
assign xor_sum[16][4] = signed_kernel[0][0] ~^ image[16][4] + signed_kernel[0][1] ~^ image[16][5] + signed_kernel[0][2] ~^ image[16][6] + signed_kernel[0][3] ~^ image[16][7] + signed_kernel[0][4] ~^ image[16][8] + signed_kernel[1][0] ~^ image[17][4] + signed_kernel[1][1] ~^ image[17][5] + signed_kernel[1][2] ~^ image[17][6] + signed_kernel[1][3] ~^ image[17][7] + signed_kernel[1][4] ~^ image[17][8] + signed_kernel[2][0] ~^ image[18][4] + signed_kernel[2][1] ~^ image[18][5] + signed_kernel[2][2] ~^ image[18][6] + signed_kernel[2][3] ~^ image[18][7] + signed_kernel[2][4] ~^ image[18][8] + signed_kernel[3][0] ~^ image[19][4] + signed_kernel[3][1] ~^ image[19][5] + signed_kernel[3][2] ~^ image[19][6] + signed_kernel[3][3] ~^ image[19][7] + signed_kernel[3][4] ~^ image[19][8] + signed_kernel[4][0] ~^ image[20][4] + signed_kernel[4][1] ~^ image[20][5] + signed_kernel[4][2] ~^ image[20][6] + signed_kernel[4][3] ~^ image[20][7] + signed_kernel[4][4] ~^ image[20][8];
assign xor_sum[16][5] = signed_kernel[0][0] ~^ image[16][5] + signed_kernel[0][1] ~^ image[16][6] + signed_kernel[0][2] ~^ image[16][7] + signed_kernel[0][3] ~^ image[16][8] + signed_kernel[0][4] ~^ image[16][9] + signed_kernel[1][0] ~^ image[17][5] + signed_kernel[1][1] ~^ image[17][6] + signed_kernel[1][2] ~^ image[17][7] + signed_kernel[1][3] ~^ image[17][8] + signed_kernel[1][4] ~^ image[17][9] + signed_kernel[2][0] ~^ image[18][5] + signed_kernel[2][1] ~^ image[18][6] + signed_kernel[2][2] ~^ image[18][7] + signed_kernel[2][3] ~^ image[18][8] + signed_kernel[2][4] ~^ image[18][9] + signed_kernel[3][0] ~^ image[19][5] + signed_kernel[3][1] ~^ image[19][6] + signed_kernel[3][2] ~^ image[19][7] + signed_kernel[3][3] ~^ image[19][8] + signed_kernel[3][4] ~^ image[19][9] + signed_kernel[4][0] ~^ image[20][5] + signed_kernel[4][1] ~^ image[20][6] + signed_kernel[4][2] ~^ image[20][7] + signed_kernel[4][3] ~^ image[20][8] + signed_kernel[4][4] ~^ image[20][9];
assign xor_sum[16][6] = signed_kernel[0][0] ~^ image[16][6] + signed_kernel[0][1] ~^ image[16][7] + signed_kernel[0][2] ~^ image[16][8] + signed_kernel[0][3] ~^ image[16][9] + signed_kernel[0][4] ~^ image[16][10] + signed_kernel[1][0] ~^ image[17][6] + signed_kernel[1][1] ~^ image[17][7] + signed_kernel[1][2] ~^ image[17][8] + signed_kernel[1][3] ~^ image[17][9] + signed_kernel[1][4] ~^ image[17][10] + signed_kernel[2][0] ~^ image[18][6] + signed_kernel[2][1] ~^ image[18][7] + signed_kernel[2][2] ~^ image[18][8] + signed_kernel[2][3] ~^ image[18][9] + signed_kernel[2][4] ~^ image[18][10] + signed_kernel[3][0] ~^ image[19][6] + signed_kernel[3][1] ~^ image[19][7] + signed_kernel[3][2] ~^ image[19][8] + signed_kernel[3][3] ~^ image[19][9] + signed_kernel[3][4] ~^ image[19][10] + signed_kernel[4][0] ~^ image[20][6] + signed_kernel[4][1] ~^ image[20][7] + signed_kernel[4][2] ~^ image[20][8] + signed_kernel[4][3] ~^ image[20][9] + signed_kernel[4][4] ~^ image[20][10];
assign xor_sum[16][7] = signed_kernel[0][0] ~^ image[16][7] + signed_kernel[0][1] ~^ image[16][8] + signed_kernel[0][2] ~^ image[16][9] + signed_kernel[0][3] ~^ image[16][10] + signed_kernel[0][4] ~^ image[16][11] + signed_kernel[1][0] ~^ image[17][7] + signed_kernel[1][1] ~^ image[17][8] + signed_kernel[1][2] ~^ image[17][9] + signed_kernel[1][3] ~^ image[17][10] + signed_kernel[1][4] ~^ image[17][11] + signed_kernel[2][0] ~^ image[18][7] + signed_kernel[2][1] ~^ image[18][8] + signed_kernel[2][2] ~^ image[18][9] + signed_kernel[2][3] ~^ image[18][10] + signed_kernel[2][4] ~^ image[18][11] + signed_kernel[3][0] ~^ image[19][7] + signed_kernel[3][1] ~^ image[19][8] + signed_kernel[3][2] ~^ image[19][9] + signed_kernel[3][3] ~^ image[19][10] + signed_kernel[3][4] ~^ image[19][11] + signed_kernel[4][0] ~^ image[20][7] + signed_kernel[4][1] ~^ image[20][8] + signed_kernel[4][2] ~^ image[20][9] + signed_kernel[4][3] ~^ image[20][10] + signed_kernel[4][4] ~^ image[20][11];
assign xor_sum[16][8] = signed_kernel[0][0] ~^ image[16][8] + signed_kernel[0][1] ~^ image[16][9] + signed_kernel[0][2] ~^ image[16][10] + signed_kernel[0][3] ~^ image[16][11] + signed_kernel[0][4] ~^ image[16][12] + signed_kernel[1][0] ~^ image[17][8] + signed_kernel[1][1] ~^ image[17][9] + signed_kernel[1][2] ~^ image[17][10] + signed_kernel[1][3] ~^ image[17][11] + signed_kernel[1][4] ~^ image[17][12] + signed_kernel[2][0] ~^ image[18][8] + signed_kernel[2][1] ~^ image[18][9] + signed_kernel[2][2] ~^ image[18][10] + signed_kernel[2][3] ~^ image[18][11] + signed_kernel[2][4] ~^ image[18][12] + signed_kernel[3][0] ~^ image[19][8] + signed_kernel[3][1] ~^ image[19][9] + signed_kernel[3][2] ~^ image[19][10] + signed_kernel[3][3] ~^ image[19][11] + signed_kernel[3][4] ~^ image[19][12] + signed_kernel[4][0] ~^ image[20][8] + signed_kernel[4][1] ~^ image[20][9] + signed_kernel[4][2] ~^ image[20][10] + signed_kernel[4][3] ~^ image[20][11] + signed_kernel[4][4] ~^ image[20][12];
assign xor_sum[16][9] = signed_kernel[0][0] ~^ image[16][9] + signed_kernel[0][1] ~^ image[16][10] + signed_kernel[0][2] ~^ image[16][11] + signed_kernel[0][3] ~^ image[16][12] + signed_kernel[0][4] ~^ image[16][13] + signed_kernel[1][0] ~^ image[17][9] + signed_kernel[1][1] ~^ image[17][10] + signed_kernel[1][2] ~^ image[17][11] + signed_kernel[1][3] ~^ image[17][12] + signed_kernel[1][4] ~^ image[17][13] + signed_kernel[2][0] ~^ image[18][9] + signed_kernel[2][1] ~^ image[18][10] + signed_kernel[2][2] ~^ image[18][11] + signed_kernel[2][3] ~^ image[18][12] + signed_kernel[2][4] ~^ image[18][13] + signed_kernel[3][0] ~^ image[19][9] + signed_kernel[3][1] ~^ image[19][10] + signed_kernel[3][2] ~^ image[19][11] + signed_kernel[3][3] ~^ image[19][12] + signed_kernel[3][4] ~^ image[19][13] + signed_kernel[4][0] ~^ image[20][9] + signed_kernel[4][1] ~^ image[20][10] + signed_kernel[4][2] ~^ image[20][11] + signed_kernel[4][3] ~^ image[20][12] + signed_kernel[4][4] ~^ image[20][13];
assign xor_sum[16][10] = signed_kernel[0][0] ~^ image[16][10] + signed_kernel[0][1] ~^ image[16][11] + signed_kernel[0][2] ~^ image[16][12] + signed_kernel[0][3] ~^ image[16][13] + signed_kernel[0][4] ~^ image[16][14] + signed_kernel[1][0] ~^ image[17][10] + signed_kernel[1][1] ~^ image[17][11] + signed_kernel[1][2] ~^ image[17][12] + signed_kernel[1][3] ~^ image[17][13] + signed_kernel[1][4] ~^ image[17][14] + signed_kernel[2][0] ~^ image[18][10] + signed_kernel[2][1] ~^ image[18][11] + signed_kernel[2][2] ~^ image[18][12] + signed_kernel[2][3] ~^ image[18][13] + signed_kernel[2][4] ~^ image[18][14] + signed_kernel[3][0] ~^ image[19][10] + signed_kernel[3][1] ~^ image[19][11] + signed_kernel[3][2] ~^ image[19][12] + signed_kernel[3][3] ~^ image[19][13] + signed_kernel[3][4] ~^ image[19][14] + signed_kernel[4][0] ~^ image[20][10] + signed_kernel[4][1] ~^ image[20][11] + signed_kernel[4][2] ~^ image[20][12] + signed_kernel[4][3] ~^ image[20][13] + signed_kernel[4][4] ~^ image[20][14];
assign xor_sum[16][11] = signed_kernel[0][0] ~^ image[16][11] + signed_kernel[0][1] ~^ image[16][12] + signed_kernel[0][2] ~^ image[16][13] + signed_kernel[0][3] ~^ image[16][14] + signed_kernel[0][4] ~^ image[16][15] + signed_kernel[1][0] ~^ image[17][11] + signed_kernel[1][1] ~^ image[17][12] + signed_kernel[1][2] ~^ image[17][13] + signed_kernel[1][3] ~^ image[17][14] + signed_kernel[1][4] ~^ image[17][15] + signed_kernel[2][0] ~^ image[18][11] + signed_kernel[2][1] ~^ image[18][12] + signed_kernel[2][2] ~^ image[18][13] + signed_kernel[2][3] ~^ image[18][14] + signed_kernel[2][4] ~^ image[18][15] + signed_kernel[3][0] ~^ image[19][11] + signed_kernel[3][1] ~^ image[19][12] + signed_kernel[3][2] ~^ image[19][13] + signed_kernel[3][3] ~^ image[19][14] + signed_kernel[3][4] ~^ image[19][15] + signed_kernel[4][0] ~^ image[20][11] + signed_kernel[4][1] ~^ image[20][12] + signed_kernel[4][2] ~^ image[20][13] + signed_kernel[4][3] ~^ image[20][14] + signed_kernel[4][4] ~^ image[20][15];
assign xor_sum[16][12] = signed_kernel[0][0] ~^ image[16][12] + signed_kernel[0][1] ~^ image[16][13] + signed_kernel[0][2] ~^ image[16][14] + signed_kernel[0][3] ~^ image[16][15] + signed_kernel[0][4] ~^ image[16][16] + signed_kernel[1][0] ~^ image[17][12] + signed_kernel[1][1] ~^ image[17][13] + signed_kernel[1][2] ~^ image[17][14] + signed_kernel[1][3] ~^ image[17][15] + signed_kernel[1][4] ~^ image[17][16] + signed_kernel[2][0] ~^ image[18][12] + signed_kernel[2][1] ~^ image[18][13] + signed_kernel[2][2] ~^ image[18][14] + signed_kernel[2][3] ~^ image[18][15] + signed_kernel[2][4] ~^ image[18][16] + signed_kernel[3][0] ~^ image[19][12] + signed_kernel[3][1] ~^ image[19][13] + signed_kernel[3][2] ~^ image[19][14] + signed_kernel[3][3] ~^ image[19][15] + signed_kernel[3][4] ~^ image[19][16] + signed_kernel[4][0] ~^ image[20][12] + signed_kernel[4][1] ~^ image[20][13] + signed_kernel[4][2] ~^ image[20][14] + signed_kernel[4][3] ~^ image[20][15] + signed_kernel[4][4] ~^ image[20][16];
assign xor_sum[16][13] = signed_kernel[0][0] ~^ image[16][13] + signed_kernel[0][1] ~^ image[16][14] + signed_kernel[0][2] ~^ image[16][15] + signed_kernel[0][3] ~^ image[16][16] + signed_kernel[0][4] ~^ image[16][17] + signed_kernel[1][0] ~^ image[17][13] + signed_kernel[1][1] ~^ image[17][14] + signed_kernel[1][2] ~^ image[17][15] + signed_kernel[1][3] ~^ image[17][16] + signed_kernel[1][4] ~^ image[17][17] + signed_kernel[2][0] ~^ image[18][13] + signed_kernel[2][1] ~^ image[18][14] + signed_kernel[2][2] ~^ image[18][15] + signed_kernel[2][3] ~^ image[18][16] + signed_kernel[2][4] ~^ image[18][17] + signed_kernel[3][0] ~^ image[19][13] + signed_kernel[3][1] ~^ image[19][14] + signed_kernel[3][2] ~^ image[19][15] + signed_kernel[3][3] ~^ image[19][16] + signed_kernel[3][4] ~^ image[19][17] + signed_kernel[4][0] ~^ image[20][13] + signed_kernel[4][1] ~^ image[20][14] + signed_kernel[4][2] ~^ image[20][15] + signed_kernel[4][3] ~^ image[20][16] + signed_kernel[4][4] ~^ image[20][17];
assign xor_sum[16][14] = signed_kernel[0][0] ~^ image[16][14] + signed_kernel[0][1] ~^ image[16][15] + signed_kernel[0][2] ~^ image[16][16] + signed_kernel[0][3] ~^ image[16][17] + signed_kernel[0][4] ~^ image[16][18] + signed_kernel[1][0] ~^ image[17][14] + signed_kernel[1][1] ~^ image[17][15] + signed_kernel[1][2] ~^ image[17][16] + signed_kernel[1][3] ~^ image[17][17] + signed_kernel[1][4] ~^ image[17][18] + signed_kernel[2][0] ~^ image[18][14] + signed_kernel[2][1] ~^ image[18][15] + signed_kernel[2][2] ~^ image[18][16] + signed_kernel[2][3] ~^ image[18][17] + signed_kernel[2][4] ~^ image[18][18] + signed_kernel[3][0] ~^ image[19][14] + signed_kernel[3][1] ~^ image[19][15] + signed_kernel[3][2] ~^ image[19][16] + signed_kernel[3][3] ~^ image[19][17] + signed_kernel[3][4] ~^ image[19][18] + signed_kernel[4][0] ~^ image[20][14] + signed_kernel[4][1] ~^ image[20][15] + signed_kernel[4][2] ~^ image[20][16] + signed_kernel[4][3] ~^ image[20][17] + signed_kernel[4][4] ~^ image[20][18];
assign xor_sum[16][15] = signed_kernel[0][0] ~^ image[16][15] + signed_kernel[0][1] ~^ image[16][16] + signed_kernel[0][2] ~^ image[16][17] + signed_kernel[0][3] ~^ image[16][18] + signed_kernel[0][4] ~^ image[16][19] + signed_kernel[1][0] ~^ image[17][15] + signed_kernel[1][1] ~^ image[17][16] + signed_kernel[1][2] ~^ image[17][17] + signed_kernel[1][3] ~^ image[17][18] + signed_kernel[1][4] ~^ image[17][19] + signed_kernel[2][0] ~^ image[18][15] + signed_kernel[2][1] ~^ image[18][16] + signed_kernel[2][2] ~^ image[18][17] + signed_kernel[2][3] ~^ image[18][18] + signed_kernel[2][4] ~^ image[18][19] + signed_kernel[3][0] ~^ image[19][15] + signed_kernel[3][1] ~^ image[19][16] + signed_kernel[3][2] ~^ image[19][17] + signed_kernel[3][3] ~^ image[19][18] + signed_kernel[3][4] ~^ image[19][19] + signed_kernel[4][0] ~^ image[20][15] + signed_kernel[4][1] ~^ image[20][16] + signed_kernel[4][2] ~^ image[20][17] + signed_kernel[4][3] ~^ image[20][18] + signed_kernel[4][4] ~^ image[20][19];
assign xor_sum[16][16] = signed_kernel[0][0] ~^ image[16][16] + signed_kernel[0][1] ~^ image[16][17] + signed_kernel[0][2] ~^ image[16][18] + signed_kernel[0][3] ~^ image[16][19] + signed_kernel[0][4] ~^ image[16][20] + signed_kernel[1][0] ~^ image[17][16] + signed_kernel[1][1] ~^ image[17][17] + signed_kernel[1][2] ~^ image[17][18] + signed_kernel[1][3] ~^ image[17][19] + signed_kernel[1][4] ~^ image[17][20] + signed_kernel[2][0] ~^ image[18][16] + signed_kernel[2][1] ~^ image[18][17] + signed_kernel[2][2] ~^ image[18][18] + signed_kernel[2][3] ~^ image[18][19] + signed_kernel[2][4] ~^ image[18][20] + signed_kernel[3][0] ~^ image[19][16] + signed_kernel[3][1] ~^ image[19][17] + signed_kernel[3][2] ~^ image[19][18] + signed_kernel[3][3] ~^ image[19][19] + signed_kernel[3][4] ~^ image[19][20] + signed_kernel[4][0] ~^ image[20][16] + signed_kernel[4][1] ~^ image[20][17] + signed_kernel[4][2] ~^ image[20][18] + signed_kernel[4][3] ~^ image[20][19] + signed_kernel[4][4] ~^ image[20][20];
assign xor_sum[16][17] = signed_kernel[0][0] ~^ image[16][17] + signed_kernel[0][1] ~^ image[16][18] + signed_kernel[0][2] ~^ image[16][19] + signed_kernel[0][3] ~^ image[16][20] + signed_kernel[0][4] ~^ image[16][21] + signed_kernel[1][0] ~^ image[17][17] + signed_kernel[1][1] ~^ image[17][18] + signed_kernel[1][2] ~^ image[17][19] + signed_kernel[1][3] ~^ image[17][20] + signed_kernel[1][4] ~^ image[17][21] + signed_kernel[2][0] ~^ image[18][17] + signed_kernel[2][1] ~^ image[18][18] + signed_kernel[2][2] ~^ image[18][19] + signed_kernel[2][3] ~^ image[18][20] + signed_kernel[2][4] ~^ image[18][21] + signed_kernel[3][0] ~^ image[19][17] + signed_kernel[3][1] ~^ image[19][18] + signed_kernel[3][2] ~^ image[19][19] + signed_kernel[3][3] ~^ image[19][20] + signed_kernel[3][4] ~^ image[19][21] + signed_kernel[4][0] ~^ image[20][17] + signed_kernel[4][1] ~^ image[20][18] + signed_kernel[4][2] ~^ image[20][19] + signed_kernel[4][3] ~^ image[20][20] + signed_kernel[4][4] ~^ image[20][21];
assign xor_sum[16][18] = signed_kernel[0][0] ~^ image[16][18] + signed_kernel[0][1] ~^ image[16][19] + signed_kernel[0][2] ~^ image[16][20] + signed_kernel[0][3] ~^ image[16][21] + signed_kernel[0][4] ~^ image[16][22] + signed_kernel[1][0] ~^ image[17][18] + signed_kernel[1][1] ~^ image[17][19] + signed_kernel[1][2] ~^ image[17][20] + signed_kernel[1][3] ~^ image[17][21] + signed_kernel[1][4] ~^ image[17][22] + signed_kernel[2][0] ~^ image[18][18] + signed_kernel[2][1] ~^ image[18][19] + signed_kernel[2][2] ~^ image[18][20] + signed_kernel[2][3] ~^ image[18][21] + signed_kernel[2][4] ~^ image[18][22] + signed_kernel[3][0] ~^ image[19][18] + signed_kernel[3][1] ~^ image[19][19] + signed_kernel[3][2] ~^ image[19][20] + signed_kernel[3][3] ~^ image[19][21] + signed_kernel[3][4] ~^ image[19][22] + signed_kernel[4][0] ~^ image[20][18] + signed_kernel[4][1] ~^ image[20][19] + signed_kernel[4][2] ~^ image[20][20] + signed_kernel[4][3] ~^ image[20][21] + signed_kernel[4][4] ~^ image[20][22];
assign xor_sum[16][19] = signed_kernel[0][0] ~^ image[16][19] + signed_kernel[0][1] ~^ image[16][20] + signed_kernel[0][2] ~^ image[16][21] + signed_kernel[0][3] ~^ image[16][22] + signed_kernel[0][4] ~^ image[16][23] + signed_kernel[1][0] ~^ image[17][19] + signed_kernel[1][1] ~^ image[17][20] + signed_kernel[1][2] ~^ image[17][21] + signed_kernel[1][3] ~^ image[17][22] + signed_kernel[1][4] ~^ image[17][23] + signed_kernel[2][0] ~^ image[18][19] + signed_kernel[2][1] ~^ image[18][20] + signed_kernel[2][2] ~^ image[18][21] + signed_kernel[2][3] ~^ image[18][22] + signed_kernel[2][4] ~^ image[18][23] + signed_kernel[3][0] ~^ image[19][19] + signed_kernel[3][1] ~^ image[19][20] + signed_kernel[3][2] ~^ image[19][21] + signed_kernel[3][3] ~^ image[19][22] + signed_kernel[3][4] ~^ image[19][23] + signed_kernel[4][0] ~^ image[20][19] + signed_kernel[4][1] ~^ image[20][20] + signed_kernel[4][2] ~^ image[20][21] + signed_kernel[4][3] ~^ image[20][22] + signed_kernel[4][4] ~^ image[20][23];
assign xor_sum[16][20] = signed_kernel[0][0] ~^ image[16][20] + signed_kernel[0][1] ~^ image[16][21] + signed_kernel[0][2] ~^ image[16][22] + signed_kernel[0][3] ~^ image[16][23] + signed_kernel[0][4] ~^ image[16][24] + signed_kernel[1][0] ~^ image[17][20] + signed_kernel[1][1] ~^ image[17][21] + signed_kernel[1][2] ~^ image[17][22] + signed_kernel[1][3] ~^ image[17][23] + signed_kernel[1][4] ~^ image[17][24] + signed_kernel[2][0] ~^ image[18][20] + signed_kernel[2][1] ~^ image[18][21] + signed_kernel[2][2] ~^ image[18][22] + signed_kernel[2][3] ~^ image[18][23] + signed_kernel[2][4] ~^ image[18][24] + signed_kernel[3][0] ~^ image[19][20] + signed_kernel[3][1] ~^ image[19][21] + signed_kernel[3][2] ~^ image[19][22] + signed_kernel[3][3] ~^ image[19][23] + signed_kernel[3][4] ~^ image[19][24] + signed_kernel[4][0] ~^ image[20][20] + signed_kernel[4][1] ~^ image[20][21] + signed_kernel[4][2] ~^ image[20][22] + signed_kernel[4][3] ~^ image[20][23] + signed_kernel[4][4] ~^ image[20][24];
assign xor_sum[16][21] = signed_kernel[0][0] ~^ image[16][21] + signed_kernel[0][1] ~^ image[16][22] + signed_kernel[0][2] ~^ image[16][23] + signed_kernel[0][3] ~^ image[16][24] + signed_kernel[0][4] ~^ image[16][25] + signed_kernel[1][0] ~^ image[17][21] + signed_kernel[1][1] ~^ image[17][22] + signed_kernel[1][2] ~^ image[17][23] + signed_kernel[1][3] ~^ image[17][24] + signed_kernel[1][4] ~^ image[17][25] + signed_kernel[2][0] ~^ image[18][21] + signed_kernel[2][1] ~^ image[18][22] + signed_kernel[2][2] ~^ image[18][23] + signed_kernel[2][3] ~^ image[18][24] + signed_kernel[2][4] ~^ image[18][25] + signed_kernel[3][0] ~^ image[19][21] + signed_kernel[3][1] ~^ image[19][22] + signed_kernel[3][2] ~^ image[19][23] + signed_kernel[3][3] ~^ image[19][24] + signed_kernel[3][4] ~^ image[19][25] + signed_kernel[4][0] ~^ image[20][21] + signed_kernel[4][1] ~^ image[20][22] + signed_kernel[4][2] ~^ image[20][23] + signed_kernel[4][3] ~^ image[20][24] + signed_kernel[4][4] ~^ image[20][25];
assign xor_sum[16][22] = signed_kernel[0][0] ~^ image[16][22] + signed_kernel[0][1] ~^ image[16][23] + signed_kernel[0][2] ~^ image[16][24] + signed_kernel[0][3] ~^ image[16][25] + signed_kernel[0][4] ~^ image[16][26] + signed_kernel[1][0] ~^ image[17][22] + signed_kernel[1][1] ~^ image[17][23] + signed_kernel[1][2] ~^ image[17][24] + signed_kernel[1][3] ~^ image[17][25] + signed_kernel[1][4] ~^ image[17][26] + signed_kernel[2][0] ~^ image[18][22] + signed_kernel[2][1] ~^ image[18][23] + signed_kernel[2][2] ~^ image[18][24] + signed_kernel[2][3] ~^ image[18][25] + signed_kernel[2][4] ~^ image[18][26] + signed_kernel[3][0] ~^ image[19][22] + signed_kernel[3][1] ~^ image[19][23] + signed_kernel[3][2] ~^ image[19][24] + signed_kernel[3][3] ~^ image[19][25] + signed_kernel[3][4] ~^ image[19][26] + signed_kernel[4][0] ~^ image[20][22] + signed_kernel[4][1] ~^ image[20][23] + signed_kernel[4][2] ~^ image[20][24] + signed_kernel[4][3] ~^ image[20][25] + signed_kernel[4][4] ~^ image[20][26];
assign xor_sum[16][23] = signed_kernel[0][0] ~^ image[16][23] + signed_kernel[0][1] ~^ image[16][24] + signed_kernel[0][2] ~^ image[16][25] + signed_kernel[0][3] ~^ image[16][26] + signed_kernel[0][4] ~^ image[16][27] + signed_kernel[1][0] ~^ image[17][23] + signed_kernel[1][1] ~^ image[17][24] + signed_kernel[1][2] ~^ image[17][25] + signed_kernel[1][3] ~^ image[17][26] + signed_kernel[1][4] ~^ image[17][27] + signed_kernel[2][0] ~^ image[18][23] + signed_kernel[2][1] ~^ image[18][24] + signed_kernel[2][2] ~^ image[18][25] + signed_kernel[2][3] ~^ image[18][26] + signed_kernel[2][4] ~^ image[18][27] + signed_kernel[3][0] ~^ image[19][23] + signed_kernel[3][1] ~^ image[19][24] + signed_kernel[3][2] ~^ image[19][25] + signed_kernel[3][3] ~^ image[19][26] + signed_kernel[3][4] ~^ image[19][27] + signed_kernel[4][0] ~^ image[20][23] + signed_kernel[4][1] ~^ image[20][24] + signed_kernel[4][2] ~^ image[20][25] + signed_kernel[4][3] ~^ image[20][26] + signed_kernel[4][4] ~^ image[20][27];
assign xor_sum[17][0] = signed_kernel[0][0] ~^ image[17][0] + signed_kernel[0][1] ~^ image[17][1] + signed_kernel[0][2] ~^ image[17][2] + signed_kernel[0][3] ~^ image[17][3] + signed_kernel[0][4] ~^ image[17][4] + signed_kernel[1][0] ~^ image[18][0] + signed_kernel[1][1] ~^ image[18][1] + signed_kernel[1][2] ~^ image[18][2] + signed_kernel[1][3] ~^ image[18][3] + signed_kernel[1][4] ~^ image[18][4] + signed_kernel[2][0] ~^ image[19][0] + signed_kernel[2][1] ~^ image[19][1] + signed_kernel[2][2] ~^ image[19][2] + signed_kernel[2][3] ~^ image[19][3] + signed_kernel[2][4] ~^ image[19][4] + signed_kernel[3][0] ~^ image[20][0] + signed_kernel[3][1] ~^ image[20][1] + signed_kernel[3][2] ~^ image[20][2] + signed_kernel[3][3] ~^ image[20][3] + signed_kernel[3][4] ~^ image[20][4] + signed_kernel[4][0] ~^ image[21][0] + signed_kernel[4][1] ~^ image[21][1] + signed_kernel[4][2] ~^ image[21][2] + signed_kernel[4][3] ~^ image[21][3] + signed_kernel[4][4] ~^ image[21][4];
assign xor_sum[17][1] = signed_kernel[0][0] ~^ image[17][1] + signed_kernel[0][1] ~^ image[17][2] + signed_kernel[0][2] ~^ image[17][3] + signed_kernel[0][3] ~^ image[17][4] + signed_kernel[0][4] ~^ image[17][5] + signed_kernel[1][0] ~^ image[18][1] + signed_kernel[1][1] ~^ image[18][2] + signed_kernel[1][2] ~^ image[18][3] + signed_kernel[1][3] ~^ image[18][4] + signed_kernel[1][4] ~^ image[18][5] + signed_kernel[2][0] ~^ image[19][1] + signed_kernel[2][1] ~^ image[19][2] + signed_kernel[2][2] ~^ image[19][3] + signed_kernel[2][3] ~^ image[19][4] + signed_kernel[2][4] ~^ image[19][5] + signed_kernel[3][0] ~^ image[20][1] + signed_kernel[3][1] ~^ image[20][2] + signed_kernel[3][2] ~^ image[20][3] + signed_kernel[3][3] ~^ image[20][4] + signed_kernel[3][4] ~^ image[20][5] + signed_kernel[4][0] ~^ image[21][1] + signed_kernel[4][1] ~^ image[21][2] + signed_kernel[4][2] ~^ image[21][3] + signed_kernel[4][3] ~^ image[21][4] + signed_kernel[4][4] ~^ image[21][5];
assign xor_sum[17][2] = signed_kernel[0][0] ~^ image[17][2] + signed_kernel[0][1] ~^ image[17][3] + signed_kernel[0][2] ~^ image[17][4] + signed_kernel[0][3] ~^ image[17][5] + signed_kernel[0][4] ~^ image[17][6] + signed_kernel[1][0] ~^ image[18][2] + signed_kernel[1][1] ~^ image[18][3] + signed_kernel[1][2] ~^ image[18][4] + signed_kernel[1][3] ~^ image[18][5] + signed_kernel[1][4] ~^ image[18][6] + signed_kernel[2][0] ~^ image[19][2] + signed_kernel[2][1] ~^ image[19][3] + signed_kernel[2][2] ~^ image[19][4] + signed_kernel[2][3] ~^ image[19][5] + signed_kernel[2][4] ~^ image[19][6] + signed_kernel[3][0] ~^ image[20][2] + signed_kernel[3][1] ~^ image[20][3] + signed_kernel[3][2] ~^ image[20][4] + signed_kernel[3][3] ~^ image[20][5] + signed_kernel[3][4] ~^ image[20][6] + signed_kernel[4][0] ~^ image[21][2] + signed_kernel[4][1] ~^ image[21][3] + signed_kernel[4][2] ~^ image[21][4] + signed_kernel[4][3] ~^ image[21][5] + signed_kernel[4][4] ~^ image[21][6];
assign xor_sum[17][3] = signed_kernel[0][0] ~^ image[17][3] + signed_kernel[0][1] ~^ image[17][4] + signed_kernel[0][2] ~^ image[17][5] + signed_kernel[0][3] ~^ image[17][6] + signed_kernel[0][4] ~^ image[17][7] + signed_kernel[1][0] ~^ image[18][3] + signed_kernel[1][1] ~^ image[18][4] + signed_kernel[1][2] ~^ image[18][5] + signed_kernel[1][3] ~^ image[18][6] + signed_kernel[1][4] ~^ image[18][7] + signed_kernel[2][0] ~^ image[19][3] + signed_kernel[2][1] ~^ image[19][4] + signed_kernel[2][2] ~^ image[19][5] + signed_kernel[2][3] ~^ image[19][6] + signed_kernel[2][4] ~^ image[19][7] + signed_kernel[3][0] ~^ image[20][3] + signed_kernel[3][1] ~^ image[20][4] + signed_kernel[3][2] ~^ image[20][5] + signed_kernel[3][3] ~^ image[20][6] + signed_kernel[3][4] ~^ image[20][7] + signed_kernel[4][0] ~^ image[21][3] + signed_kernel[4][1] ~^ image[21][4] + signed_kernel[4][2] ~^ image[21][5] + signed_kernel[4][3] ~^ image[21][6] + signed_kernel[4][4] ~^ image[21][7];
assign xor_sum[17][4] = signed_kernel[0][0] ~^ image[17][4] + signed_kernel[0][1] ~^ image[17][5] + signed_kernel[0][2] ~^ image[17][6] + signed_kernel[0][3] ~^ image[17][7] + signed_kernel[0][4] ~^ image[17][8] + signed_kernel[1][0] ~^ image[18][4] + signed_kernel[1][1] ~^ image[18][5] + signed_kernel[1][2] ~^ image[18][6] + signed_kernel[1][3] ~^ image[18][7] + signed_kernel[1][4] ~^ image[18][8] + signed_kernel[2][0] ~^ image[19][4] + signed_kernel[2][1] ~^ image[19][5] + signed_kernel[2][2] ~^ image[19][6] + signed_kernel[2][3] ~^ image[19][7] + signed_kernel[2][4] ~^ image[19][8] + signed_kernel[3][0] ~^ image[20][4] + signed_kernel[3][1] ~^ image[20][5] + signed_kernel[3][2] ~^ image[20][6] + signed_kernel[3][3] ~^ image[20][7] + signed_kernel[3][4] ~^ image[20][8] + signed_kernel[4][0] ~^ image[21][4] + signed_kernel[4][1] ~^ image[21][5] + signed_kernel[4][2] ~^ image[21][6] + signed_kernel[4][3] ~^ image[21][7] + signed_kernel[4][4] ~^ image[21][8];
assign xor_sum[17][5] = signed_kernel[0][0] ~^ image[17][5] + signed_kernel[0][1] ~^ image[17][6] + signed_kernel[0][2] ~^ image[17][7] + signed_kernel[0][3] ~^ image[17][8] + signed_kernel[0][4] ~^ image[17][9] + signed_kernel[1][0] ~^ image[18][5] + signed_kernel[1][1] ~^ image[18][6] + signed_kernel[1][2] ~^ image[18][7] + signed_kernel[1][3] ~^ image[18][8] + signed_kernel[1][4] ~^ image[18][9] + signed_kernel[2][0] ~^ image[19][5] + signed_kernel[2][1] ~^ image[19][6] + signed_kernel[2][2] ~^ image[19][7] + signed_kernel[2][3] ~^ image[19][8] + signed_kernel[2][4] ~^ image[19][9] + signed_kernel[3][0] ~^ image[20][5] + signed_kernel[3][1] ~^ image[20][6] + signed_kernel[3][2] ~^ image[20][7] + signed_kernel[3][3] ~^ image[20][8] + signed_kernel[3][4] ~^ image[20][9] + signed_kernel[4][0] ~^ image[21][5] + signed_kernel[4][1] ~^ image[21][6] + signed_kernel[4][2] ~^ image[21][7] + signed_kernel[4][3] ~^ image[21][8] + signed_kernel[4][4] ~^ image[21][9];
assign xor_sum[17][6] = signed_kernel[0][0] ~^ image[17][6] + signed_kernel[0][1] ~^ image[17][7] + signed_kernel[0][2] ~^ image[17][8] + signed_kernel[0][3] ~^ image[17][9] + signed_kernel[0][4] ~^ image[17][10] + signed_kernel[1][0] ~^ image[18][6] + signed_kernel[1][1] ~^ image[18][7] + signed_kernel[1][2] ~^ image[18][8] + signed_kernel[1][3] ~^ image[18][9] + signed_kernel[1][4] ~^ image[18][10] + signed_kernel[2][0] ~^ image[19][6] + signed_kernel[2][1] ~^ image[19][7] + signed_kernel[2][2] ~^ image[19][8] + signed_kernel[2][3] ~^ image[19][9] + signed_kernel[2][4] ~^ image[19][10] + signed_kernel[3][0] ~^ image[20][6] + signed_kernel[3][1] ~^ image[20][7] + signed_kernel[3][2] ~^ image[20][8] + signed_kernel[3][3] ~^ image[20][9] + signed_kernel[3][4] ~^ image[20][10] + signed_kernel[4][0] ~^ image[21][6] + signed_kernel[4][1] ~^ image[21][7] + signed_kernel[4][2] ~^ image[21][8] + signed_kernel[4][3] ~^ image[21][9] + signed_kernel[4][4] ~^ image[21][10];
assign xor_sum[17][7] = signed_kernel[0][0] ~^ image[17][7] + signed_kernel[0][1] ~^ image[17][8] + signed_kernel[0][2] ~^ image[17][9] + signed_kernel[0][3] ~^ image[17][10] + signed_kernel[0][4] ~^ image[17][11] + signed_kernel[1][0] ~^ image[18][7] + signed_kernel[1][1] ~^ image[18][8] + signed_kernel[1][2] ~^ image[18][9] + signed_kernel[1][3] ~^ image[18][10] + signed_kernel[1][4] ~^ image[18][11] + signed_kernel[2][0] ~^ image[19][7] + signed_kernel[2][1] ~^ image[19][8] + signed_kernel[2][2] ~^ image[19][9] + signed_kernel[2][3] ~^ image[19][10] + signed_kernel[2][4] ~^ image[19][11] + signed_kernel[3][0] ~^ image[20][7] + signed_kernel[3][1] ~^ image[20][8] + signed_kernel[3][2] ~^ image[20][9] + signed_kernel[3][3] ~^ image[20][10] + signed_kernel[3][4] ~^ image[20][11] + signed_kernel[4][0] ~^ image[21][7] + signed_kernel[4][1] ~^ image[21][8] + signed_kernel[4][2] ~^ image[21][9] + signed_kernel[4][3] ~^ image[21][10] + signed_kernel[4][4] ~^ image[21][11];
assign xor_sum[17][8] = signed_kernel[0][0] ~^ image[17][8] + signed_kernel[0][1] ~^ image[17][9] + signed_kernel[0][2] ~^ image[17][10] + signed_kernel[0][3] ~^ image[17][11] + signed_kernel[0][4] ~^ image[17][12] + signed_kernel[1][0] ~^ image[18][8] + signed_kernel[1][1] ~^ image[18][9] + signed_kernel[1][2] ~^ image[18][10] + signed_kernel[1][3] ~^ image[18][11] + signed_kernel[1][4] ~^ image[18][12] + signed_kernel[2][0] ~^ image[19][8] + signed_kernel[2][1] ~^ image[19][9] + signed_kernel[2][2] ~^ image[19][10] + signed_kernel[2][3] ~^ image[19][11] + signed_kernel[2][4] ~^ image[19][12] + signed_kernel[3][0] ~^ image[20][8] + signed_kernel[3][1] ~^ image[20][9] + signed_kernel[3][2] ~^ image[20][10] + signed_kernel[3][3] ~^ image[20][11] + signed_kernel[3][4] ~^ image[20][12] + signed_kernel[4][0] ~^ image[21][8] + signed_kernel[4][1] ~^ image[21][9] + signed_kernel[4][2] ~^ image[21][10] + signed_kernel[4][3] ~^ image[21][11] + signed_kernel[4][4] ~^ image[21][12];
assign xor_sum[17][9] = signed_kernel[0][0] ~^ image[17][9] + signed_kernel[0][1] ~^ image[17][10] + signed_kernel[0][2] ~^ image[17][11] + signed_kernel[0][3] ~^ image[17][12] + signed_kernel[0][4] ~^ image[17][13] + signed_kernel[1][0] ~^ image[18][9] + signed_kernel[1][1] ~^ image[18][10] + signed_kernel[1][2] ~^ image[18][11] + signed_kernel[1][3] ~^ image[18][12] + signed_kernel[1][4] ~^ image[18][13] + signed_kernel[2][0] ~^ image[19][9] + signed_kernel[2][1] ~^ image[19][10] + signed_kernel[2][2] ~^ image[19][11] + signed_kernel[2][3] ~^ image[19][12] + signed_kernel[2][4] ~^ image[19][13] + signed_kernel[3][0] ~^ image[20][9] + signed_kernel[3][1] ~^ image[20][10] + signed_kernel[3][2] ~^ image[20][11] + signed_kernel[3][3] ~^ image[20][12] + signed_kernel[3][4] ~^ image[20][13] + signed_kernel[4][0] ~^ image[21][9] + signed_kernel[4][1] ~^ image[21][10] + signed_kernel[4][2] ~^ image[21][11] + signed_kernel[4][3] ~^ image[21][12] + signed_kernel[4][4] ~^ image[21][13];
assign xor_sum[17][10] = signed_kernel[0][0] ~^ image[17][10] + signed_kernel[0][1] ~^ image[17][11] + signed_kernel[0][2] ~^ image[17][12] + signed_kernel[0][3] ~^ image[17][13] + signed_kernel[0][4] ~^ image[17][14] + signed_kernel[1][0] ~^ image[18][10] + signed_kernel[1][1] ~^ image[18][11] + signed_kernel[1][2] ~^ image[18][12] + signed_kernel[1][3] ~^ image[18][13] + signed_kernel[1][4] ~^ image[18][14] + signed_kernel[2][0] ~^ image[19][10] + signed_kernel[2][1] ~^ image[19][11] + signed_kernel[2][2] ~^ image[19][12] + signed_kernel[2][3] ~^ image[19][13] + signed_kernel[2][4] ~^ image[19][14] + signed_kernel[3][0] ~^ image[20][10] + signed_kernel[3][1] ~^ image[20][11] + signed_kernel[3][2] ~^ image[20][12] + signed_kernel[3][3] ~^ image[20][13] + signed_kernel[3][4] ~^ image[20][14] + signed_kernel[4][0] ~^ image[21][10] + signed_kernel[4][1] ~^ image[21][11] + signed_kernel[4][2] ~^ image[21][12] + signed_kernel[4][3] ~^ image[21][13] + signed_kernel[4][4] ~^ image[21][14];
assign xor_sum[17][11] = signed_kernel[0][0] ~^ image[17][11] + signed_kernel[0][1] ~^ image[17][12] + signed_kernel[0][2] ~^ image[17][13] + signed_kernel[0][3] ~^ image[17][14] + signed_kernel[0][4] ~^ image[17][15] + signed_kernel[1][0] ~^ image[18][11] + signed_kernel[1][1] ~^ image[18][12] + signed_kernel[1][2] ~^ image[18][13] + signed_kernel[1][3] ~^ image[18][14] + signed_kernel[1][4] ~^ image[18][15] + signed_kernel[2][0] ~^ image[19][11] + signed_kernel[2][1] ~^ image[19][12] + signed_kernel[2][2] ~^ image[19][13] + signed_kernel[2][3] ~^ image[19][14] + signed_kernel[2][4] ~^ image[19][15] + signed_kernel[3][0] ~^ image[20][11] + signed_kernel[3][1] ~^ image[20][12] + signed_kernel[3][2] ~^ image[20][13] + signed_kernel[3][3] ~^ image[20][14] + signed_kernel[3][4] ~^ image[20][15] + signed_kernel[4][0] ~^ image[21][11] + signed_kernel[4][1] ~^ image[21][12] + signed_kernel[4][2] ~^ image[21][13] + signed_kernel[4][3] ~^ image[21][14] + signed_kernel[4][4] ~^ image[21][15];
assign xor_sum[17][12] = signed_kernel[0][0] ~^ image[17][12] + signed_kernel[0][1] ~^ image[17][13] + signed_kernel[0][2] ~^ image[17][14] + signed_kernel[0][3] ~^ image[17][15] + signed_kernel[0][4] ~^ image[17][16] + signed_kernel[1][0] ~^ image[18][12] + signed_kernel[1][1] ~^ image[18][13] + signed_kernel[1][2] ~^ image[18][14] + signed_kernel[1][3] ~^ image[18][15] + signed_kernel[1][4] ~^ image[18][16] + signed_kernel[2][0] ~^ image[19][12] + signed_kernel[2][1] ~^ image[19][13] + signed_kernel[2][2] ~^ image[19][14] + signed_kernel[2][3] ~^ image[19][15] + signed_kernel[2][4] ~^ image[19][16] + signed_kernel[3][0] ~^ image[20][12] + signed_kernel[3][1] ~^ image[20][13] + signed_kernel[3][2] ~^ image[20][14] + signed_kernel[3][3] ~^ image[20][15] + signed_kernel[3][4] ~^ image[20][16] + signed_kernel[4][0] ~^ image[21][12] + signed_kernel[4][1] ~^ image[21][13] + signed_kernel[4][2] ~^ image[21][14] + signed_kernel[4][3] ~^ image[21][15] + signed_kernel[4][4] ~^ image[21][16];
assign xor_sum[17][13] = signed_kernel[0][0] ~^ image[17][13] + signed_kernel[0][1] ~^ image[17][14] + signed_kernel[0][2] ~^ image[17][15] + signed_kernel[0][3] ~^ image[17][16] + signed_kernel[0][4] ~^ image[17][17] + signed_kernel[1][0] ~^ image[18][13] + signed_kernel[1][1] ~^ image[18][14] + signed_kernel[1][2] ~^ image[18][15] + signed_kernel[1][3] ~^ image[18][16] + signed_kernel[1][4] ~^ image[18][17] + signed_kernel[2][0] ~^ image[19][13] + signed_kernel[2][1] ~^ image[19][14] + signed_kernel[2][2] ~^ image[19][15] + signed_kernel[2][3] ~^ image[19][16] + signed_kernel[2][4] ~^ image[19][17] + signed_kernel[3][0] ~^ image[20][13] + signed_kernel[3][1] ~^ image[20][14] + signed_kernel[3][2] ~^ image[20][15] + signed_kernel[3][3] ~^ image[20][16] + signed_kernel[3][4] ~^ image[20][17] + signed_kernel[4][0] ~^ image[21][13] + signed_kernel[4][1] ~^ image[21][14] + signed_kernel[4][2] ~^ image[21][15] + signed_kernel[4][3] ~^ image[21][16] + signed_kernel[4][4] ~^ image[21][17];
assign xor_sum[17][14] = signed_kernel[0][0] ~^ image[17][14] + signed_kernel[0][1] ~^ image[17][15] + signed_kernel[0][2] ~^ image[17][16] + signed_kernel[0][3] ~^ image[17][17] + signed_kernel[0][4] ~^ image[17][18] + signed_kernel[1][0] ~^ image[18][14] + signed_kernel[1][1] ~^ image[18][15] + signed_kernel[1][2] ~^ image[18][16] + signed_kernel[1][3] ~^ image[18][17] + signed_kernel[1][4] ~^ image[18][18] + signed_kernel[2][0] ~^ image[19][14] + signed_kernel[2][1] ~^ image[19][15] + signed_kernel[2][2] ~^ image[19][16] + signed_kernel[2][3] ~^ image[19][17] + signed_kernel[2][4] ~^ image[19][18] + signed_kernel[3][0] ~^ image[20][14] + signed_kernel[3][1] ~^ image[20][15] + signed_kernel[3][2] ~^ image[20][16] + signed_kernel[3][3] ~^ image[20][17] + signed_kernel[3][4] ~^ image[20][18] + signed_kernel[4][0] ~^ image[21][14] + signed_kernel[4][1] ~^ image[21][15] + signed_kernel[4][2] ~^ image[21][16] + signed_kernel[4][3] ~^ image[21][17] + signed_kernel[4][4] ~^ image[21][18];
assign xor_sum[17][15] = signed_kernel[0][0] ~^ image[17][15] + signed_kernel[0][1] ~^ image[17][16] + signed_kernel[0][2] ~^ image[17][17] + signed_kernel[0][3] ~^ image[17][18] + signed_kernel[0][4] ~^ image[17][19] + signed_kernel[1][0] ~^ image[18][15] + signed_kernel[1][1] ~^ image[18][16] + signed_kernel[1][2] ~^ image[18][17] + signed_kernel[1][3] ~^ image[18][18] + signed_kernel[1][4] ~^ image[18][19] + signed_kernel[2][0] ~^ image[19][15] + signed_kernel[2][1] ~^ image[19][16] + signed_kernel[2][2] ~^ image[19][17] + signed_kernel[2][3] ~^ image[19][18] + signed_kernel[2][4] ~^ image[19][19] + signed_kernel[3][0] ~^ image[20][15] + signed_kernel[3][1] ~^ image[20][16] + signed_kernel[3][2] ~^ image[20][17] + signed_kernel[3][3] ~^ image[20][18] + signed_kernel[3][4] ~^ image[20][19] + signed_kernel[4][0] ~^ image[21][15] + signed_kernel[4][1] ~^ image[21][16] + signed_kernel[4][2] ~^ image[21][17] + signed_kernel[4][3] ~^ image[21][18] + signed_kernel[4][4] ~^ image[21][19];
assign xor_sum[17][16] = signed_kernel[0][0] ~^ image[17][16] + signed_kernel[0][1] ~^ image[17][17] + signed_kernel[0][2] ~^ image[17][18] + signed_kernel[0][3] ~^ image[17][19] + signed_kernel[0][4] ~^ image[17][20] + signed_kernel[1][0] ~^ image[18][16] + signed_kernel[1][1] ~^ image[18][17] + signed_kernel[1][2] ~^ image[18][18] + signed_kernel[1][3] ~^ image[18][19] + signed_kernel[1][4] ~^ image[18][20] + signed_kernel[2][0] ~^ image[19][16] + signed_kernel[2][1] ~^ image[19][17] + signed_kernel[2][2] ~^ image[19][18] + signed_kernel[2][3] ~^ image[19][19] + signed_kernel[2][4] ~^ image[19][20] + signed_kernel[3][0] ~^ image[20][16] + signed_kernel[3][1] ~^ image[20][17] + signed_kernel[3][2] ~^ image[20][18] + signed_kernel[3][3] ~^ image[20][19] + signed_kernel[3][4] ~^ image[20][20] + signed_kernel[4][0] ~^ image[21][16] + signed_kernel[4][1] ~^ image[21][17] + signed_kernel[4][2] ~^ image[21][18] + signed_kernel[4][3] ~^ image[21][19] + signed_kernel[4][4] ~^ image[21][20];
assign xor_sum[17][17] = signed_kernel[0][0] ~^ image[17][17] + signed_kernel[0][1] ~^ image[17][18] + signed_kernel[0][2] ~^ image[17][19] + signed_kernel[0][3] ~^ image[17][20] + signed_kernel[0][4] ~^ image[17][21] + signed_kernel[1][0] ~^ image[18][17] + signed_kernel[1][1] ~^ image[18][18] + signed_kernel[1][2] ~^ image[18][19] + signed_kernel[1][3] ~^ image[18][20] + signed_kernel[1][4] ~^ image[18][21] + signed_kernel[2][0] ~^ image[19][17] + signed_kernel[2][1] ~^ image[19][18] + signed_kernel[2][2] ~^ image[19][19] + signed_kernel[2][3] ~^ image[19][20] + signed_kernel[2][4] ~^ image[19][21] + signed_kernel[3][0] ~^ image[20][17] + signed_kernel[3][1] ~^ image[20][18] + signed_kernel[3][2] ~^ image[20][19] + signed_kernel[3][3] ~^ image[20][20] + signed_kernel[3][4] ~^ image[20][21] + signed_kernel[4][0] ~^ image[21][17] + signed_kernel[4][1] ~^ image[21][18] + signed_kernel[4][2] ~^ image[21][19] + signed_kernel[4][3] ~^ image[21][20] + signed_kernel[4][4] ~^ image[21][21];
assign xor_sum[17][18] = signed_kernel[0][0] ~^ image[17][18] + signed_kernel[0][1] ~^ image[17][19] + signed_kernel[0][2] ~^ image[17][20] + signed_kernel[0][3] ~^ image[17][21] + signed_kernel[0][4] ~^ image[17][22] + signed_kernel[1][0] ~^ image[18][18] + signed_kernel[1][1] ~^ image[18][19] + signed_kernel[1][2] ~^ image[18][20] + signed_kernel[1][3] ~^ image[18][21] + signed_kernel[1][4] ~^ image[18][22] + signed_kernel[2][0] ~^ image[19][18] + signed_kernel[2][1] ~^ image[19][19] + signed_kernel[2][2] ~^ image[19][20] + signed_kernel[2][3] ~^ image[19][21] + signed_kernel[2][4] ~^ image[19][22] + signed_kernel[3][0] ~^ image[20][18] + signed_kernel[3][1] ~^ image[20][19] + signed_kernel[3][2] ~^ image[20][20] + signed_kernel[3][3] ~^ image[20][21] + signed_kernel[3][4] ~^ image[20][22] + signed_kernel[4][0] ~^ image[21][18] + signed_kernel[4][1] ~^ image[21][19] + signed_kernel[4][2] ~^ image[21][20] + signed_kernel[4][3] ~^ image[21][21] + signed_kernel[4][4] ~^ image[21][22];
assign xor_sum[17][19] = signed_kernel[0][0] ~^ image[17][19] + signed_kernel[0][1] ~^ image[17][20] + signed_kernel[0][2] ~^ image[17][21] + signed_kernel[0][3] ~^ image[17][22] + signed_kernel[0][4] ~^ image[17][23] + signed_kernel[1][0] ~^ image[18][19] + signed_kernel[1][1] ~^ image[18][20] + signed_kernel[1][2] ~^ image[18][21] + signed_kernel[1][3] ~^ image[18][22] + signed_kernel[1][4] ~^ image[18][23] + signed_kernel[2][0] ~^ image[19][19] + signed_kernel[2][1] ~^ image[19][20] + signed_kernel[2][2] ~^ image[19][21] + signed_kernel[2][3] ~^ image[19][22] + signed_kernel[2][4] ~^ image[19][23] + signed_kernel[3][0] ~^ image[20][19] + signed_kernel[3][1] ~^ image[20][20] + signed_kernel[3][2] ~^ image[20][21] + signed_kernel[3][3] ~^ image[20][22] + signed_kernel[3][4] ~^ image[20][23] + signed_kernel[4][0] ~^ image[21][19] + signed_kernel[4][1] ~^ image[21][20] + signed_kernel[4][2] ~^ image[21][21] + signed_kernel[4][3] ~^ image[21][22] + signed_kernel[4][4] ~^ image[21][23];
assign xor_sum[17][20] = signed_kernel[0][0] ~^ image[17][20] + signed_kernel[0][1] ~^ image[17][21] + signed_kernel[0][2] ~^ image[17][22] + signed_kernel[0][3] ~^ image[17][23] + signed_kernel[0][4] ~^ image[17][24] + signed_kernel[1][0] ~^ image[18][20] + signed_kernel[1][1] ~^ image[18][21] + signed_kernel[1][2] ~^ image[18][22] + signed_kernel[1][3] ~^ image[18][23] + signed_kernel[1][4] ~^ image[18][24] + signed_kernel[2][0] ~^ image[19][20] + signed_kernel[2][1] ~^ image[19][21] + signed_kernel[2][2] ~^ image[19][22] + signed_kernel[2][3] ~^ image[19][23] + signed_kernel[2][4] ~^ image[19][24] + signed_kernel[3][0] ~^ image[20][20] + signed_kernel[3][1] ~^ image[20][21] + signed_kernel[3][2] ~^ image[20][22] + signed_kernel[3][3] ~^ image[20][23] + signed_kernel[3][4] ~^ image[20][24] + signed_kernel[4][0] ~^ image[21][20] + signed_kernel[4][1] ~^ image[21][21] + signed_kernel[4][2] ~^ image[21][22] + signed_kernel[4][3] ~^ image[21][23] + signed_kernel[4][4] ~^ image[21][24];
assign xor_sum[17][21] = signed_kernel[0][0] ~^ image[17][21] + signed_kernel[0][1] ~^ image[17][22] + signed_kernel[0][2] ~^ image[17][23] + signed_kernel[0][3] ~^ image[17][24] + signed_kernel[0][4] ~^ image[17][25] + signed_kernel[1][0] ~^ image[18][21] + signed_kernel[1][1] ~^ image[18][22] + signed_kernel[1][2] ~^ image[18][23] + signed_kernel[1][3] ~^ image[18][24] + signed_kernel[1][4] ~^ image[18][25] + signed_kernel[2][0] ~^ image[19][21] + signed_kernel[2][1] ~^ image[19][22] + signed_kernel[2][2] ~^ image[19][23] + signed_kernel[2][3] ~^ image[19][24] + signed_kernel[2][4] ~^ image[19][25] + signed_kernel[3][0] ~^ image[20][21] + signed_kernel[3][1] ~^ image[20][22] + signed_kernel[3][2] ~^ image[20][23] + signed_kernel[3][3] ~^ image[20][24] + signed_kernel[3][4] ~^ image[20][25] + signed_kernel[4][0] ~^ image[21][21] + signed_kernel[4][1] ~^ image[21][22] + signed_kernel[4][2] ~^ image[21][23] + signed_kernel[4][3] ~^ image[21][24] + signed_kernel[4][4] ~^ image[21][25];
assign xor_sum[17][22] = signed_kernel[0][0] ~^ image[17][22] + signed_kernel[0][1] ~^ image[17][23] + signed_kernel[0][2] ~^ image[17][24] + signed_kernel[0][3] ~^ image[17][25] + signed_kernel[0][4] ~^ image[17][26] + signed_kernel[1][0] ~^ image[18][22] + signed_kernel[1][1] ~^ image[18][23] + signed_kernel[1][2] ~^ image[18][24] + signed_kernel[1][3] ~^ image[18][25] + signed_kernel[1][4] ~^ image[18][26] + signed_kernel[2][0] ~^ image[19][22] + signed_kernel[2][1] ~^ image[19][23] + signed_kernel[2][2] ~^ image[19][24] + signed_kernel[2][3] ~^ image[19][25] + signed_kernel[2][4] ~^ image[19][26] + signed_kernel[3][0] ~^ image[20][22] + signed_kernel[3][1] ~^ image[20][23] + signed_kernel[3][2] ~^ image[20][24] + signed_kernel[3][3] ~^ image[20][25] + signed_kernel[3][4] ~^ image[20][26] + signed_kernel[4][0] ~^ image[21][22] + signed_kernel[4][1] ~^ image[21][23] + signed_kernel[4][2] ~^ image[21][24] + signed_kernel[4][3] ~^ image[21][25] + signed_kernel[4][4] ~^ image[21][26];
assign xor_sum[17][23] = signed_kernel[0][0] ~^ image[17][23] + signed_kernel[0][1] ~^ image[17][24] + signed_kernel[0][2] ~^ image[17][25] + signed_kernel[0][3] ~^ image[17][26] + signed_kernel[0][4] ~^ image[17][27] + signed_kernel[1][0] ~^ image[18][23] + signed_kernel[1][1] ~^ image[18][24] + signed_kernel[1][2] ~^ image[18][25] + signed_kernel[1][3] ~^ image[18][26] + signed_kernel[1][4] ~^ image[18][27] + signed_kernel[2][0] ~^ image[19][23] + signed_kernel[2][1] ~^ image[19][24] + signed_kernel[2][2] ~^ image[19][25] + signed_kernel[2][3] ~^ image[19][26] + signed_kernel[2][4] ~^ image[19][27] + signed_kernel[3][0] ~^ image[20][23] + signed_kernel[3][1] ~^ image[20][24] + signed_kernel[3][2] ~^ image[20][25] + signed_kernel[3][3] ~^ image[20][26] + signed_kernel[3][4] ~^ image[20][27] + signed_kernel[4][0] ~^ image[21][23] + signed_kernel[4][1] ~^ image[21][24] + signed_kernel[4][2] ~^ image[21][25] + signed_kernel[4][3] ~^ image[21][26] + signed_kernel[4][4] ~^ image[21][27];
assign xor_sum[18][0] = signed_kernel[0][0] ~^ image[18][0] + signed_kernel[0][1] ~^ image[18][1] + signed_kernel[0][2] ~^ image[18][2] + signed_kernel[0][3] ~^ image[18][3] + signed_kernel[0][4] ~^ image[18][4] + signed_kernel[1][0] ~^ image[19][0] + signed_kernel[1][1] ~^ image[19][1] + signed_kernel[1][2] ~^ image[19][2] + signed_kernel[1][3] ~^ image[19][3] + signed_kernel[1][4] ~^ image[19][4] + signed_kernel[2][0] ~^ image[20][0] + signed_kernel[2][1] ~^ image[20][1] + signed_kernel[2][2] ~^ image[20][2] + signed_kernel[2][3] ~^ image[20][3] + signed_kernel[2][4] ~^ image[20][4] + signed_kernel[3][0] ~^ image[21][0] + signed_kernel[3][1] ~^ image[21][1] + signed_kernel[3][2] ~^ image[21][2] + signed_kernel[3][3] ~^ image[21][3] + signed_kernel[3][4] ~^ image[21][4] + signed_kernel[4][0] ~^ image[22][0] + signed_kernel[4][1] ~^ image[22][1] + signed_kernel[4][2] ~^ image[22][2] + signed_kernel[4][3] ~^ image[22][3] + signed_kernel[4][4] ~^ image[22][4];
assign xor_sum[18][1] = signed_kernel[0][0] ~^ image[18][1] + signed_kernel[0][1] ~^ image[18][2] + signed_kernel[0][2] ~^ image[18][3] + signed_kernel[0][3] ~^ image[18][4] + signed_kernel[0][4] ~^ image[18][5] + signed_kernel[1][0] ~^ image[19][1] + signed_kernel[1][1] ~^ image[19][2] + signed_kernel[1][2] ~^ image[19][3] + signed_kernel[1][3] ~^ image[19][4] + signed_kernel[1][4] ~^ image[19][5] + signed_kernel[2][0] ~^ image[20][1] + signed_kernel[2][1] ~^ image[20][2] + signed_kernel[2][2] ~^ image[20][3] + signed_kernel[2][3] ~^ image[20][4] + signed_kernel[2][4] ~^ image[20][5] + signed_kernel[3][0] ~^ image[21][1] + signed_kernel[3][1] ~^ image[21][2] + signed_kernel[3][2] ~^ image[21][3] + signed_kernel[3][3] ~^ image[21][4] + signed_kernel[3][4] ~^ image[21][5] + signed_kernel[4][0] ~^ image[22][1] + signed_kernel[4][1] ~^ image[22][2] + signed_kernel[4][2] ~^ image[22][3] + signed_kernel[4][3] ~^ image[22][4] + signed_kernel[4][4] ~^ image[22][5];
assign xor_sum[18][2] = signed_kernel[0][0] ~^ image[18][2] + signed_kernel[0][1] ~^ image[18][3] + signed_kernel[0][2] ~^ image[18][4] + signed_kernel[0][3] ~^ image[18][5] + signed_kernel[0][4] ~^ image[18][6] + signed_kernel[1][0] ~^ image[19][2] + signed_kernel[1][1] ~^ image[19][3] + signed_kernel[1][2] ~^ image[19][4] + signed_kernel[1][3] ~^ image[19][5] + signed_kernel[1][4] ~^ image[19][6] + signed_kernel[2][0] ~^ image[20][2] + signed_kernel[2][1] ~^ image[20][3] + signed_kernel[2][2] ~^ image[20][4] + signed_kernel[2][3] ~^ image[20][5] + signed_kernel[2][4] ~^ image[20][6] + signed_kernel[3][0] ~^ image[21][2] + signed_kernel[3][1] ~^ image[21][3] + signed_kernel[3][2] ~^ image[21][4] + signed_kernel[3][3] ~^ image[21][5] + signed_kernel[3][4] ~^ image[21][6] + signed_kernel[4][0] ~^ image[22][2] + signed_kernel[4][1] ~^ image[22][3] + signed_kernel[4][2] ~^ image[22][4] + signed_kernel[4][3] ~^ image[22][5] + signed_kernel[4][4] ~^ image[22][6];
assign xor_sum[18][3] = signed_kernel[0][0] ~^ image[18][3] + signed_kernel[0][1] ~^ image[18][4] + signed_kernel[0][2] ~^ image[18][5] + signed_kernel[0][3] ~^ image[18][6] + signed_kernel[0][4] ~^ image[18][7] + signed_kernel[1][0] ~^ image[19][3] + signed_kernel[1][1] ~^ image[19][4] + signed_kernel[1][2] ~^ image[19][5] + signed_kernel[1][3] ~^ image[19][6] + signed_kernel[1][4] ~^ image[19][7] + signed_kernel[2][0] ~^ image[20][3] + signed_kernel[2][1] ~^ image[20][4] + signed_kernel[2][2] ~^ image[20][5] + signed_kernel[2][3] ~^ image[20][6] + signed_kernel[2][4] ~^ image[20][7] + signed_kernel[3][0] ~^ image[21][3] + signed_kernel[3][1] ~^ image[21][4] + signed_kernel[3][2] ~^ image[21][5] + signed_kernel[3][3] ~^ image[21][6] + signed_kernel[3][4] ~^ image[21][7] + signed_kernel[4][0] ~^ image[22][3] + signed_kernel[4][1] ~^ image[22][4] + signed_kernel[4][2] ~^ image[22][5] + signed_kernel[4][3] ~^ image[22][6] + signed_kernel[4][4] ~^ image[22][7];
assign xor_sum[18][4] = signed_kernel[0][0] ~^ image[18][4] + signed_kernel[0][1] ~^ image[18][5] + signed_kernel[0][2] ~^ image[18][6] + signed_kernel[0][3] ~^ image[18][7] + signed_kernel[0][4] ~^ image[18][8] + signed_kernel[1][0] ~^ image[19][4] + signed_kernel[1][1] ~^ image[19][5] + signed_kernel[1][2] ~^ image[19][6] + signed_kernel[1][3] ~^ image[19][7] + signed_kernel[1][4] ~^ image[19][8] + signed_kernel[2][0] ~^ image[20][4] + signed_kernel[2][1] ~^ image[20][5] + signed_kernel[2][2] ~^ image[20][6] + signed_kernel[2][3] ~^ image[20][7] + signed_kernel[2][4] ~^ image[20][8] + signed_kernel[3][0] ~^ image[21][4] + signed_kernel[3][1] ~^ image[21][5] + signed_kernel[3][2] ~^ image[21][6] + signed_kernel[3][3] ~^ image[21][7] + signed_kernel[3][4] ~^ image[21][8] + signed_kernel[4][0] ~^ image[22][4] + signed_kernel[4][1] ~^ image[22][5] + signed_kernel[4][2] ~^ image[22][6] + signed_kernel[4][3] ~^ image[22][7] + signed_kernel[4][4] ~^ image[22][8];
assign xor_sum[18][5] = signed_kernel[0][0] ~^ image[18][5] + signed_kernel[0][1] ~^ image[18][6] + signed_kernel[0][2] ~^ image[18][7] + signed_kernel[0][3] ~^ image[18][8] + signed_kernel[0][4] ~^ image[18][9] + signed_kernel[1][0] ~^ image[19][5] + signed_kernel[1][1] ~^ image[19][6] + signed_kernel[1][2] ~^ image[19][7] + signed_kernel[1][3] ~^ image[19][8] + signed_kernel[1][4] ~^ image[19][9] + signed_kernel[2][0] ~^ image[20][5] + signed_kernel[2][1] ~^ image[20][6] + signed_kernel[2][2] ~^ image[20][7] + signed_kernel[2][3] ~^ image[20][8] + signed_kernel[2][4] ~^ image[20][9] + signed_kernel[3][0] ~^ image[21][5] + signed_kernel[3][1] ~^ image[21][6] + signed_kernel[3][2] ~^ image[21][7] + signed_kernel[3][3] ~^ image[21][8] + signed_kernel[3][4] ~^ image[21][9] + signed_kernel[4][0] ~^ image[22][5] + signed_kernel[4][1] ~^ image[22][6] + signed_kernel[4][2] ~^ image[22][7] + signed_kernel[4][3] ~^ image[22][8] + signed_kernel[4][4] ~^ image[22][9];
assign xor_sum[18][6] = signed_kernel[0][0] ~^ image[18][6] + signed_kernel[0][1] ~^ image[18][7] + signed_kernel[0][2] ~^ image[18][8] + signed_kernel[0][3] ~^ image[18][9] + signed_kernel[0][4] ~^ image[18][10] + signed_kernel[1][0] ~^ image[19][6] + signed_kernel[1][1] ~^ image[19][7] + signed_kernel[1][2] ~^ image[19][8] + signed_kernel[1][3] ~^ image[19][9] + signed_kernel[1][4] ~^ image[19][10] + signed_kernel[2][0] ~^ image[20][6] + signed_kernel[2][1] ~^ image[20][7] + signed_kernel[2][2] ~^ image[20][8] + signed_kernel[2][3] ~^ image[20][9] + signed_kernel[2][4] ~^ image[20][10] + signed_kernel[3][0] ~^ image[21][6] + signed_kernel[3][1] ~^ image[21][7] + signed_kernel[3][2] ~^ image[21][8] + signed_kernel[3][3] ~^ image[21][9] + signed_kernel[3][4] ~^ image[21][10] + signed_kernel[4][0] ~^ image[22][6] + signed_kernel[4][1] ~^ image[22][7] + signed_kernel[4][2] ~^ image[22][8] + signed_kernel[4][3] ~^ image[22][9] + signed_kernel[4][4] ~^ image[22][10];
assign xor_sum[18][7] = signed_kernel[0][0] ~^ image[18][7] + signed_kernel[0][1] ~^ image[18][8] + signed_kernel[0][2] ~^ image[18][9] + signed_kernel[0][3] ~^ image[18][10] + signed_kernel[0][4] ~^ image[18][11] + signed_kernel[1][0] ~^ image[19][7] + signed_kernel[1][1] ~^ image[19][8] + signed_kernel[1][2] ~^ image[19][9] + signed_kernel[1][3] ~^ image[19][10] + signed_kernel[1][4] ~^ image[19][11] + signed_kernel[2][0] ~^ image[20][7] + signed_kernel[2][1] ~^ image[20][8] + signed_kernel[2][2] ~^ image[20][9] + signed_kernel[2][3] ~^ image[20][10] + signed_kernel[2][4] ~^ image[20][11] + signed_kernel[3][0] ~^ image[21][7] + signed_kernel[3][1] ~^ image[21][8] + signed_kernel[3][2] ~^ image[21][9] + signed_kernel[3][3] ~^ image[21][10] + signed_kernel[3][4] ~^ image[21][11] + signed_kernel[4][0] ~^ image[22][7] + signed_kernel[4][1] ~^ image[22][8] + signed_kernel[4][2] ~^ image[22][9] + signed_kernel[4][3] ~^ image[22][10] + signed_kernel[4][4] ~^ image[22][11];
assign xor_sum[18][8] = signed_kernel[0][0] ~^ image[18][8] + signed_kernel[0][1] ~^ image[18][9] + signed_kernel[0][2] ~^ image[18][10] + signed_kernel[0][3] ~^ image[18][11] + signed_kernel[0][4] ~^ image[18][12] + signed_kernel[1][0] ~^ image[19][8] + signed_kernel[1][1] ~^ image[19][9] + signed_kernel[1][2] ~^ image[19][10] + signed_kernel[1][3] ~^ image[19][11] + signed_kernel[1][4] ~^ image[19][12] + signed_kernel[2][0] ~^ image[20][8] + signed_kernel[2][1] ~^ image[20][9] + signed_kernel[2][2] ~^ image[20][10] + signed_kernel[2][3] ~^ image[20][11] + signed_kernel[2][4] ~^ image[20][12] + signed_kernel[3][0] ~^ image[21][8] + signed_kernel[3][1] ~^ image[21][9] + signed_kernel[3][2] ~^ image[21][10] + signed_kernel[3][3] ~^ image[21][11] + signed_kernel[3][4] ~^ image[21][12] + signed_kernel[4][0] ~^ image[22][8] + signed_kernel[4][1] ~^ image[22][9] + signed_kernel[4][2] ~^ image[22][10] + signed_kernel[4][3] ~^ image[22][11] + signed_kernel[4][4] ~^ image[22][12];
assign xor_sum[18][9] = signed_kernel[0][0] ~^ image[18][9] + signed_kernel[0][1] ~^ image[18][10] + signed_kernel[0][2] ~^ image[18][11] + signed_kernel[0][3] ~^ image[18][12] + signed_kernel[0][4] ~^ image[18][13] + signed_kernel[1][0] ~^ image[19][9] + signed_kernel[1][1] ~^ image[19][10] + signed_kernel[1][2] ~^ image[19][11] + signed_kernel[1][3] ~^ image[19][12] + signed_kernel[1][4] ~^ image[19][13] + signed_kernel[2][0] ~^ image[20][9] + signed_kernel[2][1] ~^ image[20][10] + signed_kernel[2][2] ~^ image[20][11] + signed_kernel[2][3] ~^ image[20][12] + signed_kernel[2][4] ~^ image[20][13] + signed_kernel[3][0] ~^ image[21][9] + signed_kernel[3][1] ~^ image[21][10] + signed_kernel[3][2] ~^ image[21][11] + signed_kernel[3][3] ~^ image[21][12] + signed_kernel[3][4] ~^ image[21][13] + signed_kernel[4][0] ~^ image[22][9] + signed_kernel[4][1] ~^ image[22][10] + signed_kernel[4][2] ~^ image[22][11] + signed_kernel[4][3] ~^ image[22][12] + signed_kernel[4][4] ~^ image[22][13];
assign xor_sum[18][10] = signed_kernel[0][0] ~^ image[18][10] + signed_kernel[0][1] ~^ image[18][11] + signed_kernel[0][2] ~^ image[18][12] + signed_kernel[0][3] ~^ image[18][13] + signed_kernel[0][4] ~^ image[18][14] + signed_kernel[1][0] ~^ image[19][10] + signed_kernel[1][1] ~^ image[19][11] + signed_kernel[1][2] ~^ image[19][12] + signed_kernel[1][3] ~^ image[19][13] + signed_kernel[1][4] ~^ image[19][14] + signed_kernel[2][0] ~^ image[20][10] + signed_kernel[2][1] ~^ image[20][11] + signed_kernel[2][2] ~^ image[20][12] + signed_kernel[2][3] ~^ image[20][13] + signed_kernel[2][4] ~^ image[20][14] + signed_kernel[3][0] ~^ image[21][10] + signed_kernel[3][1] ~^ image[21][11] + signed_kernel[3][2] ~^ image[21][12] + signed_kernel[3][3] ~^ image[21][13] + signed_kernel[3][4] ~^ image[21][14] + signed_kernel[4][0] ~^ image[22][10] + signed_kernel[4][1] ~^ image[22][11] + signed_kernel[4][2] ~^ image[22][12] + signed_kernel[4][3] ~^ image[22][13] + signed_kernel[4][4] ~^ image[22][14];
assign xor_sum[18][11] = signed_kernel[0][0] ~^ image[18][11] + signed_kernel[0][1] ~^ image[18][12] + signed_kernel[0][2] ~^ image[18][13] + signed_kernel[0][3] ~^ image[18][14] + signed_kernel[0][4] ~^ image[18][15] + signed_kernel[1][0] ~^ image[19][11] + signed_kernel[1][1] ~^ image[19][12] + signed_kernel[1][2] ~^ image[19][13] + signed_kernel[1][3] ~^ image[19][14] + signed_kernel[1][4] ~^ image[19][15] + signed_kernel[2][0] ~^ image[20][11] + signed_kernel[2][1] ~^ image[20][12] + signed_kernel[2][2] ~^ image[20][13] + signed_kernel[2][3] ~^ image[20][14] + signed_kernel[2][4] ~^ image[20][15] + signed_kernel[3][0] ~^ image[21][11] + signed_kernel[3][1] ~^ image[21][12] + signed_kernel[3][2] ~^ image[21][13] + signed_kernel[3][3] ~^ image[21][14] + signed_kernel[3][4] ~^ image[21][15] + signed_kernel[4][0] ~^ image[22][11] + signed_kernel[4][1] ~^ image[22][12] + signed_kernel[4][2] ~^ image[22][13] + signed_kernel[4][3] ~^ image[22][14] + signed_kernel[4][4] ~^ image[22][15];
assign xor_sum[18][12] = signed_kernel[0][0] ~^ image[18][12] + signed_kernel[0][1] ~^ image[18][13] + signed_kernel[0][2] ~^ image[18][14] + signed_kernel[0][3] ~^ image[18][15] + signed_kernel[0][4] ~^ image[18][16] + signed_kernel[1][0] ~^ image[19][12] + signed_kernel[1][1] ~^ image[19][13] + signed_kernel[1][2] ~^ image[19][14] + signed_kernel[1][3] ~^ image[19][15] + signed_kernel[1][4] ~^ image[19][16] + signed_kernel[2][0] ~^ image[20][12] + signed_kernel[2][1] ~^ image[20][13] + signed_kernel[2][2] ~^ image[20][14] + signed_kernel[2][3] ~^ image[20][15] + signed_kernel[2][4] ~^ image[20][16] + signed_kernel[3][0] ~^ image[21][12] + signed_kernel[3][1] ~^ image[21][13] + signed_kernel[3][2] ~^ image[21][14] + signed_kernel[3][3] ~^ image[21][15] + signed_kernel[3][4] ~^ image[21][16] + signed_kernel[4][0] ~^ image[22][12] + signed_kernel[4][1] ~^ image[22][13] + signed_kernel[4][2] ~^ image[22][14] + signed_kernel[4][3] ~^ image[22][15] + signed_kernel[4][4] ~^ image[22][16];
assign xor_sum[18][13] = signed_kernel[0][0] ~^ image[18][13] + signed_kernel[0][1] ~^ image[18][14] + signed_kernel[0][2] ~^ image[18][15] + signed_kernel[0][3] ~^ image[18][16] + signed_kernel[0][4] ~^ image[18][17] + signed_kernel[1][0] ~^ image[19][13] + signed_kernel[1][1] ~^ image[19][14] + signed_kernel[1][2] ~^ image[19][15] + signed_kernel[1][3] ~^ image[19][16] + signed_kernel[1][4] ~^ image[19][17] + signed_kernel[2][0] ~^ image[20][13] + signed_kernel[2][1] ~^ image[20][14] + signed_kernel[2][2] ~^ image[20][15] + signed_kernel[2][3] ~^ image[20][16] + signed_kernel[2][4] ~^ image[20][17] + signed_kernel[3][0] ~^ image[21][13] + signed_kernel[3][1] ~^ image[21][14] + signed_kernel[3][2] ~^ image[21][15] + signed_kernel[3][3] ~^ image[21][16] + signed_kernel[3][4] ~^ image[21][17] + signed_kernel[4][0] ~^ image[22][13] + signed_kernel[4][1] ~^ image[22][14] + signed_kernel[4][2] ~^ image[22][15] + signed_kernel[4][3] ~^ image[22][16] + signed_kernel[4][4] ~^ image[22][17];
assign xor_sum[18][14] = signed_kernel[0][0] ~^ image[18][14] + signed_kernel[0][1] ~^ image[18][15] + signed_kernel[0][2] ~^ image[18][16] + signed_kernel[0][3] ~^ image[18][17] + signed_kernel[0][4] ~^ image[18][18] + signed_kernel[1][0] ~^ image[19][14] + signed_kernel[1][1] ~^ image[19][15] + signed_kernel[1][2] ~^ image[19][16] + signed_kernel[1][3] ~^ image[19][17] + signed_kernel[1][4] ~^ image[19][18] + signed_kernel[2][0] ~^ image[20][14] + signed_kernel[2][1] ~^ image[20][15] + signed_kernel[2][2] ~^ image[20][16] + signed_kernel[2][3] ~^ image[20][17] + signed_kernel[2][4] ~^ image[20][18] + signed_kernel[3][0] ~^ image[21][14] + signed_kernel[3][1] ~^ image[21][15] + signed_kernel[3][2] ~^ image[21][16] + signed_kernel[3][3] ~^ image[21][17] + signed_kernel[3][4] ~^ image[21][18] + signed_kernel[4][0] ~^ image[22][14] + signed_kernel[4][1] ~^ image[22][15] + signed_kernel[4][2] ~^ image[22][16] + signed_kernel[4][3] ~^ image[22][17] + signed_kernel[4][4] ~^ image[22][18];
assign xor_sum[18][15] = signed_kernel[0][0] ~^ image[18][15] + signed_kernel[0][1] ~^ image[18][16] + signed_kernel[0][2] ~^ image[18][17] + signed_kernel[0][3] ~^ image[18][18] + signed_kernel[0][4] ~^ image[18][19] + signed_kernel[1][0] ~^ image[19][15] + signed_kernel[1][1] ~^ image[19][16] + signed_kernel[1][2] ~^ image[19][17] + signed_kernel[1][3] ~^ image[19][18] + signed_kernel[1][4] ~^ image[19][19] + signed_kernel[2][0] ~^ image[20][15] + signed_kernel[2][1] ~^ image[20][16] + signed_kernel[2][2] ~^ image[20][17] + signed_kernel[2][3] ~^ image[20][18] + signed_kernel[2][4] ~^ image[20][19] + signed_kernel[3][0] ~^ image[21][15] + signed_kernel[3][1] ~^ image[21][16] + signed_kernel[3][2] ~^ image[21][17] + signed_kernel[3][3] ~^ image[21][18] + signed_kernel[3][4] ~^ image[21][19] + signed_kernel[4][0] ~^ image[22][15] + signed_kernel[4][1] ~^ image[22][16] + signed_kernel[4][2] ~^ image[22][17] + signed_kernel[4][3] ~^ image[22][18] + signed_kernel[4][4] ~^ image[22][19];
assign xor_sum[18][16] = signed_kernel[0][0] ~^ image[18][16] + signed_kernel[0][1] ~^ image[18][17] + signed_kernel[0][2] ~^ image[18][18] + signed_kernel[0][3] ~^ image[18][19] + signed_kernel[0][4] ~^ image[18][20] + signed_kernel[1][0] ~^ image[19][16] + signed_kernel[1][1] ~^ image[19][17] + signed_kernel[1][2] ~^ image[19][18] + signed_kernel[1][3] ~^ image[19][19] + signed_kernel[1][4] ~^ image[19][20] + signed_kernel[2][0] ~^ image[20][16] + signed_kernel[2][1] ~^ image[20][17] + signed_kernel[2][2] ~^ image[20][18] + signed_kernel[2][3] ~^ image[20][19] + signed_kernel[2][4] ~^ image[20][20] + signed_kernel[3][0] ~^ image[21][16] + signed_kernel[3][1] ~^ image[21][17] + signed_kernel[3][2] ~^ image[21][18] + signed_kernel[3][3] ~^ image[21][19] + signed_kernel[3][4] ~^ image[21][20] + signed_kernel[4][0] ~^ image[22][16] + signed_kernel[4][1] ~^ image[22][17] + signed_kernel[4][2] ~^ image[22][18] + signed_kernel[4][3] ~^ image[22][19] + signed_kernel[4][4] ~^ image[22][20];
assign xor_sum[18][17] = signed_kernel[0][0] ~^ image[18][17] + signed_kernel[0][1] ~^ image[18][18] + signed_kernel[0][2] ~^ image[18][19] + signed_kernel[0][3] ~^ image[18][20] + signed_kernel[0][4] ~^ image[18][21] + signed_kernel[1][0] ~^ image[19][17] + signed_kernel[1][1] ~^ image[19][18] + signed_kernel[1][2] ~^ image[19][19] + signed_kernel[1][3] ~^ image[19][20] + signed_kernel[1][4] ~^ image[19][21] + signed_kernel[2][0] ~^ image[20][17] + signed_kernel[2][1] ~^ image[20][18] + signed_kernel[2][2] ~^ image[20][19] + signed_kernel[2][3] ~^ image[20][20] + signed_kernel[2][4] ~^ image[20][21] + signed_kernel[3][0] ~^ image[21][17] + signed_kernel[3][1] ~^ image[21][18] + signed_kernel[3][2] ~^ image[21][19] + signed_kernel[3][3] ~^ image[21][20] + signed_kernel[3][4] ~^ image[21][21] + signed_kernel[4][0] ~^ image[22][17] + signed_kernel[4][1] ~^ image[22][18] + signed_kernel[4][2] ~^ image[22][19] + signed_kernel[4][3] ~^ image[22][20] + signed_kernel[4][4] ~^ image[22][21];
assign xor_sum[18][18] = signed_kernel[0][0] ~^ image[18][18] + signed_kernel[0][1] ~^ image[18][19] + signed_kernel[0][2] ~^ image[18][20] + signed_kernel[0][3] ~^ image[18][21] + signed_kernel[0][4] ~^ image[18][22] + signed_kernel[1][0] ~^ image[19][18] + signed_kernel[1][1] ~^ image[19][19] + signed_kernel[1][2] ~^ image[19][20] + signed_kernel[1][3] ~^ image[19][21] + signed_kernel[1][4] ~^ image[19][22] + signed_kernel[2][0] ~^ image[20][18] + signed_kernel[2][1] ~^ image[20][19] + signed_kernel[2][2] ~^ image[20][20] + signed_kernel[2][3] ~^ image[20][21] + signed_kernel[2][4] ~^ image[20][22] + signed_kernel[3][0] ~^ image[21][18] + signed_kernel[3][1] ~^ image[21][19] + signed_kernel[3][2] ~^ image[21][20] + signed_kernel[3][3] ~^ image[21][21] + signed_kernel[3][4] ~^ image[21][22] + signed_kernel[4][0] ~^ image[22][18] + signed_kernel[4][1] ~^ image[22][19] + signed_kernel[4][2] ~^ image[22][20] + signed_kernel[4][3] ~^ image[22][21] + signed_kernel[4][4] ~^ image[22][22];
assign xor_sum[18][19] = signed_kernel[0][0] ~^ image[18][19] + signed_kernel[0][1] ~^ image[18][20] + signed_kernel[0][2] ~^ image[18][21] + signed_kernel[0][3] ~^ image[18][22] + signed_kernel[0][4] ~^ image[18][23] + signed_kernel[1][0] ~^ image[19][19] + signed_kernel[1][1] ~^ image[19][20] + signed_kernel[1][2] ~^ image[19][21] + signed_kernel[1][3] ~^ image[19][22] + signed_kernel[1][4] ~^ image[19][23] + signed_kernel[2][0] ~^ image[20][19] + signed_kernel[2][1] ~^ image[20][20] + signed_kernel[2][2] ~^ image[20][21] + signed_kernel[2][3] ~^ image[20][22] + signed_kernel[2][4] ~^ image[20][23] + signed_kernel[3][0] ~^ image[21][19] + signed_kernel[3][1] ~^ image[21][20] + signed_kernel[3][2] ~^ image[21][21] + signed_kernel[3][3] ~^ image[21][22] + signed_kernel[3][4] ~^ image[21][23] + signed_kernel[4][0] ~^ image[22][19] + signed_kernel[4][1] ~^ image[22][20] + signed_kernel[4][2] ~^ image[22][21] + signed_kernel[4][3] ~^ image[22][22] + signed_kernel[4][4] ~^ image[22][23];
assign xor_sum[18][20] = signed_kernel[0][0] ~^ image[18][20] + signed_kernel[0][1] ~^ image[18][21] + signed_kernel[0][2] ~^ image[18][22] + signed_kernel[0][3] ~^ image[18][23] + signed_kernel[0][4] ~^ image[18][24] + signed_kernel[1][0] ~^ image[19][20] + signed_kernel[1][1] ~^ image[19][21] + signed_kernel[1][2] ~^ image[19][22] + signed_kernel[1][3] ~^ image[19][23] + signed_kernel[1][4] ~^ image[19][24] + signed_kernel[2][0] ~^ image[20][20] + signed_kernel[2][1] ~^ image[20][21] + signed_kernel[2][2] ~^ image[20][22] + signed_kernel[2][3] ~^ image[20][23] + signed_kernel[2][4] ~^ image[20][24] + signed_kernel[3][0] ~^ image[21][20] + signed_kernel[3][1] ~^ image[21][21] + signed_kernel[3][2] ~^ image[21][22] + signed_kernel[3][3] ~^ image[21][23] + signed_kernel[3][4] ~^ image[21][24] + signed_kernel[4][0] ~^ image[22][20] + signed_kernel[4][1] ~^ image[22][21] + signed_kernel[4][2] ~^ image[22][22] + signed_kernel[4][3] ~^ image[22][23] + signed_kernel[4][4] ~^ image[22][24];
assign xor_sum[18][21] = signed_kernel[0][0] ~^ image[18][21] + signed_kernel[0][1] ~^ image[18][22] + signed_kernel[0][2] ~^ image[18][23] + signed_kernel[0][3] ~^ image[18][24] + signed_kernel[0][4] ~^ image[18][25] + signed_kernel[1][0] ~^ image[19][21] + signed_kernel[1][1] ~^ image[19][22] + signed_kernel[1][2] ~^ image[19][23] + signed_kernel[1][3] ~^ image[19][24] + signed_kernel[1][4] ~^ image[19][25] + signed_kernel[2][0] ~^ image[20][21] + signed_kernel[2][1] ~^ image[20][22] + signed_kernel[2][2] ~^ image[20][23] + signed_kernel[2][3] ~^ image[20][24] + signed_kernel[2][4] ~^ image[20][25] + signed_kernel[3][0] ~^ image[21][21] + signed_kernel[3][1] ~^ image[21][22] + signed_kernel[3][2] ~^ image[21][23] + signed_kernel[3][3] ~^ image[21][24] + signed_kernel[3][4] ~^ image[21][25] + signed_kernel[4][0] ~^ image[22][21] + signed_kernel[4][1] ~^ image[22][22] + signed_kernel[4][2] ~^ image[22][23] + signed_kernel[4][3] ~^ image[22][24] + signed_kernel[4][4] ~^ image[22][25];
assign xor_sum[18][22] = signed_kernel[0][0] ~^ image[18][22] + signed_kernel[0][1] ~^ image[18][23] + signed_kernel[0][2] ~^ image[18][24] + signed_kernel[0][3] ~^ image[18][25] + signed_kernel[0][4] ~^ image[18][26] + signed_kernel[1][0] ~^ image[19][22] + signed_kernel[1][1] ~^ image[19][23] + signed_kernel[1][2] ~^ image[19][24] + signed_kernel[1][3] ~^ image[19][25] + signed_kernel[1][4] ~^ image[19][26] + signed_kernel[2][0] ~^ image[20][22] + signed_kernel[2][1] ~^ image[20][23] + signed_kernel[2][2] ~^ image[20][24] + signed_kernel[2][3] ~^ image[20][25] + signed_kernel[2][4] ~^ image[20][26] + signed_kernel[3][0] ~^ image[21][22] + signed_kernel[3][1] ~^ image[21][23] + signed_kernel[3][2] ~^ image[21][24] + signed_kernel[3][3] ~^ image[21][25] + signed_kernel[3][4] ~^ image[21][26] + signed_kernel[4][0] ~^ image[22][22] + signed_kernel[4][1] ~^ image[22][23] + signed_kernel[4][2] ~^ image[22][24] + signed_kernel[4][3] ~^ image[22][25] + signed_kernel[4][4] ~^ image[22][26];
assign xor_sum[18][23] = signed_kernel[0][0] ~^ image[18][23] + signed_kernel[0][1] ~^ image[18][24] + signed_kernel[0][2] ~^ image[18][25] + signed_kernel[0][3] ~^ image[18][26] + signed_kernel[0][4] ~^ image[18][27] + signed_kernel[1][0] ~^ image[19][23] + signed_kernel[1][1] ~^ image[19][24] + signed_kernel[1][2] ~^ image[19][25] + signed_kernel[1][3] ~^ image[19][26] + signed_kernel[1][4] ~^ image[19][27] + signed_kernel[2][0] ~^ image[20][23] + signed_kernel[2][1] ~^ image[20][24] + signed_kernel[2][2] ~^ image[20][25] + signed_kernel[2][3] ~^ image[20][26] + signed_kernel[2][4] ~^ image[20][27] + signed_kernel[3][0] ~^ image[21][23] + signed_kernel[3][1] ~^ image[21][24] + signed_kernel[3][2] ~^ image[21][25] + signed_kernel[3][3] ~^ image[21][26] + signed_kernel[3][4] ~^ image[21][27] + signed_kernel[4][0] ~^ image[22][23] + signed_kernel[4][1] ~^ image[22][24] + signed_kernel[4][2] ~^ image[22][25] + signed_kernel[4][3] ~^ image[22][26] + signed_kernel[4][4] ~^ image[22][27];
assign xor_sum[19][0] = signed_kernel[0][0] ~^ image[19][0] + signed_kernel[0][1] ~^ image[19][1] + signed_kernel[0][2] ~^ image[19][2] + signed_kernel[0][3] ~^ image[19][3] + signed_kernel[0][4] ~^ image[19][4] + signed_kernel[1][0] ~^ image[20][0] + signed_kernel[1][1] ~^ image[20][1] + signed_kernel[1][2] ~^ image[20][2] + signed_kernel[1][3] ~^ image[20][3] + signed_kernel[1][4] ~^ image[20][4] + signed_kernel[2][0] ~^ image[21][0] + signed_kernel[2][1] ~^ image[21][1] + signed_kernel[2][2] ~^ image[21][2] + signed_kernel[2][3] ~^ image[21][3] + signed_kernel[2][4] ~^ image[21][4] + signed_kernel[3][0] ~^ image[22][0] + signed_kernel[3][1] ~^ image[22][1] + signed_kernel[3][2] ~^ image[22][2] + signed_kernel[3][3] ~^ image[22][3] + signed_kernel[3][4] ~^ image[22][4] + signed_kernel[4][0] ~^ image[23][0] + signed_kernel[4][1] ~^ image[23][1] + signed_kernel[4][2] ~^ image[23][2] + signed_kernel[4][3] ~^ image[23][3] + signed_kernel[4][4] ~^ image[23][4];
assign xor_sum[19][1] = signed_kernel[0][0] ~^ image[19][1] + signed_kernel[0][1] ~^ image[19][2] + signed_kernel[0][2] ~^ image[19][3] + signed_kernel[0][3] ~^ image[19][4] + signed_kernel[0][4] ~^ image[19][5] + signed_kernel[1][0] ~^ image[20][1] + signed_kernel[1][1] ~^ image[20][2] + signed_kernel[1][2] ~^ image[20][3] + signed_kernel[1][3] ~^ image[20][4] + signed_kernel[1][4] ~^ image[20][5] + signed_kernel[2][0] ~^ image[21][1] + signed_kernel[2][1] ~^ image[21][2] + signed_kernel[2][2] ~^ image[21][3] + signed_kernel[2][3] ~^ image[21][4] + signed_kernel[2][4] ~^ image[21][5] + signed_kernel[3][0] ~^ image[22][1] + signed_kernel[3][1] ~^ image[22][2] + signed_kernel[3][2] ~^ image[22][3] + signed_kernel[3][3] ~^ image[22][4] + signed_kernel[3][4] ~^ image[22][5] + signed_kernel[4][0] ~^ image[23][1] + signed_kernel[4][1] ~^ image[23][2] + signed_kernel[4][2] ~^ image[23][3] + signed_kernel[4][3] ~^ image[23][4] + signed_kernel[4][4] ~^ image[23][5];
assign xor_sum[19][2] = signed_kernel[0][0] ~^ image[19][2] + signed_kernel[0][1] ~^ image[19][3] + signed_kernel[0][2] ~^ image[19][4] + signed_kernel[0][3] ~^ image[19][5] + signed_kernel[0][4] ~^ image[19][6] + signed_kernel[1][0] ~^ image[20][2] + signed_kernel[1][1] ~^ image[20][3] + signed_kernel[1][2] ~^ image[20][4] + signed_kernel[1][3] ~^ image[20][5] + signed_kernel[1][4] ~^ image[20][6] + signed_kernel[2][0] ~^ image[21][2] + signed_kernel[2][1] ~^ image[21][3] + signed_kernel[2][2] ~^ image[21][4] + signed_kernel[2][3] ~^ image[21][5] + signed_kernel[2][4] ~^ image[21][6] + signed_kernel[3][0] ~^ image[22][2] + signed_kernel[3][1] ~^ image[22][3] + signed_kernel[3][2] ~^ image[22][4] + signed_kernel[3][3] ~^ image[22][5] + signed_kernel[3][4] ~^ image[22][6] + signed_kernel[4][0] ~^ image[23][2] + signed_kernel[4][1] ~^ image[23][3] + signed_kernel[4][2] ~^ image[23][4] + signed_kernel[4][3] ~^ image[23][5] + signed_kernel[4][4] ~^ image[23][6];
assign xor_sum[19][3] = signed_kernel[0][0] ~^ image[19][3] + signed_kernel[0][1] ~^ image[19][4] + signed_kernel[0][2] ~^ image[19][5] + signed_kernel[0][3] ~^ image[19][6] + signed_kernel[0][4] ~^ image[19][7] + signed_kernel[1][0] ~^ image[20][3] + signed_kernel[1][1] ~^ image[20][4] + signed_kernel[1][2] ~^ image[20][5] + signed_kernel[1][3] ~^ image[20][6] + signed_kernel[1][4] ~^ image[20][7] + signed_kernel[2][0] ~^ image[21][3] + signed_kernel[2][1] ~^ image[21][4] + signed_kernel[2][2] ~^ image[21][5] + signed_kernel[2][3] ~^ image[21][6] + signed_kernel[2][4] ~^ image[21][7] + signed_kernel[3][0] ~^ image[22][3] + signed_kernel[3][1] ~^ image[22][4] + signed_kernel[3][2] ~^ image[22][5] + signed_kernel[3][3] ~^ image[22][6] + signed_kernel[3][4] ~^ image[22][7] + signed_kernel[4][0] ~^ image[23][3] + signed_kernel[4][1] ~^ image[23][4] + signed_kernel[4][2] ~^ image[23][5] + signed_kernel[4][3] ~^ image[23][6] + signed_kernel[4][4] ~^ image[23][7];
assign xor_sum[19][4] = signed_kernel[0][0] ~^ image[19][4] + signed_kernel[0][1] ~^ image[19][5] + signed_kernel[0][2] ~^ image[19][6] + signed_kernel[0][3] ~^ image[19][7] + signed_kernel[0][4] ~^ image[19][8] + signed_kernel[1][0] ~^ image[20][4] + signed_kernel[1][1] ~^ image[20][5] + signed_kernel[1][2] ~^ image[20][6] + signed_kernel[1][3] ~^ image[20][7] + signed_kernel[1][4] ~^ image[20][8] + signed_kernel[2][0] ~^ image[21][4] + signed_kernel[2][1] ~^ image[21][5] + signed_kernel[2][2] ~^ image[21][6] + signed_kernel[2][3] ~^ image[21][7] + signed_kernel[2][4] ~^ image[21][8] + signed_kernel[3][0] ~^ image[22][4] + signed_kernel[3][1] ~^ image[22][5] + signed_kernel[3][2] ~^ image[22][6] + signed_kernel[3][3] ~^ image[22][7] + signed_kernel[3][4] ~^ image[22][8] + signed_kernel[4][0] ~^ image[23][4] + signed_kernel[4][1] ~^ image[23][5] + signed_kernel[4][2] ~^ image[23][6] + signed_kernel[4][3] ~^ image[23][7] + signed_kernel[4][4] ~^ image[23][8];
assign xor_sum[19][5] = signed_kernel[0][0] ~^ image[19][5] + signed_kernel[0][1] ~^ image[19][6] + signed_kernel[0][2] ~^ image[19][7] + signed_kernel[0][3] ~^ image[19][8] + signed_kernel[0][4] ~^ image[19][9] + signed_kernel[1][0] ~^ image[20][5] + signed_kernel[1][1] ~^ image[20][6] + signed_kernel[1][2] ~^ image[20][7] + signed_kernel[1][3] ~^ image[20][8] + signed_kernel[1][4] ~^ image[20][9] + signed_kernel[2][0] ~^ image[21][5] + signed_kernel[2][1] ~^ image[21][6] + signed_kernel[2][2] ~^ image[21][7] + signed_kernel[2][3] ~^ image[21][8] + signed_kernel[2][4] ~^ image[21][9] + signed_kernel[3][0] ~^ image[22][5] + signed_kernel[3][1] ~^ image[22][6] + signed_kernel[3][2] ~^ image[22][7] + signed_kernel[3][3] ~^ image[22][8] + signed_kernel[3][4] ~^ image[22][9] + signed_kernel[4][0] ~^ image[23][5] + signed_kernel[4][1] ~^ image[23][6] + signed_kernel[4][2] ~^ image[23][7] + signed_kernel[4][3] ~^ image[23][8] + signed_kernel[4][4] ~^ image[23][9];
assign xor_sum[19][6] = signed_kernel[0][0] ~^ image[19][6] + signed_kernel[0][1] ~^ image[19][7] + signed_kernel[0][2] ~^ image[19][8] + signed_kernel[0][3] ~^ image[19][9] + signed_kernel[0][4] ~^ image[19][10] + signed_kernel[1][0] ~^ image[20][6] + signed_kernel[1][1] ~^ image[20][7] + signed_kernel[1][2] ~^ image[20][8] + signed_kernel[1][3] ~^ image[20][9] + signed_kernel[1][4] ~^ image[20][10] + signed_kernel[2][0] ~^ image[21][6] + signed_kernel[2][1] ~^ image[21][7] + signed_kernel[2][2] ~^ image[21][8] + signed_kernel[2][3] ~^ image[21][9] + signed_kernel[2][4] ~^ image[21][10] + signed_kernel[3][0] ~^ image[22][6] + signed_kernel[3][1] ~^ image[22][7] + signed_kernel[3][2] ~^ image[22][8] + signed_kernel[3][3] ~^ image[22][9] + signed_kernel[3][4] ~^ image[22][10] + signed_kernel[4][0] ~^ image[23][6] + signed_kernel[4][1] ~^ image[23][7] + signed_kernel[4][2] ~^ image[23][8] + signed_kernel[4][3] ~^ image[23][9] + signed_kernel[4][4] ~^ image[23][10];
assign xor_sum[19][7] = signed_kernel[0][0] ~^ image[19][7] + signed_kernel[0][1] ~^ image[19][8] + signed_kernel[0][2] ~^ image[19][9] + signed_kernel[0][3] ~^ image[19][10] + signed_kernel[0][4] ~^ image[19][11] + signed_kernel[1][0] ~^ image[20][7] + signed_kernel[1][1] ~^ image[20][8] + signed_kernel[1][2] ~^ image[20][9] + signed_kernel[1][3] ~^ image[20][10] + signed_kernel[1][4] ~^ image[20][11] + signed_kernel[2][0] ~^ image[21][7] + signed_kernel[2][1] ~^ image[21][8] + signed_kernel[2][2] ~^ image[21][9] + signed_kernel[2][3] ~^ image[21][10] + signed_kernel[2][4] ~^ image[21][11] + signed_kernel[3][0] ~^ image[22][7] + signed_kernel[3][1] ~^ image[22][8] + signed_kernel[3][2] ~^ image[22][9] + signed_kernel[3][3] ~^ image[22][10] + signed_kernel[3][4] ~^ image[22][11] + signed_kernel[4][0] ~^ image[23][7] + signed_kernel[4][1] ~^ image[23][8] + signed_kernel[4][2] ~^ image[23][9] + signed_kernel[4][3] ~^ image[23][10] + signed_kernel[4][4] ~^ image[23][11];
assign xor_sum[19][8] = signed_kernel[0][0] ~^ image[19][8] + signed_kernel[0][1] ~^ image[19][9] + signed_kernel[0][2] ~^ image[19][10] + signed_kernel[0][3] ~^ image[19][11] + signed_kernel[0][4] ~^ image[19][12] + signed_kernel[1][0] ~^ image[20][8] + signed_kernel[1][1] ~^ image[20][9] + signed_kernel[1][2] ~^ image[20][10] + signed_kernel[1][3] ~^ image[20][11] + signed_kernel[1][4] ~^ image[20][12] + signed_kernel[2][0] ~^ image[21][8] + signed_kernel[2][1] ~^ image[21][9] + signed_kernel[2][2] ~^ image[21][10] + signed_kernel[2][3] ~^ image[21][11] + signed_kernel[2][4] ~^ image[21][12] + signed_kernel[3][0] ~^ image[22][8] + signed_kernel[3][1] ~^ image[22][9] + signed_kernel[3][2] ~^ image[22][10] + signed_kernel[3][3] ~^ image[22][11] + signed_kernel[3][4] ~^ image[22][12] + signed_kernel[4][0] ~^ image[23][8] + signed_kernel[4][1] ~^ image[23][9] + signed_kernel[4][2] ~^ image[23][10] + signed_kernel[4][3] ~^ image[23][11] + signed_kernel[4][4] ~^ image[23][12];
assign xor_sum[19][9] = signed_kernel[0][0] ~^ image[19][9] + signed_kernel[0][1] ~^ image[19][10] + signed_kernel[0][2] ~^ image[19][11] + signed_kernel[0][3] ~^ image[19][12] + signed_kernel[0][4] ~^ image[19][13] + signed_kernel[1][0] ~^ image[20][9] + signed_kernel[1][1] ~^ image[20][10] + signed_kernel[1][2] ~^ image[20][11] + signed_kernel[1][3] ~^ image[20][12] + signed_kernel[1][4] ~^ image[20][13] + signed_kernel[2][0] ~^ image[21][9] + signed_kernel[2][1] ~^ image[21][10] + signed_kernel[2][2] ~^ image[21][11] + signed_kernel[2][3] ~^ image[21][12] + signed_kernel[2][4] ~^ image[21][13] + signed_kernel[3][0] ~^ image[22][9] + signed_kernel[3][1] ~^ image[22][10] + signed_kernel[3][2] ~^ image[22][11] + signed_kernel[3][3] ~^ image[22][12] + signed_kernel[3][4] ~^ image[22][13] + signed_kernel[4][0] ~^ image[23][9] + signed_kernel[4][1] ~^ image[23][10] + signed_kernel[4][2] ~^ image[23][11] + signed_kernel[4][3] ~^ image[23][12] + signed_kernel[4][4] ~^ image[23][13];
assign xor_sum[19][10] = signed_kernel[0][0] ~^ image[19][10] + signed_kernel[0][1] ~^ image[19][11] + signed_kernel[0][2] ~^ image[19][12] + signed_kernel[0][3] ~^ image[19][13] + signed_kernel[0][4] ~^ image[19][14] + signed_kernel[1][0] ~^ image[20][10] + signed_kernel[1][1] ~^ image[20][11] + signed_kernel[1][2] ~^ image[20][12] + signed_kernel[1][3] ~^ image[20][13] + signed_kernel[1][4] ~^ image[20][14] + signed_kernel[2][0] ~^ image[21][10] + signed_kernel[2][1] ~^ image[21][11] + signed_kernel[2][2] ~^ image[21][12] + signed_kernel[2][3] ~^ image[21][13] + signed_kernel[2][4] ~^ image[21][14] + signed_kernel[3][0] ~^ image[22][10] + signed_kernel[3][1] ~^ image[22][11] + signed_kernel[3][2] ~^ image[22][12] + signed_kernel[3][3] ~^ image[22][13] + signed_kernel[3][4] ~^ image[22][14] + signed_kernel[4][0] ~^ image[23][10] + signed_kernel[4][1] ~^ image[23][11] + signed_kernel[4][2] ~^ image[23][12] + signed_kernel[4][3] ~^ image[23][13] + signed_kernel[4][4] ~^ image[23][14];
assign xor_sum[19][11] = signed_kernel[0][0] ~^ image[19][11] + signed_kernel[0][1] ~^ image[19][12] + signed_kernel[0][2] ~^ image[19][13] + signed_kernel[0][3] ~^ image[19][14] + signed_kernel[0][4] ~^ image[19][15] + signed_kernel[1][0] ~^ image[20][11] + signed_kernel[1][1] ~^ image[20][12] + signed_kernel[1][2] ~^ image[20][13] + signed_kernel[1][3] ~^ image[20][14] + signed_kernel[1][4] ~^ image[20][15] + signed_kernel[2][0] ~^ image[21][11] + signed_kernel[2][1] ~^ image[21][12] + signed_kernel[2][2] ~^ image[21][13] + signed_kernel[2][3] ~^ image[21][14] + signed_kernel[2][4] ~^ image[21][15] + signed_kernel[3][0] ~^ image[22][11] + signed_kernel[3][1] ~^ image[22][12] + signed_kernel[3][2] ~^ image[22][13] + signed_kernel[3][3] ~^ image[22][14] + signed_kernel[3][4] ~^ image[22][15] + signed_kernel[4][0] ~^ image[23][11] + signed_kernel[4][1] ~^ image[23][12] + signed_kernel[4][2] ~^ image[23][13] + signed_kernel[4][3] ~^ image[23][14] + signed_kernel[4][4] ~^ image[23][15];
assign xor_sum[19][12] = signed_kernel[0][0] ~^ image[19][12] + signed_kernel[0][1] ~^ image[19][13] + signed_kernel[0][2] ~^ image[19][14] + signed_kernel[0][3] ~^ image[19][15] + signed_kernel[0][4] ~^ image[19][16] + signed_kernel[1][0] ~^ image[20][12] + signed_kernel[1][1] ~^ image[20][13] + signed_kernel[1][2] ~^ image[20][14] + signed_kernel[1][3] ~^ image[20][15] + signed_kernel[1][4] ~^ image[20][16] + signed_kernel[2][0] ~^ image[21][12] + signed_kernel[2][1] ~^ image[21][13] + signed_kernel[2][2] ~^ image[21][14] + signed_kernel[2][3] ~^ image[21][15] + signed_kernel[2][4] ~^ image[21][16] + signed_kernel[3][0] ~^ image[22][12] + signed_kernel[3][1] ~^ image[22][13] + signed_kernel[3][2] ~^ image[22][14] + signed_kernel[3][3] ~^ image[22][15] + signed_kernel[3][4] ~^ image[22][16] + signed_kernel[4][0] ~^ image[23][12] + signed_kernel[4][1] ~^ image[23][13] + signed_kernel[4][2] ~^ image[23][14] + signed_kernel[4][3] ~^ image[23][15] + signed_kernel[4][4] ~^ image[23][16];
assign xor_sum[19][13] = signed_kernel[0][0] ~^ image[19][13] + signed_kernel[0][1] ~^ image[19][14] + signed_kernel[0][2] ~^ image[19][15] + signed_kernel[0][3] ~^ image[19][16] + signed_kernel[0][4] ~^ image[19][17] + signed_kernel[1][0] ~^ image[20][13] + signed_kernel[1][1] ~^ image[20][14] + signed_kernel[1][2] ~^ image[20][15] + signed_kernel[1][3] ~^ image[20][16] + signed_kernel[1][4] ~^ image[20][17] + signed_kernel[2][0] ~^ image[21][13] + signed_kernel[2][1] ~^ image[21][14] + signed_kernel[2][2] ~^ image[21][15] + signed_kernel[2][3] ~^ image[21][16] + signed_kernel[2][4] ~^ image[21][17] + signed_kernel[3][0] ~^ image[22][13] + signed_kernel[3][1] ~^ image[22][14] + signed_kernel[3][2] ~^ image[22][15] + signed_kernel[3][3] ~^ image[22][16] + signed_kernel[3][4] ~^ image[22][17] + signed_kernel[4][0] ~^ image[23][13] + signed_kernel[4][1] ~^ image[23][14] + signed_kernel[4][2] ~^ image[23][15] + signed_kernel[4][3] ~^ image[23][16] + signed_kernel[4][4] ~^ image[23][17];
assign xor_sum[19][14] = signed_kernel[0][0] ~^ image[19][14] + signed_kernel[0][1] ~^ image[19][15] + signed_kernel[0][2] ~^ image[19][16] + signed_kernel[0][3] ~^ image[19][17] + signed_kernel[0][4] ~^ image[19][18] + signed_kernel[1][0] ~^ image[20][14] + signed_kernel[1][1] ~^ image[20][15] + signed_kernel[1][2] ~^ image[20][16] + signed_kernel[1][3] ~^ image[20][17] + signed_kernel[1][4] ~^ image[20][18] + signed_kernel[2][0] ~^ image[21][14] + signed_kernel[2][1] ~^ image[21][15] + signed_kernel[2][2] ~^ image[21][16] + signed_kernel[2][3] ~^ image[21][17] + signed_kernel[2][4] ~^ image[21][18] + signed_kernel[3][0] ~^ image[22][14] + signed_kernel[3][1] ~^ image[22][15] + signed_kernel[3][2] ~^ image[22][16] + signed_kernel[3][3] ~^ image[22][17] + signed_kernel[3][4] ~^ image[22][18] + signed_kernel[4][0] ~^ image[23][14] + signed_kernel[4][1] ~^ image[23][15] + signed_kernel[4][2] ~^ image[23][16] + signed_kernel[4][3] ~^ image[23][17] + signed_kernel[4][4] ~^ image[23][18];
assign xor_sum[19][15] = signed_kernel[0][0] ~^ image[19][15] + signed_kernel[0][1] ~^ image[19][16] + signed_kernel[0][2] ~^ image[19][17] + signed_kernel[0][3] ~^ image[19][18] + signed_kernel[0][4] ~^ image[19][19] + signed_kernel[1][0] ~^ image[20][15] + signed_kernel[1][1] ~^ image[20][16] + signed_kernel[1][2] ~^ image[20][17] + signed_kernel[1][3] ~^ image[20][18] + signed_kernel[1][4] ~^ image[20][19] + signed_kernel[2][0] ~^ image[21][15] + signed_kernel[2][1] ~^ image[21][16] + signed_kernel[2][2] ~^ image[21][17] + signed_kernel[2][3] ~^ image[21][18] + signed_kernel[2][4] ~^ image[21][19] + signed_kernel[3][0] ~^ image[22][15] + signed_kernel[3][1] ~^ image[22][16] + signed_kernel[3][2] ~^ image[22][17] + signed_kernel[3][3] ~^ image[22][18] + signed_kernel[3][4] ~^ image[22][19] + signed_kernel[4][0] ~^ image[23][15] + signed_kernel[4][1] ~^ image[23][16] + signed_kernel[4][2] ~^ image[23][17] + signed_kernel[4][3] ~^ image[23][18] + signed_kernel[4][4] ~^ image[23][19];
assign xor_sum[19][16] = signed_kernel[0][0] ~^ image[19][16] + signed_kernel[0][1] ~^ image[19][17] + signed_kernel[0][2] ~^ image[19][18] + signed_kernel[0][3] ~^ image[19][19] + signed_kernel[0][4] ~^ image[19][20] + signed_kernel[1][0] ~^ image[20][16] + signed_kernel[1][1] ~^ image[20][17] + signed_kernel[1][2] ~^ image[20][18] + signed_kernel[1][3] ~^ image[20][19] + signed_kernel[1][4] ~^ image[20][20] + signed_kernel[2][0] ~^ image[21][16] + signed_kernel[2][1] ~^ image[21][17] + signed_kernel[2][2] ~^ image[21][18] + signed_kernel[2][3] ~^ image[21][19] + signed_kernel[2][4] ~^ image[21][20] + signed_kernel[3][0] ~^ image[22][16] + signed_kernel[3][1] ~^ image[22][17] + signed_kernel[3][2] ~^ image[22][18] + signed_kernel[3][3] ~^ image[22][19] + signed_kernel[3][4] ~^ image[22][20] + signed_kernel[4][0] ~^ image[23][16] + signed_kernel[4][1] ~^ image[23][17] + signed_kernel[4][2] ~^ image[23][18] + signed_kernel[4][3] ~^ image[23][19] + signed_kernel[4][4] ~^ image[23][20];
assign xor_sum[19][17] = signed_kernel[0][0] ~^ image[19][17] + signed_kernel[0][1] ~^ image[19][18] + signed_kernel[0][2] ~^ image[19][19] + signed_kernel[0][3] ~^ image[19][20] + signed_kernel[0][4] ~^ image[19][21] + signed_kernel[1][0] ~^ image[20][17] + signed_kernel[1][1] ~^ image[20][18] + signed_kernel[1][2] ~^ image[20][19] + signed_kernel[1][3] ~^ image[20][20] + signed_kernel[1][4] ~^ image[20][21] + signed_kernel[2][0] ~^ image[21][17] + signed_kernel[2][1] ~^ image[21][18] + signed_kernel[2][2] ~^ image[21][19] + signed_kernel[2][3] ~^ image[21][20] + signed_kernel[2][4] ~^ image[21][21] + signed_kernel[3][0] ~^ image[22][17] + signed_kernel[3][1] ~^ image[22][18] + signed_kernel[3][2] ~^ image[22][19] + signed_kernel[3][3] ~^ image[22][20] + signed_kernel[3][4] ~^ image[22][21] + signed_kernel[4][0] ~^ image[23][17] + signed_kernel[4][1] ~^ image[23][18] + signed_kernel[4][2] ~^ image[23][19] + signed_kernel[4][3] ~^ image[23][20] + signed_kernel[4][4] ~^ image[23][21];
assign xor_sum[19][18] = signed_kernel[0][0] ~^ image[19][18] + signed_kernel[0][1] ~^ image[19][19] + signed_kernel[0][2] ~^ image[19][20] + signed_kernel[0][3] ~^ image[19][21] + signed_kernel[0][4] ~^ image[19][22] + signed_kernel[1][0] ~^ image[20][18] + signed_kernel[1][1] ~^ image[20][19] + signed_kernel[1][2] ~^ image[20][20] + signed_kernel[1][3] ~^ image[20][21] + signed_kernel[1][4] ~^ image[20][22] + signed_kernel[2][0] ~^ image[21][18] + signed_kernel[2][1] ~^ image[21][19] + signed_kernel[2][2] ~^ image[21][20] + signed_kernel[2][3] ~^ image[21][21] + signed_kernel[2][4] ~^ image[21][22] + signed_kernel[3][0] ~^ image[22][18] + signed_kernel[3][1] ~^ image[22][19] + signed_kernel[3][2] ~^ image[22][20] + signed_kernel[3][3] ~^ image[22][21] + signed_kernel[3][4] ~^ image[22][22] + signed_kernel[4][0] ~^ image[23][18] + signed_kernel[4][1] ~^ image[23][19] + signed_kernel[4][2] ~^ image[23][20] + signed_kernel[4][3] ~^ image[23][21] + signed_kernel[4][4] ~^ image[23][22];
assign xor_sum[19][19] = signed_kernel[0][0] ~^ image[19][19] + signed_kernel[0][1] ~^ image[19][20] + signed_kernel[0][2] ~^ image[19][21] + signed_kernel[0][3] ~^ image[19][22] + signed_kernel[0][4] ~^ image[19][23] + signed_kernel[1][0] ~^ image[20][19] + signed_kernel[1][1] ~^ image[20][20] + signed_kernel[1][2] ~^ image[20][21] + signed_kernel[1][3] ~^ image[20][22] + signed_kernel[1][4] ~^ image[20][23] + signed_kernel[2][0] ~^ image[21][19] + signed_kernel[2][1] ~^ image[21][20] + signed_kernel[2][2] ~^ image[21][21] + signed_kernel[2][3] ~^ image[21][22] + signed_kernel[2][4] ~^ image[21][23] + signed_kernel[3][0] ~^ image[22][19] + signed_kernel[3][1] ~^ image[22][20] + signed_kernel[3][2] ~^ image[22][21] + signed_kernel[3][3] ~^ image[22][22] + signed_kernel[3][4] ~^ image[22][23] + signed_kernel[4][0] ~^ image[23][19] + signed_kernel[4][1] ~^ image[23][20] + signed_kernel[4][2] ~^ image[23][21] + signed_kernel[4][3] ~^ image[23][22] + signed_kernel[4][4] ~^ image[23][23];
assign xor_sum[19][20] = signed_kernel[0][0] ~^ image[19][20] + signed_kernel[0][1] ~^ image[19][21] + signed_kernel[0][2] ~^ image[19][22] + signed_kernel[0][3] ~^ image[19][23] + signed_kernel[0][4] ~^ image[19][24] + signed_kernel[1][0] ~^ image[20][20] + signed_kernel[1][1] ~^ image[20][21] + signed_kernel[1][2] ~^ image[20][22] + signed_kernel[1][3] ~^ image[20][23] + signed_kernel[1][4] ~^ image[20][24] + signed_kernel[2][0] ~^ image[21][20] + signed_kernel[2][1] ~^ image[21][21] + signed_kernel[2][2] ~^ image[21][22] + signed_kernel[2][3] ~^ image[21][23] + signed_kernel[2][4] ~^ image[21][24] + signed_kernel[3][0] ~^ image[22][20] + signed_kernel[3][1] ~^ image[22][21] + signed_kernel[3][2] ~^ image[22][22] + signed_kernel[3][3] ~^ image[22][23] + signed_kernel[3][4] ~^ image[22][24] + signed_kernel[4][0] ~^ image[23][20] + signed_kernel[4][1] ~^ image[23][21] + signed_kernel[4][2] ~^ image[23][22] + signed_kernel[4][3] ~^ image[23][23] + signed_kernel[4][4] ~^ image[23][24];
assign xor_sum[19][21] = signed_kernel[0][0] ~^ image[19][21] + signed_kernel[0][1] ~^ image[19][22] + signed_kernel[0][2] ~^ image[19][23] + signed_kernel[0][3] ~^ image[19][24] + signed_kernel[0][4] ~^ image[19][25] + signed_kernel[1][0] ~^ image[20][21] + signed_kernel[1][1] ~^ image[20][22] + signed_kernel[1][2] ~^ image[20][23] + signed_kernel[1][3] ~^ image[20][24] + signed_kernel[1][4] ~^ image[20][25] + signed_kernel[2][0] ~^ image[21][21] + signed_kernel[2][1] ~^ image[21][22] + signed_kernel[2][2] ~^ image[21][23] + signed_kernel[2][3] ~^ image[21][24] + signed_kernel[2][4] ~^ image[21][25] + signed_kernel[3][0] ~^ image[22][21] + signed_kernel[3][1] ~^ image[22][22] + signed_kernel[3][2] ~^ image[22][23] + signed_kernel[3][3] ~^ image[22][24] + signed_kernel[3][4] ~^ image[22][25] + signed_kernel[4][0] ~^ image[23][21] + signed_kernel[4][1] ~^ image[23][22] + signed_kernel[4][2] ~^ image[23][23] + signed_kernel[4][3] ~^ image[23][24] + signed_kernel[4][4] ~^ image[23][25];
assign xor_sum[19][22] = signed_kernel[0][0] ~^ image[19][22] + signed_kernel[0][1] ~^ image[19][23] + signed_kernel[0][2] ~^ image[19][24] + signed_kernel[0][3] ~^ image[19][25] + signed_kernel[0][4] ~^ image[19][26] + signed_kernel[1][0] ~^ image[20][22] + signed_kernel[1][1] ~^ image[20][23] + signed_kernel[1][2] ~^ image[20][24] + signed_kernel[1][3] ~^ image[20][25] + signed_kernel[1][4] ~^ image[20][26] + signed_kernel[2][0] ~^ image[21][22] + signed_kernel[2][1] ~^ image[21][23] + signed_kernel[2][2] ~^ image[21][24] + signed_kernel[2][3] ~^ image[21][25] + signed_kernel[2][4] ~^ image[21][26] + signed_kernel[3][0] ~^ image[22][22] + signed_kernel[3][1] ~^ image[22][23] + signed_kernel[3][2] ~^ image[22][24] + signed_kernel[3][3] ~^ image[22][25] + signed_kernel[3][4] ~^ image[22][26] + signed_kernel[4][0] ~^ image[23][22] + signed_kernel[4][1] ~^ image[23][23] + signed_kernel[4][2] ~^ image[23][24] + signed_kernel[4][3] ~^ image[23][25] + signed_kernel[4][4] ~^ image[23][26];
assign xor_sum[19][23] = signed_kernel[0][0] ~^ image[19][23] + signed_kernel[0][1] ~^ image[19][24] + signed_kernel[0][2] ~^ image[19][25] + signed_kernel[0][3] ~^ image[19][26] + signed_kernel[0][4] ~^ image[19][27] + signed_kernel[1][0] ~^ image[20][23] + signed_kernel[1][1] ~^ image[20][24] + signed_kernel[1][2] ~^ image[20][25] + signed_kernel[1][3] ~^ image[20][26] + signed_kernel[1][4] ~^ image[20][27] + signed_kernel[2][0] ~^ image[21][23] + signed_kernel[2][1] ~^ image[21][24] + signed_kernel[2][2] ~^ image[21][25] + signed_kernel[2][3] ~^ image[21][26] + signed_kernel[2][4] ~^ image[21][27] + signed_kernel[3][0] ~^ image[22][23] + signed_kernel[3][1] ~^ image[22][24] + signed_kernel[3][2] ~^ image[22][25] + signed_kernel[3][3] ~^ image[22][26] + signed_kernel[3][4] ~^ image[22][27] + signed_kernel[4][0] ~^ image[23][23] + signed_kernel[4][1] ~^ image[23][24] + signed_kernel[4][2] ~^ image[23][25] + signed_kernel[4][3] ~^ image[23][26] + signed_kernel[4][4] ~^ image[23][27];
assign xor_sum[20][0] = signed_kernel[0][0] ~^ image[20][0] + signed_kernel[0][1] ~^ image[20][1] + signed_kernel[0][2] ~^ image[20][2] + signed_kernel[0][3] ~^ image[20][3] + signed_kernel[0][4] ~^ image[20][4] + signed_kernel[1][0] ~^ image[21][0] + signed_kernel[1][1] ~^ image[21][1] + signed_kernel[1][2] ~^ image[21][2] + signed_kernel[1][3] ~^ image[21][3] + signed_kernel[1][4] ~^ image[21][4] + signed_kernel[2][0] ~^ image[22][0] + signed_kernel[2][1] ~^ image[22][1] + signed_kernel[2][2] ~^ image[22][2] + signed_kernel[2][3] ~^ image[22][3] + signed_kernel[2][4] ~^ image[22][4] + signed_kernel[3][0] ~^ image[23][0] + signed_kernel[3][1] ~^ image[23][1] + signed_kernel[3][2] ~^ image[23][2] + signed_kernel[3][3] ~^ image[23][3] + signed_kernel[3][4] ~^ image[23][4] + signed_kernel[4][0] ~^ image[24][0] + signed_kernel[4][1] ~^ image[24][1] + signed_kernel[4][2] ~^ image[24][2] + signed_kernel[4][3] ~^ image[24][3] + signed_kernel[4][4] ~^ image[24][4];
assign xor_sum[20][1] = signed_kernel[0][0] ~^ image[20][1] + signed_kernel[0][1] ~^ image[20][2] + signed_kernel[0][2] ~^ image[20][3] + signed_kernel[0][3] ~^ image[20][4] + signed_kernel[0][4] ~^ image[20][5] + signed_kernel[1][0] ~^ image[21][1] + signed_kernel[1][1] ~^ image[21][2] + signed_kernel[1][2] ~^ image[21][3] + signed_kernel[1][3] ~^ image[21][4] + signed_kernel[1][4] ~^ image[21][5] + signed_kernel[2][0] ~^ image[22][1] + signed_kernel[2][1] ~^ image[22][2] + signed_kernel[2][2] ~^ image[22][3] + signed_kernel[2][3] ~^ image[22][4] + signed_kernel[2][4] ~^ image[22][5] + signed_kernel[3][0] ~^ image[23][1] + signed_kernel[3][1] ~^ image[23][2] + signed_kernel[3][2] ~^ image[23][3] + signed_kernel[3][3] ~^ image[23][4] + signed_kernel[3][4] ~^ image[23][5] + signed_kernel[4][0] ~^ image[24][1] + signed_kernel[4][1] ~^ image[24][2] + signed_kernel[4][2] ~^ image[24][3] + signed_kernel[4][3] ~^ image[24][4] + signed_kernel[4][4] ~^ image[24][5];
assign xor_sum[20][2] = signed_kernel[0][0] ~^ image[20][2] + signed_kernel[0][1] ~^ image[20][3] + signed_kernel[0][2] ~^ image[20][4] + signed_kernel[0][3] ~^ image[20][5] + signed_kernel[0][4] ~^ image[20][6] + signed_kernel[1][0] ~^ image[21][2] + signed_kernel[1][1] ~^ image[21][3] + signed_kernel[1][2] ~^ image[21][4] + signed_kernel[1][3] ~^ image[21][5] + signed_kernel[1][4] ~^ image[21][6] + signed_kernel[2][0] ~^ image[22][2] + signed_kernel[2][1] ~^ image[22][3] + signed_kernel[2][2] ~^ image[22][4] + signed_kernel[2][3] ~^ image[22][5] + signed_kernel[2][4] ~^ image[22][6] + signed_kernel[3][0] ~^ image[23][2] + signed_kernel[3][1] ~^ image[23][3] + signed_kernel[3][2] ~^ image[23][4] + signed_kernel[3][3] ~^ image[23][5] + signed_kernel[3][4] ~^ image[23][6] + signed_kernel[4][0] ~^ image[24][2] + signed_kernel[4][1] ~^ image[24][3] + signed_kernel[4][2] ~^ image[24][4] + signed_kernel[4][3] ~^ image[24][5] + signed_kernel[4][4] ~^ image[24][6];
assign xor_sum[20][3] = signed_kernel[0][0] ~^ image[20][3] + signed_kernel[0][1] ~^ image[20][4] + signed_kernel[0][2] ~^ image[20][5] + signed_kernel[0][3] ~^ image[20][6] + signed_kernel[0][4] ~^ image[20][7] + signed_kernel[1][0] ~^ image[21][3] + signed_kernel[1][1] ~^ image[21][4] + signed_kernel[1][2] ~^ image[21][5] + signed_kernel[1][3] ~^ image[21][6] + signed_kernel[1][4] ~^ image[21][7] + signed_kernel[2][0] ~^ image[22][3] + signed_kernel[2][1] ~^ image[22][4] + signed_kernel[2][2] ~^ image[22][5] + signed_kernel[2][3] ~^ image[22][6] + signed_kernel[2][4] ~^ image[22][7] + signed_kernel[3][0] ~^ image[23][3] + signed_kernel[3][1] ~^ image[23][4] + signed_kernel[3][2] ~^ image[23][5] + signed_kernel[3][3] ~^ image[23][6] + signed_kernel[3][4] ~^ image[23][7] + signed_kernel[4][0] ~^ image[24][3] + signed_kernel[4][1] ~^ image[24][4] + signed_kernel[4][2] ~^ image[24][5] + signed_kernel[4][3] ~^ image[24][6] + signed_kernel[4][4] ~^ image[24][7];
assign xor_sum[20][4] = signed_kernel[0][0] ~^ image[20][4] + signed_kernel[0][1] ~^ image[20][5] + signed_kernel[0][2] ~^ image[20][6] + signed_kernel[0][3] ~^ image[20][7] + signed_kernel[0][4] ~^ image[20][8] + signed_kernel[1][0] ~^ image[21][4] + signed_kernel[1][1] ~^ image[21][5] + signed_kernel[1][2] ~^ image[21][6] + signed_kernel[1][3] ~^ image[21][7] + signed_kernel[1][4] ~^ image[21][8] + signed_kernel[2][0] ~^ image[22][4] + signed_kernel[2][1] ~^ image[22][5] + signed_kernel[2][2] ~^ image[22][6] + signed_kernel[2][3] ~^ image[22][7] + signed_kernel[2][4] ~^ image[22][8] + signed_kernel[3][0] ~^ image[23][4] + signed_kernel[3][1] ~^ image[23][5] + signed_kernel[3][2] ~^ image[23][6] + signed_kernel[3][3] ~^ image[23][7] + signed_kernel[3][4] ~^ image[23][8] + signed_kernel[4][0] ~^ image[24][4] + signed_kernel[4][1] ~^ image[24][5] + signed_kernel[4][2] ~^ image[24][6] + signed_kernel[4][3] ~^ image[24][7] + signed_kernel[4][4] ~^ image[24][8];
assign xor_sum[20][5] = signed_kernel[0][0] ~^ image[20][5] + signed_kernel[0][1] ~^ image[20][6] + signed_kernel[0][2] ~^ image[20][7] + signed_kernel[0][3] ~^ image[20][8] + signed_kernel[0][4] ~^ image[20][9] + signed_kernel[1][0] ~^ image[21][5] + signed_kernel[1][1] ~^ image[21][6] + signed_kernel[1][2] ~^ image[21][7] + signed_kernel[1][3] ~^ image[21][8] + signed_kernel[1][4] ~^ image[21][9] + signed_kernel[2][0] ~^ image[22][5] + signed_kernel[2][1] ~^ image[22][6] + signed_kernel[2][2] ~^ image[22][7] + signed_kernel[2][3] ~^ image[22][8] + signed_kernel[2][4] ~^ image[22][9] + signed_kernel[3][0] ~^ image[23][5] + signed_kernel[3][1] ~^ image[23][6] + signed_kernel[3][2] ~^ image[23][7] + signed_kernel[3][3] ~^ image[23][8] + signed_kernel[3][4] ~^ image[23][9] + signed_kernel[4][0] ~^ image[24][5] + signed_kernel[4][1] ~^ image[24][6] + signed_kernel[4][2] ~^ image[24][7] + signed_kernel[4][3] ~^ image[24][8] + signed_kernel[4][4] ~^ image[24][9];
assign xor_sum[20][6] = signed_kernel[0][0] ~^ image[20][6] + signed_kernel[0][1] ~^ image[20][7] + signed_kernel[0][2] ~^ image[20][8] + signed_kernel[0][3] ~^ image[20][9] + signed_kernel[0][4] ~^ image[20][10] + signed_kernel[1][0] ~^ image[21][6] + signed_kernel[1][1] ~^ image[21][7] + signed_kernel[1][2] ~^ image[21][8] + signed_kernel[1][3] ~^ image[21][9] + signed_kernel[1][4] ~^ image[21][10] + signed_kernel[2][0] ~^ image[22][6] + signed_kernel[2][1] ~^ image[22][7] + signed_kernel[2][2] ~^ image[22][8] + signed_kernel[2][3] ~^ image[22][9] + signed_kernel[2][4] ~^ image[22][10] + signed_kernel[3][0] ~^ image[23][6] + signed_kernel[3][1] ~^ image[23][7] + signed_kernel[3][2] ~^ image[23][8] + signed_kernel[3][3] ~^ image[23][9] + signed_kernel[3][4] ~^ image[23][10] + signed_kernel[4][0] ~^ image[24][6] + signed_kernel[4][1] ~^ image[24][7] + signed_kernel[4][2] ~^ image[24][8] + signed_kernel[4][3] ~^ image[24][9] + signed_kernel[4][4] ~^ image[24][10];
assign xor_sum[20][7] = signed_kernel[0][0] ~^ image[20][7] + signed_kernel[0][1] ~^ image[20][8] + signed_kernel[0][2] ~^ image[20][9] + signed_kernel[0][3] ~^ image[20][10] + signed_kernel[0][4] ~^ image[20][11] + signed_kernel[1][0] ~^ image[21][7] + signed_kernel[1][1] ~^ image[21][8] + signed_kernel[1][2] ~^ image[21][9] + signed_kernel[1][3] ~^ image[21][10] + signed_kernel[1][4] ~^ image[21][11] + signed_kernel[2][0] ~^ image[22][7] + signed_kernel[2][1] ~^ image[22][8] + signed_kernel[2][2] ~^ image[22][9] + signed_kernel[2][3] ~^ image[22][10] + signed_kernel[2][4] ~^ image[22][11] + signed_kernel[3][0] ~^ image[23][7] + signed_kernel[3][1] ~^ image[23][8] + signed_kernel[3][2] ~^ image[23][9] + signed_kernel[3][3] ~^ image[23][10] + signed_kernel[3][4] ~^ image[23][11] + signed_kernel[4][0] ~^ image[24][7] + signed_kernel[4][1] ~^ image[24][8] + signed_kernel[4][2] ~^ image[24][9] + signed_kernel[4][3] ~^ image[24][10] + signed_kernel[4][4] ~^ image[24][11];
assign xor_sum[20][8] = signed_kernel[0][0] ~^ image[20][8] + signed_kernel[0][1] ~^ image[20][9] + signed_kernel[0][2] ~^ image[20][10] + signed_kernel[0][3] ~^ image[20][11] + signed_kernel[0][4] ~^ image[20][12] + signed_kernel[1][0] ~^ image[21][8] + signed_kernel[1][1] ~^ image[21][9] + signed_kernel[1][2] ~^ image[21][10] + signed_kernel[1][3] ~^ image[21][11] + signed_kernel[1][4] ~^ image[21][12] + signed_kernel[2][0] ~^ image[22][8] + signed_kernel[2][1] ~^ image[22][9] + signed_kernel[2][2] ~^ image[22][10] + signed_kernel[2][3] ~^ image[22][11] + signed_kernel[2][4] ~^ image[22][12] + signed_kernel[3][0] ~^ image[23][8] + signed_kernel[3][1] ~^ image[23][9] + signed_kernel[3][2] ~^ image[23][10] + signed_kernel[3][3] ~^ image[23][11] + signed_kernel[3][4] ~^ image[23][12] + signed_kernel[4][0] ~^ image[24][8] + signed_kernel[4][1] ~^ image[24][9] + signed_kernel[4][2] ~^ image[24][10] + signed_kernel[4][3] ~^ image[24][11] + signed_kernel[4][4] ~^ image[24][12];
assign xor_sum[20][9] = signed_kernel[0][0] ~^ image[20][9] + signed_kernel[0][1] ~^ image[20][10] + signed_kernel[0][2] ~^ image[20][11] + signed_kernel[0][3] ~^ image[20][12] + signed_kernel[0][4] ~^ image[20][13] + signed_kernel[1][0] ~^ image[21][9] + signed_kernel[1][1] ~^ image[21][10] + signed_kernel[1][2] ~^ image[21][11] + signed_kernel[1][3] ~^ image[21][12] + signed_kernel[1][4] ~^ image[21][13] + signed_kernel[2][0] ~^ image[22][9] + signed_kernel[2][1] ~^ image[22][10] + signed_kernel[2][2] ~^ image[22][11] + signed_kernel[2][3] ~^ image[22][12] + signed_kernel[2][4] ~^ image[22][13] + signed_kernel[3][0] ~^ image[23][9] + signed_kernel[3][1] ~^ image[23][10] + signed_kernel[3][2] ~^ image[23][11] + signed_kernel[3][3] ~^ image[23][12] + signed_kernel[3][4] ~^ image[23][13] + signed_kernel[4][0] ~^ image[24][9] + signed_kernel[4][1] ~^ image[24][10] + signed_kernel[4][2] ~^ image[24][11] + signed_kernel[4][3] ~^ image[24][12] + signed_kernel[4][4] ~^ image[24][13];
assign xor_sum[20][10] = signed_kernel[0][0] ~^ image[20][10] + signed_kernel[0][1] ~^ image[20][11] + signed_kernel[0][2] ~^ image[20][12] + signed_kernel[0][3] ~^ image[20][13] + signed_kernel[0][4] ~^ image[20][14] + signed_kernel[1][0] ~^ image[21][10] + signed_kernel[1][1] ~^ image[21][11] + signed_kernel[1][2] ~^ image[21][12] + signed_kernel[1][3] ~^ image[21][13] + signed_kernel[1][4] ~^ image[21][14] + signed_kernel[2][0] ~^ image[22][10] + signed_kernel[2][1] ~^ image[22][11] + signed_kernel[2][2] ~^ image[22][12] + signed_kernel[2][3] ~^ image[22][13] + signed_kernel[2][4] ~^ image[22][14] + signed_kernel[3][0] ~^ image[23][10] + signed_kernel[3][1] ~^ image[23][11] + signed_kernel[3][2] ~^ image[23][12] + signed_kernel[3][3] ~^ image[23][13] + signed_kernel[3][4] ~^ image[23][14] + signed_kernel[4][0] ~^ image[24][10] + signed_kernel[4][1] ~^ image[24][11] + signed_kernel[4][2] ~^ image[24][12] + signed_kernel[4][3] ~^ image[24][13] + signed_kernel[4][4] ~^ image[24][14];
assign xor_sum[20][11] = signed_kernel[0][0] ~^ image[20][11] + signed_kernel[0][1] ~^ image[20][12] + signed_kernel[0][2] ~^ image[20][13] + signed_kernel[0][3] ~^ image[20][14] + signed_kernel[0][4] ~^ image[20][15] + signed_kernel[1][0] ~^ image[21][11] + signed_kernel[1][1] ~^ image[21][12] + signed_kernel[1][2] ~^ image[21][13] + signed_kernel[1][3] ~^ image[21][14] + signed_kernel[1][4] ~^ image[21][15] + signed_kernel[2][0] ~^ image[22][11] + signed_kernel[2][1] ~^ image[22][12] + signed_kernel[2][2] ~^ image[22][13] + signed_kernel[2][3] ~^ image[22][14] + signed_kernel[2][4] ~^ image[22][15] + signed_kernel[3][0] ~^ image[23][11] + signed_kernel[3][1] ~^ image[23][12] + signed_kernel[3][2] ~^ image[23][13] + signed_kernel[3][3] ~^ image[23][14] + signed_kernel[3][4] ~^ image[23][15] + signed_kernel[4][0] ~^ image[24][11] + signed_kernel[4][1] ~^ image[24][12] + signed_kernel[4][2] ~^ image[24][13] + signed_kernel[4][3] ~^ image[24][14] + signed_kernel[4][4] ~^ image[24][15];
assign xor_sum[20][12] = signed_kernel[0][0] ~^ image[20][12] + signed_kernel[0][1] ~^ image[20][13] + signed_kernel[0][2] ~^ image[20][14] + signed_kernel[0][3] ~^ image[20][15] + signed_kernel[0][4] ~^ image[20][16] + signed_kernel[1][0] ~^ image[21][12] + signed_kernel[1][1] ~^ image[21][13] + signed_kernel[1][2] ~^ image[21][14] + signed_kernel[1][3] ~^ image[21][15] + signed_kernel[1][4] ~^ image[21][16] + signed_kernel[2][0] ~^ image[22][12] + signed_kernel[2][1] ~^ image[22][13] + signed_kernel[2][2] ~^ image[22][14] + signed_kernel[2][3] ~^ image[22][15] + signed_kernel[2][4] ~^ image[22][16] + signed_kernel[3][0] ~^ image[23][12] + signed_kernel[3][1] ~^ image[23][13] + signed_kernel[3][2] ~^ image[23][14] + signed_kernel[3][3] ~^ image[23][15] + signed_kernel[3][4] ~^ image[23][16] + signed_kernel[4][0] ~^ image[24][12] + signed_kernel[4][1] ~^ image[24][13] + signed_kernel[4][2] ~^ image[24][14] + signed_kernel[4][3] ~^ image[24][15] + signed_kernel[4][4] ~^ image[24][16];
assign xor_sum[20][13] = signed_kernel[0][0] ~^ image[20][13] + signed_kernel[0][1] ~^ image[20][14] + signed_kernel[0][2] ~^ image[20][15] + signed_kernel[0][3] ~^ image[20][16] + signed_kernel[0][4] ~^ image[20][17] + signed_kernel[1][0] ~^ image[21][13] + signed_kernel[1][1] ~^ image[21][14] + signed_kernel[1][2] ~^ image[21][15] + signed_kernel[1][3] ~^ image[21][16] + signed_kernel[1][4] ~^ image[21][17] + signed_kernel[2][0] ~^ image[22][13] + signed_kernel[2][1] ~^ image[22][14] + signed_kernel[2][2] ~^ image[22][15] + signed_kernel[2][3] ~^ image[22][16] + signed_kernel[2][4] ~^ image[22][17] + signed_kernel[3][0] ~^ image[23][13] + signed_kernel[3][1] ~^ image[23][14] + signed_kernel[3][2] ~^ image[23][15] + signed_kernel[3][3] ~^ image[23][16] + signed_kernel[3][4] ~^ image[23][17] + signed_kernel[4][0] ~^ image[24][13] + signed_kernel[4][1] ~^ image[24][14] + signed_kernel[4][2] ~^ image[24][15] + signed_kernel[4][3] ~^ image[24][16] + signed_kernel[4][4] ~^ image[24][17];
assign xor_sum[20][14] = signed_kernel[0][0] ~^ image[20][14] + signed_kernel[0][1] ~^ image[20][15] + signed_kernel[0][2] ~^ image[20][16] + signed_kernel[0][3] ~^ image[20][17] + signed_kernel[0][4] ~^ image[20][18] + signed_kernel[1][0] ~^ image[21][14] + signed_kernel[1][1] ~^ image[21][15] + signed_kernel[1][2] ~^ image[21][16] + signed_kernel[1][3] ~^ image[21][17] + signed_kernel[1][4] ~^ image[21][18] + signed_kernel[2][0] ~^ image[22][14] + signed_kernel[2][1] ~^ image[22][15] + signed_kernel[2][2] ~^ image[22][16] + signed_kernel[2][3] ~^ image[22][17] + signed_kernel[2][4] ~^ image[22][18] + signed_kernel[3][0] ~^ image[23][14] + signed_kernel[3][1] ~^ image[23][15] + signed_kernel[3][2] ~^ image[23][16] + signed_kernel[3][3] ~^ image[23][17] + signed_kernel[3][4] ~^ image[23][18] + signed_kernel[4][0] ~^ image[24][14] + signed_kernel[4][1] ~^ image[24][15] + signed_kernel[4][2] ~^ image[24][16] + signed_kernel[4][3] ~^ image[24][17] + signed_kernel[4][4] ~^ image[24][18];
assign xor_sum[20][15] = signed_kernel[0][0] ~^ image[20][15] + signed_kernel[0][1] ~^ image[20][16] + signed_kernel[0][2] ~^ image[20][17] + signed_kernel[0][3] ~^ image[20][18] + signed_kernel[0][4] ~^ image[20][19] + signed_kernel[1][0] ~^ image[21][15] + signed_kernel[1][1] ~^ image[21][16] + signed_kernel[1][2] ~^ image[21][17] + signed_kernel[1][3] ~^ image[21][18] + signed_kernel[1][4] ~^ image[21][19] + signed_kernel[2][0] ~^ image[22][15] + signed_kernel[2][1] ~^ image[22][16] + signed_kernel[2][2] ~^ image[22][17] + signed_kernel[2][3] ~^ image[22][18] + signed_kernel[2][4] ~^ image[22][19] + signed_kernel[3][0] ~^ image[23][15] + signed_kernel[3][1] ~^ image[23][16] + signed_kernel[3][2] ~^ image[23][17] + signed_kernel[3][3] ~^ image[23][18] + signed_kernel[3][4] ~^ image[23][19] + signed_kernel[4][0] ~^ image[24][15] + signed_kernel[4][1] ~^ image[24][16] + signed_kernel[4][2] ~^ image[24][17] + signed_kernel[4][3] ~^ image[24][18] + signed_kernel[4][4] ~^ image[24][19];
assign xor_sum[20][16] = signed_kernel[0][0] ~^ image[20][16] + signed_kernel[0][1] ~^ image[20][17] + signed_kernel[0][2] ~^ image[20][18] + signed_kernel[0][3] ~^ image[20][19] + signed_kernel[0][4] ~^ image[20][20] + signed_kernel[1][0] ~^ image[21][16] + signed_kernel[1][1] ~^ image[21][17] + signed_kernel[1][2] ~^ image[21][18] + signed_kernel[1][3] ~^ image[21][19] + signed_kernel[1][4] ~^ image[21][20] + signed_kernel[2][0] ~^ image[22][16] + signed_kernel[2][1] ~^ image[22][17] + signed_kernel[2][2] ~^ image[22][18] + signed_kernel[2][3] ~^ image[22][19] + signed_kernel[2][4] ~^ image[22][20] + signed_kernel[3][0] ~^ image[23][16] + signed_kernel[3][1] ~^ image[23][17] + signed_kernel[3][2] ~^ image[23][18] + signed_kernel[3][3] ~^ image[23][19] + signed_kernel[3][4] ~^ image[23][20] + signed_kernel[4][0] ~^ image[24][16] + signed_kernel[4][1] ~^ image[24][17] + signed_kernel[4][2] ~^ image[24][18] + signed_kernel[4][3] ~^ image[24][19] + signed_kernel[4][4] ~^ image[24][20];
assign xor_sum[20][17] = signed_kernel[0][0] ~^ image[20][17] + signed_kernel[0][1] ~^ image[20][18] + signed_kernel[0][2] ~^ image[20][19] + signed_kernel[0][3] ~^ image[20][20] + signed_kernel[0][4] ~^ image[20][21] + signed_kernel[1][0] ~^ image[21][17] + signed_kernel[1][1] ~^ image[21][18] + signed_kernel[1][2] ~^ image[21][19] + signed_kernel[1][3] ~^ image[21][20] + signed_kernel[1][4] ~^ image[21][21] + signed_kernel[2][0] ~^ image[22][17] + signed_kernel[2][1] ~^ image[22][18] + signed_kernel[2][2] ~^ image[22][19] + signed_kernel[2][3] ~^ image[22][20] + signed_kernel[2][4] ~^ image[22][21] + signed_kernel[3][0] ~^ image[23][17] + signed_kernel[3][1] ~^ image[23][18] + signed_kernel[3][2] ~^ image[23][19] + signed_kernel[3][3] ~^ image[23][20] + signed_kernel[3][4] ~^ image[23][21] + signed_kernel[4][0] ~^ image[24][17] + signed_kernel[4][1] ~^ image[24][18] + signed_kernel[4][2] ~^ image[24][19] + signed_kernel[4][3] ~^ image[24][20] + signed_kernel[4][4] ~^ image[24][21];
assign xor_sum[20][18] = signed_kernel[0][0] ~^ image[20][18] + signed_kernel[0][1] ~^ image[20][19] + signed_kernel[0][2] ~^ image[20][20] + signed_kernel[0][3] ~^ image[20][21] + signed_kernel[0][4] ~^ image[20][22] + signed_kernel[1][0] ~^ image[21][18] + signed_kernel[1][1] ~^ image[21][19] + signed_kernel[1][2] ~^ image[21][20] + signed_kernel[1][3] ~^ image[21][21] + signed_kernel[1][4] ~^ image[21][22] + signed_kernel[2][0] ~^ image[22][18] + signed_kernel[2][1] ~^ image[22][19] + signed_kernel[2][2] ~^ image[22][20] + signed_kernel[2][3] ~^ image[22][21] + signed_kernel[2][4] ~^ image[22][22] + signed_kernel[3][0] ~^ image[23][18] + signed_kernel[3][1] ~^ image[23][19] + signed_kernel[3][2] ~^ image[23][20] + signed_kernel[3][3] ~^ image[23][21] + signed_kernel[3][4] ~^ image[23][22] + signed_kernel[4][0] ~^ image[24][18] + signed_kernel[4][1] ~^ image[24][19] + signed_kernel[4][2] ~^ image[24][20] + signed_kernel[4][3] ~^ image[24][21] + signed_kernel[4][4] ~^ image[24][22];
assign xor_sum[20][19] = signed_kernel[0][0] ~^ image[20][19] + signed_kernel[0][1] ~^ image[20][20] + signed_kernel[0][2] ~^ image[20][21] + signed_kernel[0][3] ~^ image[20][22] + signed_kernel[0][4] ~^ image[20][23] + signed_kernel[1][0] ~^ image[21][19] + signed_kernel[1][1] ~^ image[21][20] + signed_kernel[1][2] ~^ image[21][21] + signed_kernel[1][3] ~^ image[21][22] + signed_kernel[1][4] ~^ image[21][23] + signed_kernel[2][0] ~^ image[22][19] + signed_kernel[2][1] ~^ image[22][20] + signed_kernel[2][2] ~^ image[22][21] + signed_kernel[2][3] ~^ image[22][22] + signed_kernel[2][4] ~^ image[22][23] + signed_kernel[3][0] ~^ image[23][19] + signed_kernel[3][1] ~^ image[23][20] + signed_kernel[3][2] ~^ image[23][21] + signed_kernel[3][3] ~^ image[23][22] + signed_kernel[3][4] ~^ image[23][23] + signed_kernel[4][0] ~^ image[24][19] + signed_kernel[4][1] ~^ image[24][20] + signed_kernel[4][2] ~^ image[24][21] + signed_kernel[4][3] ~^ image[24][22] + signed_kernel[4][4] ~^ image[24][23];
assign xor_sum[20][20] = signed_kernel[0][0] ~^ image[20][20] + signed_kernel[0][1] ~^ image[20][21] + signed_kernel[0][2] ~^ image[20][22] + signed_kernel[0][3] ~^ image[20][23] + signed_kernel[0][4] ~^ image[20][24] + signed_kernel[1][0] ~^ image[21][20] + signed_kernel[1][1] ~^ image[21][21] + signed_kernel[1][2] ~^ image[21][22] + signed_kernel[1][3] ~^ image[21][23] + signed_kernel[1][4] ~^ image[21][24] + signed_kernel[2][0] ~^ image[22][20] + signed_kernel[2][1] ~^ image[22][21] + signed_kernel[2][2] ~^ image[22][22] + signed_kernel[2][3] ~^ image[22][23] + signed_kernel[2][4] ~^ image[22][24] + signed_kernel[3][0] ~^ image[23][20] + signed_kernel[3][1] ~^ image[23][21] + signed_kernel[3][2] ~^ image[23][22] + signed_kernel[3][3] ~^ image[23][23] + signed_kernel[3][4] ~^ image[23][24] + signed_kernel[4][0] ~^ image[24][20] + signed_kernel[4][1] ~^ image[24][21] + signed_kernel[4][2] ~^ image[24][22] + signed_kernel[4][3] ~^ image[24][23] + signed_kernel[4][4] ~^ image[24][24];
assign xor_sum[20][21] = signed_kernel[0][0] ~^ image[20][21] + signed_kernel[0][1] ~^ image[20][22] + signed_kernel[0][2] ~^ image[20][23] + signed_kernel[0][3] ~^ image[20][24] + signed_kernel[0][4] ~^ image[20][25] + signed_kernel[1][0] ~^ image[21][21] + signed_kernel[1][1] ~^ image[21][22] + signed_kernel[1][2] ~^ image[21][23] + signed_kernel[1][3] ~^ image[21][24] + signed_kernel[1][4] ~^ image[21][25] + signed_kernel[2][0] ~^ image[22][21] + signed_kernel[2][1] ~^ image[22][22] + signed_kernel[2][2] ~^ image[22][23] + signed_kernel[2][3] ~^ image[22][24] + signed_kernel[2][4] ~^ image[22][25] + signed_kernel[3][0] ~^ image[23][21] + signed_kernel[3][1] ~^ image[23][22] + signed_kernel[3][2] ~^ image[23][23] + signed_kernel[3][3] ~^ image[23][24] + signed_kernel[3][4] ~^ image[23][25] + signed_kernel[4][0] ~^ image[24][21] + signed_kernel[4][1] ~^ image[24][22] + signed_kernel[4][2] ~^ image[24][23] + signed_kernel[4][3] ~^ image[24][24] + signed_kernel[4][4] ~^ image[24][25];
assign xor_sum[20][22] = signed_kernel[0][0] ~^ image[20][22] + signed_kernel[0][1] ~^ image[20][23] + signed_kernel[0][2] ~^ image[20][24] + signed_kernel[0][3] ~^ image[20][25] + signed_kernel[0][4] ~^ image[20][26] + signed_kernel[1][0] ~^ image[21][22] + signed_kernel[1][1] ~^ image[21][23] + signed_kernel[1][2] ~^ image[21][24] + signed_kernel[1][3] ~^ image[21][25] + signed_kernel[1][4] ~^ image[21][26] + signed_kernel[2][0] ~^ image[22][22] + signed_kernel[2][1] ~^ image[22][23] + signed_kernel[2][2] ~^ image[22][24] + signed_kernel[2][3] ~^ image[22][25] + signed_kernel[2][4] ~^ image[22][26] + signed_kernel[3][0] ~^ image[23][22] + signed_kernel[3][1] ~^ image[23][23] + signed_kernel[3][2] ~^ image[23][24] + signed_kernel[3][3] ~^ image[23][25] + signed_kernel[3][4] ~^ image[23][26] + signed_kernel[4][0] ~^ image[24][22] + signed_kernel[4][1] ~^ image[24][23] + signed_kernel[4][2] ~^ image[24][24] + signed_kernel[4][3] ~^ image[24][25] + signed_kernel[4][4] ~^ image[24][26];
assign xor_sum[20][23] = signed_kernel[0][0] ~^ image[20][23] + signed_kernel[0][1] ~^ image[20][24] + signed_kernel[0][2] ~^ image[20][25] + signed_kernel[0][3] ~^ image[20][26] + signed_kernel[0][4] ~^ image[20][27] + signed_kernel[1][0] ~^ image[21][23] + signed_kernel[1][1] ~^ image[21][24] + signed_kernel[1][2] ~^ image[21][25] + signed_kernel[1][3] ~^ image[21][26] + signed_kernel[1][4] ~^ image[21][27] + signed_kernel[2][0] ~^ image[22][23] + signed_kernel[2][1] ~^ image[22][24] + signed_kernel[2][2] ~^ image[22][25] + signed_kernel[2][3] ~^ image[22][26] + signed_kernel[2][4] ~^ image[22][27] + signed_kernel[3][0] ~^ image[23][23] + signed_kernel[3][1] ~^ image[23][24] + signed_kernel[3][2] ~^ image[23][25] + signed_kernel[3][3] ~^ image[23][26] + signed_kernel[3][4] ~^ image[23][27] + signed_kernel[4][0] ~^ image[24][23] + signed_kernel[4][1] ~^ image[24][24] + signed_kernel[4][2] ~^ image[24][25] + signed_kernel[4][3] ~^ image[24][26] + signed_kernel[4][4] ~^ image[24][27];
assign xor_sum[21][0] = signed_kernel[0][0] ~^ image[21][0] + signed_kernel[0][1] ~^ image[21][1] + signed_kernel[0][2] ~^ image[21][2] + signed_kernel[0][3] ~^ image[21][3] + signed_kernel[0][4] ~^ image[21][4] + signed_kernel[1][0] ~^ image[22][0] + signed_kernel[1][1] ~^ image[22][1] + signed_kernel[1][2] ~^ image[22][2] + signed_kernel[1][3] ~^ image[22][3] + signed_kernel[1][4] ~^ image[22][4] + signed_kernel[2][0] ~^ image[23][0] + signed_kernel[2][1] ~^ image[23][1] + signed_kernel[2][2] ~^ image[23][2] + signed_kernel[2][3] ~^ image[23][3] + signed_kernel[2][4] ~^ image[23][4] + signed_kernel[3][0] ~^ image[24][0] + signed_kernel[3][1] ~^ image[24][1] + signed_kernel[3][2] ~^ image[24][2] + signed_kernel[3][3] ~^ image[24][3] + signed_kernel[3][4] ~^ image[24][4] + signed_kernel[4][0] ~^ image[25][0] + signed_kernel[4][1] ~^ image[25][1] + signed_kernel[4][2] ~^ image[25][2] + signed_kernel[4][3] ~^ image[25][3] + signed_kernel[4][4] ~^ image[25][4];
assign xor_sum[21][1] = signed_kernel[0][0] ~^ image[21][1] + signed_kernel[0][1] ~^ image[21][2] + signed_kernel[0][2] ~^ image[21][3] + signed_kernel[0][3] ~^ image[21][4] + signed_kernel[0][4] ~^ image[21][5] + signed_kernel[1][0] ~^ image[22][1] + signed_kernel[1][1] ~^ image[22][2] + signed_kernel[1][2] ~^ image[22][3] + signed_kernel[1][3] ~^ image[22][4] + signed_kernel[1][4] ~^ image[22][5] + signed_kernel[2][0] ~^ image[23][1] + signed_kernel[2][1] ~^ image[23][2] + signed_kernel[2][2] ~^ image[23][3] + signed_kernel[2][3] ~^ image[23][4] + signed_kernel[2][4] ~^ image[23][5] + signed_kernel[3][0] ~^ image[24][1] + signed_kernel[3][1] ~^ image[24][2] + signed_kernel[3][2] ~^ image[24][3] + signed_kernel[3][3] ~^ image[24][4] + signed_kernel[3][4] ~^ image[24][5] + signed_kernel[4][0] ~^ image[25][1] + signed_kernel[4][1] ~^ image[25][2] + signed_kernel[4][2] ~^ image[25][3] + signed_kernel[4][3] ~^ image[25][4] + signed_kernel[4][4] ~^ image[25][5];
assign xor_sum[21][2] = signed_kernel[0][0] ~^ image[21][2] + signed_kernel[0][1] ~^ image[21][3] + signed_kernel[0][2] ~^ image[21][4] + signed_kernel[0][3] ~^ image[21][5] + signed_kernel[0][4] ~^ image[21][6] + signed_kernel[1][0] ~^ image[22][2] + signed_kernel[1][1] ~^ image[22][3] + signed_kernel[1][2] ~^ image[22][4] + signed_kernel[1][3] ~^ image[22][5] + signed_kernel[1][4] ~^ image[22][6] + signed_kernel[2][0] ~^ image[23][2] + signed_kernel[2][1] ~^ image[23][3] + signed_kernel[2][2] ~^ image[23][4] + signed_kernel[2][3] ~^ image[23][5] + signed_kernel[2][4] ~^ image[23][6] + signed_kernel[3][0] ~^ image[24][2] + signed_kernel[3][1] ~^ image[24][3] + signed_kernel[3][2] ~^ image[24][4] + signed_kernel[3][3] ~^ image[24][5] + signed_kernel[3][4] ~^ image[24][6] + signed_kernel[4][0] ~^ image[25][2] + signed_kernel[4][1] ~^ image[25][3] + signed_kernel[4][2] ~^ image[25][4] + signed_kernel[4][3] ~^ image[25][5] + signed_kernel[4][4] ~^ image[25][6];
assign xor_sum[21][3] = signed_kernel[0][0] ~^ image[21][3] + signed_kernel[0][1] ~^ image[21][4] + signed_kernel[0][2] ~^ image[21][5] + signed_kernel[0][3] ~^ image[21][6] + signed_kernel[0][4] ~^ image[21][7] + signed_kernel[1][0] ~^ image[22][3] + signed_kernel[1][1] ~^ image[22][4] + signed_kernel[1][2] ~^ image[22][5] + signed_kernel[1][3] ~^ image[22][6] + signed_kernel[1][4] ~^ image[22][7] + signed_kernel[2][0] ~^ image[23][3] + signed_kernel[2][1] ~^ image[23][4] + signed_kernel[2][2] ~^ image[23][5] + signed_kernel[2][3] ~^ image[23][6] + signed_kernel[2][4] ~^ image[23][7] + signed_kernel[3][0] ~^ image[24][3] + signed_kernel[3][1] ~^ image[24][4] + signed_kernel[3][2] ~^ image[24][5] + signed_kernel[3][3] ~^ image[24][6] + signed_kernel[3][4] ~^ image[24][7] + signed_kernel[4][0] ~^ image[25][3] + signed_kernel[4][1] ~^ image[25][4] + signed_kernel[4][2] ~^ image[25][5] + signed_kernel[4][3] ~^ image[25][6] + signed_kernel[4][4] ~^ image[25][7];
assign xor_sum[21][4] = signed_kernel[0][0] ~^ image[21][4] + signed_kernel[0][1] ~^ image[21][5] + signed_kernel[0][2] ~^ image[21][6] + signed_kernel[0][3] ~^ image[21][7] + signed_kernel[0][4] ~^ image[21][8] + signed_kernel[1][0] ~^ image[22][4] + signed_kernel[1][1] ~^ image[22][5] + signed_kernel[1][2] ~^ image[22][6] + signed_kernel[1][3] ~^ image[22][7] + signed_kernel[1][4] ~^ image[22][8] + signed_kernel[2][0] ~^ image[23][4] + signed_kernel[2][1] ~^ image[23][5] + signed_kernel[2][2] ~^ image[23][6] + signed_kernel[2][3] ~^ image[23][7] + signed_kernel[2][4] ~^ image[23][8] + signed_kernel[3][0] ~^ image[24][4] + signed_kernel[3][1] ~^ image[24][5] + signed_kernel[3][2] ~^ image[24][6] + signed_kernel[3][3] ~^ image[24][7] + signed_kernel[3][4] ~^ image[24][8] + signed_kernel[4][0] ~^ image[25][4] + signed_kernel[4][1] ~^ image[25][5] + signed_kernel[4][2] ~^ image[25][6] + signed_kernel[4][3] ~^ image[25][7] + signed_kernel[4][4] ~^ image[25][8];
assign xor_sum[21][5] = signed_kernel[0][0] ~^ image[21][5] + signed_kernel[0][1] ~^ image[21][6] + signed_kernel[0][2] ~^ image[21][7] + signed_kernel[0][3] ~^ image[21][8] + signed_kernel[0][4] ~^ image[21][9] + signed_kernel[1][0] ~^ image[22][5] + signed_kernel[1][1] ~^ image[22][6] + signed_kernel[1][2] ~^ image[22][7] + signed_kernel[1][3] ~^ image[22][8] + signed_kernel[1][4] ~^ image[22][9] + signed_kernel[2][0] ~^ image[23][5] + signed_kernel[2][1] ~^ image[23][6] + signed_kernel[2][2] ~^ image[23][7] + signed_kernel[2][3] ~^ image[23][8] + signed_kernel[2][4] ~^ image[23][9] + signed_kernel[3][0] ~^ image[24][5] + signed_kernel[3][1] ~^ image[24][6] + signed_kernel[3][2] ~^ image[24][7] + signed_kernel[3][3] ~^ image[24][8] + signed_kernel[3][4] ~^ image[24][9] + signed_kernel[4][0] ~^ image[25][5] + signed_kernel[4][1] ~^ image[25][6] + signed_kernel[4][2] ~^ image[25][7] + signed_kernel[4][3] ~^ image[25][8] + signed_kernel[4][4] ~^ image[25][9];
assign xor_sum[21][6] = signed_kernel[0][0] ~^ image[21][6] + signed_kernel[0][1] ~^ image[21][7] + signed_kernel[0][2] ~^ image[21][8] + signed_kernel[0][3] ~^ image[21][9] + signed_kernel[0][4] ~^ image[21][10] + signed_kernel[1][0] ~^ image[22][6] + signed_kernel[1][1] ~^ image[22][7] + signed_kernel[1][2] ~^ image[22][8] + signed_kernel[1][3] ~^ image[22][9] + signed_kernel[1][4] ~^ image[22][10] + signed_kernel[2][0] ~^ image[23][6] + signed_kernel[2][1] ~^ image[23][7] + signed_kernel[2][2] ~^ image[23][8] + signed_kernel[2][3] ~^ image[23][9] + signed_kernel[2][4] ~^ image[23][10] + signed_kernel[3][0] ~^ image[24][6] + signed_kernel[3][1] ~^ image[24][7] + signed_kernel[3][2] ~^ image[24][8] + signed_kernel[3][3] ~^ image[24][9] + signed_kernel[3][4] ~^ image[24][10] + signed_kernel[4][0] ~^ image[25][6] + signed_kernel[4][1] ~^ image[25][7] + signed_kernel[4][2] ~^ image[25][8] + signed_kernel[4][3] ~^ image[25][9] + signed_kernel[4][4] ~^ image[25][10];
assign xor_sum[21][7] = signed_kernel[0][0] ~^ image[21][7] + signed_kernel[0][1] ~^ image[21][8] + signed_kernel[0][2] ~^ image[21][9] + signed_kernel[0][3] ~^ image[21][10] + signed_kernel[0][4] ~^ image[21][11] + signed_kernel[1][0] ~^ image[22][7] + signed_kernel[1][1] ~^ image[22][8] + signed_kernel[1][2] ~^ image[22][9] + signed_kernel[1][3] ~^ image[22][10] + signed_kernel[1][4] ~^ image[22][11] + signed_kernel[2][0] ~^ image[23][7] + signed_kernel[2][1] ~^ image[23][8] + signed_kernel[2][2] ~^ image[23][9] + signed_kernel[2][3] ~^ image[23][10] + signed_kernel[2][4] ~^ image[23][11] + signed_kernel[3][0] ~^ image[24][7] + signed_kernel[3][1] ~^ image[24][8] + signed_kernel[3][2] ~^ image[24][9] + signed_kernel[3][3] ~^ image[24][10] + signed_kernel[3][4] ~^ image[24][11] + signed_kernel[4][0] ~^ image[25][7] + signed_kernel[4][1] ~^ image[25][8] + signed_kernel[4][2] ~^ image[25][9] + signed_kernel[4][3] ~^ image[25][10] + signed_kernel[4][4] ~^ image[25][11];
assign xor_sum[21][8] = signed_kernel[0][0] ~^ image[21][8] + signed_kernel[0][1] ~^ image[21][9] + signed_kernel[0][2] ~^ image[21][10] + signed_kernel[0][3] ~^ image[21][11] + signed_kernel[0][4] ~^ image[21][12] + signed_kernel[1][0] ~^ image[22][8] + signed_kernel[1][1] ~^ image[22][9] + signed_kernel[1][2] ~^ image[22][10] + signed_kernel[1][3] ~^ image[22][11] + signed_kernel[1][4] ~^ image[22][12] + signed_kernel[2][0] ~^ image[23][8] + signed_kernel[2][1] ~^ image[23][9] + signed_kernel[2][2] ~^ image[23][10] + signed_kernel[2][3] ~^ image[23][11] + signed_kernel[2][4] ~^ image[23][12] + signed_kernel[3][0] ~^ image[24][8] + signed_kernel[3][1] ~^ image[24][9] + signed_kernel[3][2] ~^ image[24][10] + signed_kernel[3][3] ~^ image[24][11] + signed_kernel[3][4] ~^ image[24][12] + signed_kernel[4][0] ~^ image[25][8] + signed_kernel[4][1] ~^ image[25][9] + signed_kernel[4][2] ~^ image[25][10] + signed_kernel[4][3] ~^ image[25][11] + signed_kernel[4][4] ~^ image[25][12];
assign xor_sum[21][9] = signed_kernel[0][0] ~^ image[21][9] + signed_kernel[0][1] ~^ image[21][10] + signed_kernel[0][2] ~^ image[21][11] + signed_kernel[0][3] ~^ image[21][12] + signed_kernel[0][4] ~^ image[21][13] + signed_kernel[1][0] ~^ image[22][9] + signed_kernel[1][1] ~^ image[22][10] + signed_kernel[1][2] ~^ image[22][11] + signed_kernel[1][3] ~^ image[22][12] + signed_kernel[1][4] ~^ image[22][13] + signed_kernel[2][0] ~^ image[23][9] + signed_kernel[2][1] ~^ image[23][10] + signed_kernel[2][2] ~^ image[23][11] + signed_kernel[2][3] ~^ image[23][12] + signed_kernel[2][4] ~^ image[23][13] + signed_kernel[3][0] ~^ image[24][9] + signed_kernel[3][1] ~^ image[24][10] + signed_kernel[3][2] ~^ image[24][11] + signed_kernel[3][3] ~^ image[24][12] + signed_kernel[3][4] ~^ image[24][13] + signed_kernel[4][0] ~^ image[25][9] + signed_kernel[4][1] ~^ image[25][10] + signed_kernel[4][2] ~^ image[25][11] + signed_kernel[4][3] ~^ image[25][12] + signed_kernel[4][4] ~^ image[25][13];
assign xor_sum[21][10] = signed_kernel[0][0] ~^ image[21][10] + signed_kernel[0][1] ~^ image[21][11] + signed_kernel[0][2] ~^ image[21][12] + signed_kernel[0][3] ~^ image[21][13] + signed_kernel[0][4] ~^ image[21][14] + signed_kernel[1][0] ~^ image[22][10] + signed_kernel[1][1] ~^ image[22][11] + signed_kernel[1][2] ~^ image[22][12] + signed_kernel[1][3] ~^ image[22][13] + signed_kernel[1][4] ~^ image[22][14] + signed_kernel[2][0] ~^ image[23][10] + signed_kernel[2][1] ~^ image[23][11] + signed_kernel[2][2] ~^ image[23][12] + signed_kernel[2][3] ~^ image[23][13] + signed_kernel[2][4] ~^ image[23][14] + signed_kernel[3][0] ~^ image[24][10] + signed_kernel[3][1] ~^ image[24][11] + signed_kernel[3][2] ~^ image[24][12] + signed_kernel[3][3] ~^ image[24][13] + signed_kernel[3][4] ~^ image[24][14] + signed_kernel[4][0] ~^ image[25][10] + signed_kernel[4][1] ~^ image[25][11] + signed_kernel[4][2] ~^ image[25][12] + signed_kernel[4][3] ~^ image[25][13] + signed_kernel[4][4] ~^ image[25][14];
assign xor_sum[21][11] = signed_kernel[0][0] ~^ image[21][11] + signed_kernel[0][1] ~^ image[21][12] + signed_kernel[0][2] ~^ image[21][13] + signed_kernel[0][3] ~^ image[21][14] + signed_kernel[0][4] ~^ image[21][15] + signed_kernel[1][0] ~^ image[22][11] + signed_kernel[1][1] ~^ image[22][12] + signed_kernel[1][2] ~^ image[22][13] + signed_kernel[1][3] ~^ image[22][14] + signed_kernel[1][4] ~^ image[22][15] + signed_kernel[2][0] ~^ image[23][11] + signed_kernel[2][1] ~^ image[23][12] + signed_kernel[2][2] ~^ image[23][13] + signed_kernel[2][3] ~^ image[23][14] + signed_kernel[2][4] ~^ image[23][15] + signed_kernel[3][0] ~^ image[24][11] + signed_kernel[3][1] ~^ image[24][12] + signed_kernel[3][2] ~^ image[24][13] + signed_kernel[3][3] ~^ image[24][14] + signed_kernel[3][4] ~^ image[24][15] + signed_kernel[4][0] ~^ image[25][11] + signed_kernel[4][1] ~^ image[25][12] + signed_kernel[4][2] ~^ image[25][13] + signed_kernel[4][3] ~^ image[25][14] + signed_kernel[4][4] ~^ image[25][15];
assign xor_sum[21][12] = signed_kernel[0][0] ~^ image[21][12] + signed_kernel[0][1] ~^ image[21][13] + signed_kernel[0][2] ~^ image[21][14] + signed_kernel[0][3] ~^ image[21][15] + signed_kernel[0][4] ~^ image[21][16] + signed_kernel[1][0] ~^ image[22][12] + signed_kernel[1][1] ~^ image[22][13] + signed_kernel[1][2] ~^ image[22][14] + signed_kernel[1][3] ~^ image[22][15] + signed_kernel[1][4] ~^ image[22][16] + signed_kernel[2][0] ~^ image[23][12] + signed_kernel[2][1] ~^ image[23][13] + signed_kernel[2][2] ~^ image[23][14] + signed_kernel[2][3] ~^ image[23][15] + signed_kernel[2][4] ~^ image[23][16] + signed_kernel[3][0] ~^ image[24][12] + signed_kernel[3][1] ~^ image[24][13] + signed_kernel[3][2] ~^ image[24][14] + signed_kernel[3][3] ~^ image[24][15] + signed_kernel[3][4] ~^ image[24][16] + signed_kernel[4][0] ~^ image[25][12] + signed_kernel[4][1] ~^ image[25][13] + signed_kernel[4][2] ~^ image[25][14] + signed_kernel[4][3] ~^ image[25][15] + signed_kernel[4][4] ~^ image[25][16];
assign xor_sum[21][13] = signed_kernel[0][0] ~^ image[21][13] + signed_kernel[0][1] ~^ image[21][14] + signed_kernel[0][2] ~^ image[21][15] + signed_kernel[0][3] ~^ image[21][16] + signed_kernel[0][4] ~^ image[21][17] + signed_kernel[1][0] ~^ image[22][13] + signed_kernel[1][1] ~^ image[22][14] + signed_kernel[1][2] ~^ image[22][15] + signed_kernel[1][3] ~^ image[22][16] + signed_kernel[1][4] ~^ image[22][17] + signed_kernel[2][0] ~^ image[23][13] + signed_kernel[2][1] ~^ image[23][14] + signed_kernel[2][2] ~^ image[23][15] + signed_kernel[2][3] ~^ image[23][16] + signed_kernel[2][4] ~^ image[23][17] + signed_kernel[3][0] ~^ image[24][13] + signed_kernel[3][1] ~^ image[24][14] + signed_kernel[3][2] ~^ image[24][15] + signed_kernel[3][3] ~^ image[24][16] + signed_kernel[3][4] ~^ image[24][17] + signed_kernel[4][0] ~^ image[25][13] + signed_kernel[4][1] ~^ image[25][14] + signed_kernel[4][2] ~^ image[25][15] + signed_kernel[4][3] ~^ image[25][16] + signed_kernel[4][4] ~^ image[25][17];
assign xor_sum[21][14] = signed_kernel[0][0] ~^ image[21][14] + signed_kernel[0][1] ~^ image[21][15] + signed_kernel[0][2] ~^ image[21][16] + signed_kernel[0][3] ~^ image[21][17] + signed_kernel[0][4] ~^ image[21][18] + signed_kernel[1][0] ~^ image[22][14] + signed_kernel[1][1] ~^ image[22][15] + signed_kernel[1][2] ~^ image[22][16] + signed_kernel[1][3] ~^ image[22][17] + signed_kernel[1][4] ~^ image[22][18] + signed_kernel[2][0] ~^ image[23][14] + signed_kernel[2][1] ~^ image[23][15] + signed_kernel[2][2] ~^ image[23][16] + signed_kernel[2][3] ~^ image[23][17] + signed_kernel[2][4] ~^ image[23][18] + signed_kernel[3][0] ~^ image[24][14] + signed_kernel[3][1] ~^ image[24][15] + signed_kernel[3][2] ~^ image[24][16] + signed_kernel[3][3] ~^ image[24][17] + signed_kernel[3][4] ~^ image[24][18] + signed_kernel[4][0] ~^ image[25][14] + signed_kernel[4][1] ~^ image[25][15] + signed_kernel[4][2] ~^ image[25][16] + signed_kernel[4][3] ~^ image[25][17] + signed_kernel[4][4] ~^ image[25][18];
assign xor_sum[21][15] = signed_kernel[0][0] ~^ image[21][15] + signed_kernel[0][1] ~^ image[21][16] + signed_kernel[0][2] ~^ image[21][17] + signed_kernel[0][3] ~^ image[21][18] + signed_kernel[0][4] ~^ image[21][19] + signed_kernel[1][0] ~^ image[22][15] + signed_kernel[1][1] ~^ image[22][16] + signed_kernel[1][2] ~^ image[22][17] + signed_kernel[1][3] ~^ image[22][18] + signed_kernel[1][4] ~^ image[22][19] + signed_kernel[2][0] ~^ image[23][15] + signed_kernel[2][1] ~^ image[23][16] + signed_kernel[2][2] ~^ image[23][17] + signed_kernel[2][3] ~^ image[23][18] + signed_kernel[2][4] ~^ image[23][19] + signed_kernel[3][0] ~^ image[24][15] + signed_kernel[3][1] ~^ image[24][16] + signed_kernel[3][2] ~^ image[24][17] + signed_kernel[3][3] ~^ image[24][18] + signed_kernel[3][4] ~^ image[24][19] + signed_kernel[4][0] ~^ image[25][15] + signed_kernel[4][1] ~^ image[25][16] + signed_kernel[4][2] ~^ image[25][17] + signed_kernel[4][3] ~^ image[25][18] + signed_kernel[4][4] ~^ image[25][19];
assign xor_sum[21][16] = signed_kernel[0][0] ~^ image[21][16] + signed_kernel[0][1] ~^ image[21][17] + signed_kernel[0][2] ~^ image[21][18] + signed_kernel[0][3] ~^ image[21][19] + signed_kernel[0][4] ~^ image[21][20] + signed_kernel[1][0] ~^ image[22][16] + signed_kernel[1][1] ~^ image[22][17] + signed_kernel[1][2] ~^ image[22][18] + signed_kernel[1][3] ~^ image[22][19] + signed_kernel[1][4] ~^ image[22][20] + signed_kernel[2][0] ~^ image[23][16] + signed_kernel[2][1] ~^ image[23][17] + signed_kernel[2][2] ~^ image[23][18] + signed_kernel[2][3] ~^ image[23][19] + signed_kernel[2][4] ~^ image[23][20] + signed_kernel[3][0] ~^ image[24][16] + signed_kernel[3][1] ~^ image[24][17] + signed_kernel[3][2] ~^ image[24][18] + signed_kernel[3][3] ~^ image[24][19] + signed_kernel[3][4] ~^ image[24][20] + signed_kernel[4][0] ~^ image[25][16] + signed_kernel[4][1] ~^ image[25][17] + signed_kernel[4][2] ~^ image[25][18] + signed_kernel[4][3] ~^ image[25][19] + signed_kernel[4][4] ~^ image[25][20];
assign xor_sum[21][17] = signed_kernel[0][0] ~^ image[21][17] + signed_kernel[0][1] ~^ image[21][18] + signed_kernel[0][2] ~^ image[21][19] + signed_kernel[0][3] ~^ image[21][20] + signed_kernel[0][4] ~^ image[21][21] + signed_kernel[1][0] ~^ image[22][17] + signed_kernel[1][1] ~^ image[22][18] + signed_kernel[1][2] ~^ image[22][19] + signed_kernel[1][3] ~^ image[22][20] + signed_kernel[1][4] ~^ image[22][21] + signed_kernel[2][0] ~^ image[23][17] + signed_kernel[2][1] ~^ image[23][18] + signed_kernel[2][2] ~^ image[23][19] + signed_kernel[2][3] ~^ image[23][20] + signed_kernel[2][4] ~^ image[23][21] + signed_kernel[3][0] ~^ image[24][17] + signed_kernel[3][1] ~^ image[24][18] + signed_kernel[3][2] ~^ image[24][19] + signed_kernel[3][3] ~^ image[24][20] + signed_kernel[3][4] ~^ image[24][21] + signed_kernel[4][0] ~^ image[25][17] + signed_kernel[4][1] ~^ image[25][18] + signed_kernel[4][2] ~^ image[25][19] + signed_kernel[4][3] ~^ image[25][20] + signed_kernel[4][4] ~^ image[25][21];
assign xor_sum[21][18] = signed_kernel[0][0] ~^ image[21][18] + signed_kernel[0][1] ~^ image[21][19] + signed_kernel[0][2] ~^ image[21][20] + signed_kernel[0][3] ~^ image[21][21] + signed_kernel[0][4] ~^ image[21][22] + signed_kernel[1][0] ~^ image[22][18] + signed_kernel[1][1] ~^ image[22][19] + signed_kernel[1][2] ~^ image[22][20] + signed_kernel[1][3] ~^ image[22][21] + signed_kernel[1][4] ~^ image[22][22] + signed_kernel[2][0] ~^ image[23][18] + signed_kernel[2][1] ~^ image[23][19] + signed_kernel[2][2] ~^ image[23][20] + signed_kernel[2][3] ~^ image[23][21] + signed_kernel[2][4] ~^ image[23][22] + signed_kernel[3][0] ~^ image[24][18] + signed_kernel[3][1] ~^ image[24][19] + signed_kernel[3][2] ~^ image[24][20] + signed_kernel[3][3] ~^ image[24][21] + signed_kernel[3][4] ~^ image[24][22] + signed_kernel[4][0] ~^ image[25][18] + signed_kernel[4][1] ~^ image[25][19] + signed_kernel[4][2] ~^ image[25][20] + signed_kernel[4][3] ~^ image[25][21] + signed_kernel[4][4] ~^ image[25][22];
assign xor_sum[21][19] = signed_kernel[0][0] ~^ image[21][19] + signed_kernel[0][1] ~^ image[21][20] + signed_kernel[0][2] ~^ image[21][21] + signed_kernel[0][3] ~^ image[21][22] + signed_kernel[0][4] ~^ image[21][23] + signed_kernel[1][0] ~^ image[22][19] + signed_kernel[1][1] ~^ image[22][20] + signed_kernel[1][2] ~^ image[22][21] + signed_kernel[1][3] ~^ image[22][22] + signed_kernel[1][4] ~^ image[22][23] + signed_kernel[2][0] ~^ image[23][19] + signed_kernel[2][1] ~^ image[23][20] + signed_kernel[2][2] ~^ image[23][21] + signed_kernel[2][3] ~^ image[23][22] + signed_kernel[2][4] ~^ image[23][23] + signed_kernel[3][0] ~^ image[24][19] + signed_kernel[3][1] ~^ image[24][20] + signed_kernel[3][2] ~^ image[24][21] + signed_kernel[3][3] ~^ image[24][22] + signed_kernel[3][4] ~^ image[24][23] + signed_kernel[4][0] ~^ image[25][19] + signed_kernel[4][1] ~^ image[25][20] + signed_kernel[4][2] ~^ image[25][21] + signed_kernel[4][3] ~^ image[25][22] + signed_kernel[4][4] ~^ image[25][23];
assign xor_sum[21][20] = signed_kernel[0][0] ~^ image[21][20] + signed_kernel[0][1] ~^ image[21][21] + signed_kernel[0][2] ~^ image[21][22] + signed_kernel[0][3] ~^ image[21][23] + signed_kernel[0][4] ~^ image[21][24] + signed_kernel[1][0] ~^ image[22][20] + signed_kernel[1][1] ~^ image[22][21] + signed_kernel[1][2] ~^ image[22][22] + signed_kernel[1][3] ~^ image[22][23] + signed_kernel[1][4] ~^ image[22][24] + signed_kernel[2][0] ~^ image[23][20] + signed_kernel[2][1] ~^ image[23][21] + signed_kernel[2][2] ~^ image[23][22] + signed_kernel[2][3] ~^ image[23][23] + signed_kernel[2][4] ~^ image[23][24] + signed_kernel[3][0] ~^ image[24][20] + signed_kernel[3][1] ~^ image[24][21] + signed_kernel[3][2] ~^ image[24][22] + signed_kernel[3][3] ~^ image[24][23] + signed_kernel[3][4] ~^ image[24][24] + signed_kernel[4][0] ~^ image[25][20] + signed_kernel[4][1] ~^ image[25][21] + signed_kernel[4][2] ~^ image[25][22] + signed_kernel[4][3] ~^ image[25][23] + signed_kernel[4][4] ~^ image[25][24];
assign xor_sum[21][21] = signed_kernel[0][0] ~^ image[21][21] + signed_kernel[0][1] ~^ image[21][22] + signed_kernel[0][2] ~^ image[21][23] + signed_kernel[0][3] ~^ image[21][24] + signed_kernel[0][4] ~^ image[21][25] + signed_kernel[1][0] ~^ image[22][21] + signed_kernel[1][1] ~^ image[22][22] + signed_kernel[1][2] ~^ image[22][23] + signed_kernel[1][3] ~^ image[22][24] + signed_kernel[1][4] ~^ image[22][25] + signed_kernel[2][0] ~^ image[23][21] + signed_kernel[2][1] ~^ image[23][22] + signed_kernel[2][2] ~^ image[23][23] + signed_kernel[2][3] ~^ image[23][24] + signed_kernel[2][4] ~^ image[23][25] + signed_kernel[3][0] ~^ image[24][21] + signed_kernel[3][1] ~^ image[24][22] + signed_kernel[3][2] ~^ image[24][23] + signed_kernel[3][3] ~^ image[24][24] + signed_kernel[3][4] ~^ image[24][25] + signed_kernel[4][0] ~^ image[25][21] + signed_kernel[4][1] ~^ image[25][22] + signed_kernel[4][2] ~^ image[25][23] + signed_kernel[4][3] ~^ image[25][24] + signed_kernel[4][4] ~^ image[25][25];
assign xor_sum[21][22] = signed_kernel[0][0] ~^ image[21][22] + signed_kernel[0][1] ~^ image[21][23] + signed_kernel[0][2] ~^ image[21][24] + signed_kernel[0][3] ~^ image[21][25] + signed_kernel[0][4] ~^ image[21][26] + signed_kernel[1][0] ~^ image[22][22] + signed_kernel[1][1] ~^ image[22][23] + signed_kernel[1][2] ~^ image[22][24] + signed_kernel[1][3] ~^ image[22][25] + signed_kernel[1][4] ~^ image[22][26] + signed_kernel[2][0] ~^ image[23][22] + signed_kernel[2][1] ~^ image[23][23] + signed_kernel[2][2] ~^ image[23][24] + signed_kernel[2][3] ~^ image[23][25] + signed_kernel[2][4] ~^ image[23][26] + signed_kernel[3][0] ~^ image[24][22] + signed_kernel[3][1] ~^ image[24][23] + signed_kernel[3][2] ~^ image[24][24] + signed_kernel[3][3] ~^ image[24][25] + signed_kernel[3][4] ~^ image[24][26] + signed_kernel[4][0] ~^ image[25][22] + signed_kernel[4][1] ~^ image[25][23] + signed_kernel[4][2] ~^ image[25][24] + signed_kernel[4][3] ~^ image[25][25] + signed_kernel[4][4] ~^ image[25][26];
assign xor_sum[21][23] = signed_kernel[0][0] ~^ image[21][23] + signed_kernel[0][1] ~^ image[21][24] + signed_kernel[0][2] ~^ image[21][25] + signed_kernel[0][3] ~^ image[21][26] + signed_kernel[0][4] ~^ image[21][27] + signed_kernel[1][0] ~^ image[22][23] + signed_kernel[1][1] ~^ image[22][24] + signed_kernel[1][2] ~^ image[22][25] + signed_kernel[1][3] ~^ image[22][26] + signed_kernel[1][4] ~^ image[22][27] + signed_kernel[2][0] ~^ image[23][23] + signed_kernel[2][1] ~^ image[23][24] + signed_kernel[2][2] ~^ image[23][25] + signed_kernel[2][3] ~^ image[23][26] + signed_kernel[2][4] ~^ image[23][27] + signed_kernel[3][0] ~^ image[24][23] + signed_kernel[3][1] ~^ image[24][24] + signed_kernel[3][2] ~^ image[24][25] + signed_kernel[3][3] ~^ image[24][26] + signed_kernel[3][4] ~^ image[24][27] + signed_kernel[4][0] ~^ image[25][23] + signed_kernel[4][1] ~^ image[25][24] + signed_kernel[4][2] ~^ image[25][25] + signed_kernel[4][3] ~^ image[25][26] + signed_kernel[4][4] ~^ image[25][27];
assign xor_sum[22][0] = signed_kernel[0][0] ~^ image[22][0] + signed_kernel[0][1] ~^ image[22][1] + signed_kernel[0][2] ~^ image[22][2] + signed_kernel[0][3] ~^ image[22][3] + signed_kernel[0][4] ~^ image[22][4] + signed_kernel[1][0] ~^ image[23][0] + signed_kernel[1][1] ~^ image[23][1] + signed_kernel[1][2] ~^ image[23][2] + signed_kernel[1][3] ~^ image[23][3] + signed_kernel[1][4] ~^ image[23][4] + signed_kernel[2][0] ~^ image[24][0] + signed_kernel[2][1] ~^ image[24][1] + signed_kernel[2][2] ~^ image[24][2] + signed_kernel[2][3] ~^ image[24][3] + signed_kernel[2][4] ~^ image[24][4] + signed_kernel[3][0] ~^ image[25][0] + signed_kernel[3][1] ~^ image[25][1] + signed_kernel[3][2] ~^ image[25][2] + signed_kernel[3][3] ~^ image[25][3] + signed_kernel[3][4] ~^ image[25][4] + signed_kernel[4][0] ~^ image[26][0] + signed_kernel[4][1] ~^ image[26][1] + signed_kernel[4][2] ~^ image[26][2] + signed_kernel[4][3] ~^ image[26][3] + signed_kernel[4][4] ~^ image[26][4];
assign xor_sum[22][1] = signed_kernel[0][0] ~^ image[22][1] + signed_kernel[0][1] ~^ image[22][2] + signed_kernel[0][2] ~^ image[22][3] + signed_kernel[0][3] ~^ image[22][4] + signed_kernel[0][4] ~^ image[22][5] + signed_kernel[1][0] ~^ image[23][1] + signed_kernel[1][1] ~^ image[23][2] + signed_kernel[1][2] ~^ image[23][3] + signed_kernel[1][3] ~^ image[23][4] + signed_kernel[1][4] ~^ image[23][5] + signed_kernel[2][0] ~^ image[24][1] + signed_kernel[2][1] ~^ image[24][2] + signed_kernel[2][2] ~^ image[24][3] + signed_kernel[2][3] ~^ image[24][4] + signed_kernel[2][4] ~^ image[24][5] + signed_kernel[3][0] ~^ image[25][1] + signed_kernel[3][1] ~^ image[25][2] + signed_kernel[3][2] ~^ image[25][3] + signed_kernel[3][3] ~^ image[25][4] + signed_kernel[3][4] ~^ image[25][5] + signed_kernel[4][0] ~^ image[26][1] + signed_kernel[4][1] ~^ image[26][2] + signed_kernel[4][2] ~^ image[26][3] + signed_kernel[4][3] ~^ image[26][4] + signed_kernel[4][4] ~^ image[26][5];
assign xor_sum[22][2] = signed_kernel[0][0] ~^ image[22][2] + signed_kernel[0][1] ~^ image[22][3] + signed_kernel[0][2] ~^ image[22][4] + signed_kernel[0][3] ~^ image[22][5] + signed_kernel[0][4] ~^ image[22][6] + signed_kernel[1][0] ~^ image[23][2] + signed_kernel[1][1] ~^ image[23][3] + signed_kernel[1][2] ~^ image[23][4] + signed_kernel[1][3] ~^ image[23][5] + signed_kernel[1][4] ~^ image[23][6] + signed_kernel[2][0] ~^ image[24][2] + signed_kernel[2][1] ~^ image[24][3] + signed_kernel[2][2] ~^ image[24][4] + signed_kernel[2][3] ~^ image[24][5] + signed_kernel[2][4] ~^ image[24][6] + signed_kernel[3][0] ~^ image[25][2] + signed_kernel[3][1] ~^ image[25][3] + signed_kernel[3][2] ~^ image[25][4] + signed_kernel[3][3] ~^ image[25][5] + signed_kernel[3][4] ~^ image[25][6] + signed_kernel[4][0] ~^ image[26][2] + signed_kernel[4][1] ~^ image[26][3] + signed_kernel[4][2] ~^ image[26][4] + signed_kernel[4][3] ~^ image[26][5] + signed_kernel[4][4] ~^ image[26][6];
assign xor_sum[22][3] = signed_kernel[0][0] ~^ image[22][3] + signed_kernel[0][1] ~^ image[22][4] + signed_kernel[0][2] ~^ image[22][5] + signed_kernel[0][3] ~^ image[22][6] + signed_kernel[0][4] ~^ image[22][7] + signed_kernel[1][0] ~^ image[23][3] + signed_kernel[1][1] ~^ image[23][4] + signed_kernel[1][2] ~^ image[23][5] + signed_kernel[1][3] ~^ image[23][6] + signed_kernel[1][4] ~^ image[23][7] + signed_kernel[2][0] ~^ image[24][3] + signed_kernel[2][1] ~^ image[24][4] + signed_kernel[2][2] ~^ image[24][5] + signed_kernel[2][3] ~^ image[24][6] + signed_kernel[2][4] ~^ image[24][7] + signed_kernel[3][0] ~^ image[25][3] + signed_kernel[3][1] ~^ image[25][4] + signed_kernel[3][2] ~^ image[25][5] + signed_kernel[3][3] ~^ image[25][6] + signed_kernel[3][4] ~^ image[25][7] + signed_kernel[4][0] ~^ image[26][3] + signed_kernel[4][1] ~^ image[26][4] + signed_kernel[4][2] ~^ image[26][5] + signed_kernel[4][3] ~^ image[26][6] + signed_kernel[4][4] ~^ image[26][7];
assign xor_sum[22][4] = signed_kernel[0][0] ~^ image[22][4] + signed_kernel[0][1] ~^ image[22][5] + signed_kernel[0][2] ~^ image[22][6] + signed_kernel[0][3] ~^ image[22][7] + signed_kernel[0][4] ~^ image[22][8] + signed_kernel[1][0] ~^ image[23][4] + signed_kernel[1][1] ~^ image[23][5] + signed_kernel[1][2] ~^ image[23][6] + signed_kernel[1][3] ~^ image[23][7] + signed_kernel[1][4] ~^ image[23][8] + signed_kernel[2][0] ~^ image[24][4] + signed_kernel[2][1] ~^ image[24][5] + signed_kernel[2][2] ~^ image[24][6] + signed_kernel[2][3] ~^ image[24][7] + signed_kernel[2][4] ~^ image[24][8] + signed_kernel[3][0] ~^ image[25][4] + signed_kernel[3][1] ~^ image[25][5] + signed_kernel[3][2] ~^ image[25][6] + signed_kernel[3][3] ~^ image[25][7] + signed_kernel[3][4] ~^ image[25][8] + signed_kernel[4][0] ~^ image[26][4] + signed_kernel[4][1] ~^ image[26][5] + signed_kernel[4][2] ~^ image[26][6] + signed_kernel[4][3] ~^ image[26][7] + signed_kernel[4][4] ~^ image[26][8];
assign xor_sum[22][5] = signed_kernel[0][0] ~^ image[22][5] + signed_kernel[0][1] ~^ image[22][6] + signed_kernel[0][2] ~^ image[22][7] + signed_kernel[0][3] ~^ image[22][8] + signed_kernel[0][4] ~^ image[22][9] + signed_kernel[1][0] ~^ image[23][5] + signed_kernel[1][1] ~^ image[23][6] + signed_kernel[1][2] ~^ image[23][7] + signed_kernel[1][3] ~^ image[23][8] + signed_kernel[1][4] ~^ image[23][9] + signed_kernel[2][0] ~^ image[24][5] + signed_kernel[2][1] ~^ image[24][6] + signed_kernel[2][2] ~^ image[24][7] + signed_kernel[2][3] ~^ image[24][8] + signed_kernel[2][4] ~^ image[24][9] + signed_kernel[3][0] ~^ image[25][5] + signed_kernel[3][1] ~^ image[25][6] + signed_kernel[3][2] ~^ image[25][7] + signed_kernel[3][3] ~^ image[25][8] + signed_kernel[3][4] ~^ image[25][9] + signed_kernel[4][0] ~^ image[26][5] + signed_kernel[4][1] ~^ image[26][6] + signed_kernel[4][2] ~^ image[26][7] + signed_kernel[4][3] ~^ image[26][8] + signed_kernel[4][4] ~^ image[26][9];
assign xor_sum[22][6] = signed_kernel[0][0] ~^ image[22][6] + signed_kernel[0][1] ~^ image[22][7] + signed_kernel[0][2] ~^ image[22][8] + signed_kernel[0][3] ~^ image[22][9] + signed_kernel[0][4] ~^ image[22][10] + signed_kernel[1][0] ~^ image[23][6] + signed_kernel[1][1] ~^ image[23][7] + signed_kernel[1][2] ~^ image[23][8] + signed_kernel[1][3] ~^ image[23][9] + signed_kernel[1][4] ~^ image[23][10] + signed_kernel[2][0] ~^ image[24][6] + signed_kernel[2][1] ~^ image[24][7] + signed_kernel[2][2] ~^ image[24][8] + signed_kernel[2][3] ~^ image[24][9] + signed_kernel[2][4] ~^ image[24][10] + signed_kernel[3][0] ~^ image[25][6] + signed_kernel[3][1] ~^ image[25][7] + signed_kernel[3][2] ~^ image[25][8] + signed_kernel[3][3] ~^ image[25][9] + signed_kernel[3][4] ~^ image[25][10] + signed_kernel[4][0] ~^ image[26][6] + signed_kernel[4][1] ~^ image[26][7] + signed_kernel[4][2] ~^ image[26][8] + signed_kernel[4][3] ~^ image[26][9] + signed_kernel[4][4] ~^ image[26][10];
assign xor_sum[22][7] = signed_kernel[0][0] ~^ image[22][7] + signed_kernel[0][1] ~^ image[22][8] + signed_kernel[0][2] ~^ image[22][9] + signed_kernel[0][3] ~^ image[22][10] + signed_kernel[0][4] ~^ image[22][11] + signed_kernel[1][0] ~^ image[23][7] + signed_kernel[1][1] ~^ image[23][8] + signed_kernel[1][2] ~^ image[23][9] + signed_kernel[1][3] ~^ image[23][10] + signed_kernel[1][4] ~^ image[23][11] + signed_kernel[2][0] ~^ image[24][7] + signed_kernel[2][1] ~^ image[24][8] + signed_kernel[2][2] ~^ image[24][9] + signed_kernel[2][3] ~^ image[24][10] + signed_kernel[2][4] ~^ image[24][11] + signed_kernel[3][0] ~^ image[25][7] + signed_kernel[3][1] ~^ image[25][8] + signed_kernel[3][2] ~^ image[25][9] + signed_kernel[3][3] ~^ image[25][10] + signed_kernel[3][4] ~^ image[25][11] + signed_kernel[4][0] ~^ image[26][7] + signed_kernel[4][1] ~^ image[26][8] + signed_kernel[4][2] ~^ image[26][9] + signed_kernel[4][3] ~^ image[26][10] + signed_kernel[4][4] ~^ image[26][11];
assign xor_sum[22][8] = signed_kernel[0][0] ~^ image[22][8] + signed_kernel[0][1] ~^ image[22][9] + signed_kernel[0][2] ~^ image[22][10] + signed_kernel[0][3] ~^ image[22][11] + signed_kernel[0][4] ~^ image[22][12] + signed_kernel[1][0] ~^ image[23][8] + signed_kernel[1][1] ~^ image[23][9] + signed_kernel[1][2] ~^ image[23][10] + signed_kernel[1][3] ~^ image[23][11] + signed_kernel[1][4] ~^ image[23][12] + signed_kernel[2][0] ~^ image[24][8] + signed_kernel[2][1] ~^ image[24][9] + signed_kernel[2][2] ~^ image[24][10] + signed_kernel[2][3] ~^ image[24][11] + signed_kernel[2][4] ~^ image[24][12] + signed_kernel[3][0] ~^ image[25][8] + signed_kernel[3][1] ~^ image[25][9] + signed_kernel[3][2] ~^ image[25][10] + signed_kernel[3][3] ~^ image[25][11] + signed_kernel[3][4] ~^ image[25][12] + signed_kernel[4][0] ~^ image[26][8] + signed_kernel[4][1] ~^ image[26][9] + signed_kernel[4][2] ~^ image[26][10] + signed_kernel[4][3] ~^ image[26][11] + signed_kernel[4][4] ~^ image[26][12];
assign xor_sum[22][9] = signed_kernel[0][0] ~^ image[22][9] + signed_kernel[0][1] ~^ image[22][10] + signed_kernel[0][2] ~^ image[22][11] + signed_kernel[0][3] ~^ image[22][12] + signed_kernel[0][4] ~^ image[22][13] + signed_kernel[1][0] ~^ image[23][9] + signed_kernel[1][1] ~^ image[23][10] + signed_kernel[1][2] ~^ image[23][11] + signed_kernel[1][3] ~^ image[23][12] + signed_kernel[1][4] ~^ image[23][13] + signed_kernel[2][0] ~^ image[24][9] + signed_kernel[2][1] ~^ image[24][10] + signed_kernel[2][2] ~^ image[24][11] + signed_kernel[2][3] ~^ image[24][12] + signed_kernel[2][4] ~^ image[24][13] + signed_kernel[3][0] ~^ image[25][9] + signed_kernel[3][1] ~^ image[25][10] + signed_kernel[3][2] ~^ image[25][11] + signed_kernel[3][3] ~^ image[25][12] + signed_kernel[3][4] ~^ image[25][13] + signed_kernel[4][0] ~^ image[26][9] + signed_kernel[4][1] ~^ image[26][10] + signed_kernel[4][2] ~^ image[26][11] + signed_kernel[4][3] ~^ image[26][12] + signed_kernel[4][4] ~^ image[26][13];
assign xor_sum[22][10] = signed_kernel[0][0] ~^ image[22][10] + signed_kernel[0][1] ~^ image[22][11] + signed_kernel[0][2] ~^ image[22][12] + signed_kernel[0][3] ~^ image[22][13] + signed_kernel[0][4] ~^ image[22][14] + signed_kernel[1][0] ~^ image[23][10] + signed_kernel[1][1] ~^ image[23][11] + signed_kernel[1][2] ~^ image[23][12] + signed_kernel[1][3] ~^ image[23][13] + signed_kernel[1][4] ~^ image[23][14] + signed_kernel[2][0] ~^ image[24][10] + signed_kernel[2][1] ~^ image[24][11] + signed_kernel[2][2] ~^ image[24][12] + signed_kernel[2][3] ~^ image[24][13] + signed_kernel[2][4] ~^ image[24][14] + signed_kernel[3][0] ~^ image[25][10] + signed_kernel[3][1] ~^ image[25][11] + signed_kernel[3][2] ~^ image[25][12] + signed_kernel[3][3] ~^ image[25][13] + signed_kernel[3][4] ~^ image[25][14] + signed_kernel[4][0] ~^ image[26][10] + signed_kernel[4][1] ~^ image[26][11] + signed_kernel[4][2] ~^ image[26][12] + signed_kernel[4][3] ~^ image[26][13] + signed_kernel[4][4] ~^ image[26][14];
assign xor_sum[22][11] = signed_kernel[0][0] ~^ image[22][11] + signed_kernel[0][1] ~^ image[22][12] + signed_kernel[0][2] ~^ image[22][13] + signed_kernel[0][3] ~^ image[22][14] + signed_kernel[0][4] ~^ image[22][15] + signed_kernel[1][0] ~^ image[23][11] + signed_kernel[1][1] ~^ image[23][12] + signed_kernel[1][2] ~^ image[23][13] + signed_kernel[1][3] ~^ image[23][14] + signed_kernel[1][4] ~^ image[23][15] + signed_kernel[2][0] ~^ image[24][11] + signed_kernel[2][1] ~^ image[24][12] + signed_kernel[2][2] ~^ image[24][13] + signed_kernel[2][3] ~^ image[24][14] + signed_kernel[2][4] ~^ image[24][15] + signed_kernel[3][0] ~^ image[25][11] + signed_kernel[3][1] ~^ image[25][12] + signed_kernel[3][2] ~^ image[25][13] + signed_kernel[3][3] ~^ image[25][14] + signed_kernel[3][4] ~^ image[25][15] + signed_kernel[4][0] ~^ image[26][11] + signed_kernel[4][1] ~^ image[26][12] + signed_kernel[4][2] ~^ image[26][13] + signed_kernel[4][3] ~^ image[26][14] + signed_kernel[4][4] ~^ image[26][15];
assign xor_sum[22][12] = signed_kernel[0][0] ~^ image[22][12] + signed_kernel[0][1] ~^ image[22][13] + signed_kernel[0][2] ~^ image[22][14] + signed_kernel[0][3] ~^ image[22][15] + signed_kernel[0][4] ~^ image[22][16] + signed_kernel[1][0] ~^ image[23][12] + signed_kernel[1][1] ~^ image[23][13] + signed_kernel[1][2] ~^ image[23][14] + signed_kernel[1][3] ~^ image[23][15] + signed_kernel[1][4] ~^ image[23][16] + signed_kernel[2][0] ~^ image[24][12] + signed_kernel[2][1] ~^ image[24][13] + signed_kernel[2][2] ~^ image[24][14] + signed_kernel[2][3] ~^ image[24][15] + signed_kernel[2][4] ~^ image[24][16] + signed_kernel[3][0] ~^ image[25][12] + signed_kernel[3][1] ~^ image[25][13] + signed_kernel[3][2] ~^ image[25][14] + signed_kernel[3][3] ~^ image[25][15] + signed_kernel[3][4] ~^ image[25][16] + signed_kernel[4][0] ~^ image[26][12] + signed_kernel[4][1] ~^ image[26][13] + signed_kernel[4][2] ~^ image[26][14] + signed_kernel[4][3] ~^ image[26][15] + signed_kernel[4][4] ~^ image[26][16];
assign xor_sum[22][13] = signed_kernel[0][0] ~^ image[22][13] + signed_kernel[0][1] ~^ image[22][14] + signed_kernel[0][2] ~^ image[22][15] + signed_kernel[0][3] ~^ image[22][16] + signed_kernel[0][4] ~^ image[22][17] + signed_kernel[1][0] ~^ image[23][13] + signed_kernel[1][1] ~^ image[23][14] + signed_kernel[1][2] ~^ image[23][15] + signed_kernel[1][3] ~^ image[23][16] + signed_kernel[1][4] ~^ image[23][17] + signed_kernel[2][0] ~^ image[24][13] + signed_kernel[2][1] ~^ image[24][14] + signed_kernel[2][2] ~^ image[24][15] + signed_kernel[2][3] ~^ image[24][16] + signed_kernel[2][4] ~^ image[24][17] + signed_kernel[3][0] ~^ image[25][13] + signed_kernel[3][1] ~^ image[25][14] + signed_kernel[3][2] ~^ image[25][15] + signed_kernel[3][3] ~^ image[25][16] + signed_kernel[3][4] ~^ image[25][17] + signed_kernel[4][0] ~^ image[26][13] + signed_kernel[4][1] ~^ image[26][14] + signed_kernel[4][2] ~^ image[26][15] + signed_kernel[4][3] ~^ image[26][16] + signed_kernel[4][4] ~^ image[26][17];
assign xor_sum[22][14] = signed_kernel[0][0] ~^ image[22][14] + signed_kernel[0][1] ~^ image[22][15] + signed_kernel[0][2] ~^ image[22][16] + signed_kernel[0][3] ~^ image[22][17] + signed_kernel[0][4] ~^ image[22][18] + signed_kernel[1][0] ~^ image[23][14] + signed_kernel[1][1] ~^ image[23][15] + signed_kernel[1][2] ~^ image[23][16] + signed_kernel[1][3] ~^ image[23][17] + signed_kernel[1][4] ~^ image[23][18] + signed_kernel[2][0] ~^ image[24][14] + signed_kernel[2][1] ~^ image[24][15] + signed_kernel[2][2] ~^ image[24][16] + signed_kernel[2][3] ~^ image[24][17] + signed_kernel[2][4] ~^ image[24][18] + signed_kernel[3][0] ~^ image[25][14] + signed_kernel[3][1] ~^ image[25][15] + signed_kernel[3][2] ~^ image[25][16] + signed_kernel[3][3] ~^ image[25][17] + signed_kernel[3][4] ~^ image[25][18] + signed_kernel[4][0] ~^ image[26][14] + signed_kernel[4][1] ~^ image[26][15] + signed_kernel[4][2] ~^ image[26][16] + signed_kernel[4][3] ~^ image[26][17] + signed_kernel[4][4] ~^ image[26][18];
assign xor_sum[22][15] = signed_kernel[0][0] ~^ image[22][15] + signed_kernel[0][1] ~^ image[22][16] + signed_kernel[0][2] ~^ image[22][17] + signed_kernel[0][3] ~^ image[22][18] + signed_kernel[0][4] ~^ image[22][19] + signed_kernel[1][0] ~^ image[23][15] + signed_kernel[1][1] ~^ image[23][16] + signed_kernel[1][2] ~^ image[23][17] + signed_kernel[1][3] ~^ image[23][18] + signed_kernel[1][4] ~^ image[23][19] + signed_kernel[2][0] ~^ image[24][15] + signed_kernel[2][1] ~^ image[24][16] + signed_kernel[2][2] ~^ image[24][17] + signed_kernel[2][3] ~^ image[24][18] + signed_kernel[2][4] ~^ image[24][19] + signed_kernel[3][0] ~^ image[25][15] + signed_kernel[3][1] ~^ image[25][16] + signed_kernel[3][2] ~^ image[25][17] + signed_kernel[3][3] ~^ image[25][18] + signed_kernel[3][4] ~^ image[25][19] + signed_kernel[4][0] ~^ image[26][15] + signed_kernel[4][1] ~^ image[26][16] + signed_kernel[4][2] ~^ image[26][17] + signed_kernel[4][3] ~^ image[26][18] + signed_kernel[4][4] ~^ image[26][19];
assign xor_sum[22][16] = signed_kernel[0][0] ~^ image[22][16] + signed_kernel[0][1] ~^ image[22][17] + signed_kernel[0][2] ~^ image[22][18] + signed_kernel[0][3] ~^ image[22][19] + signed_kernel[0][4] ~^ image[22][20] + signed_kernel[1][0] ~^ image[23][16] + signed_kernel[1][1] ~^ image[23][17] + signed_kernel[1][2] ~^ image[23][18] + signed_kernel[1][3] ~^ image[23][19] + signed_kernel[1][4] ~^ image[23][20] + signed_kernel[2][0] ~^ image[24][16] + signed_kernel[2][1] ~^ image[24][17] + signed_kernel[2][2] ~^ image[24][18] + signed_kernel[2][3] ~^ image[24][19] + signed_kernel[2][4] ~^ image[24][20] + signed_kernel[3][0] ~^ image[25][16] + signed_kernel[3][1] ~^ image[25][17] + signed_kernel[3][2] ~^ image[25][18] + signed_kernel[3][3] ~^ image[25][19] + signed_kernel[3][4] ~^ image[25][20] + signed_kernel[4][0] ~^ image[26][16] + signed_kernel[4][1] ~^ image[26][17] + signed_kernel[4][2] ~^ image[26][18] + signed_kernel[4][3] ~^ image[26][19] + signed_kernel[4][4] ~^ image[26][20];
assign xor_sum[22][17] = signed_kernel[0][0] ~^ image[22][17] + signed_kernel[0][1] ~^ image[22][18] + signed_kernel[0][2] ~^ image[22][19] + signed_kernel[0][3] ~^ image[22][20] + signed_kernel[0][4] ~^ image[22][21] + signed_kernel[1][0] ~^ image[23][17] + signed_kernel[1][1] ~^ image[23][18] + signed_kernel[1][2] ~^ image[23][19] + signed_kernel[1][3] ~^ image[23][20] + signed_kernel[1][4] ~^ image[23][21] + signed_kernel[2][0] ~^ image[24][17] + signed_kernel[2][1] ~^ image[24][18] + signed_kernel[2][2] ~^ image[24][19] + signed_kernel[2][3] ~^ image[24][20] + signed_kernel[2][4] ~^ image[24][21] + signed_kernel[3][0] ~^ image[25][17] + signed_kernel[3][1] ~^ image[25][18] + signed_kernel[3][2] ~^ image[25][19] + signed_kernel[3][3] ~^ image[25][20] + signed_kernel[3][4] ~^ image[25][21] + signed_kernel[4][0] ~^ image[26][17] + signed_kernel[4][1] ~^ image[26][18] + signed_kernel[4][2] ~^ image[26][19] + signed_kernel[4][3] ~^ image[26][20] + signed_kernel[4][4] ~^ image[26][21];
assign xor_sum[22][18] = signed_kernel[0][0] ~^ image[22][18] + signed_kernel[0][1] ~^ image[22][19] + signed_kernel[0][2] ~^ image[22][20] + signed_kernel[0][3] ~^ image[22][21] + signed_kernel[0][4] ~^ image[22][22] + signed_kernel[1][0] ~^ image[23][18] + signed_kernel[1][1] ~^ image[23][19] + signed_kernel[1][2] ~^ image[23][20] + signed_kernel[1][3] ~^ image[23][21] + signed_kernel[1][4] ~^ image[23][22] + signed_kernel[2][0] ~^ image[24][18] + signed_kernel[2][1] ~^ image[24][19] + signed_kernel[2][2] ~^ image[24][20] + signed_kernel[2][3] ~^ image[24][21] + signed_kernel[2][4] ~^ image[24][22] + signed_kernel[3][0] ~^ image[25][18] + signed_kernel[3][1] ~^ image[25][19] + signed_kernel[3][2] ~^ image[25][20] + signed_kernel[3][3] ~^ image[25][21] + signed_kernel[3][4] ~^ image[25][22] + signed_kernel[4][0] ~^ image[26][18] + signed_kernel[4][1] ~^ image[26][19] + signed_kernel[4][2] ~^ image[26][20] + signed_kernel[4][3] ~^ image[26][21] + signed_kernel[4][4] ~^ image[26][22];
assign xor_sum[22][19] = signed_kernel[0][0] ~^ image[22][19] + signed_kernel[0][1] ~^ image[22][20] + signed_kernel[0][2] ~^ image[22][21] + signed_kernel[0][3] ~^ image[22][22] + signed_kernel[0][4] ~^ image[22][23] + signed_kernel[1][0] ~^ image[23][19] + signed_kernel[1][1] ~^ image[23][20] + signed_kernel[1][2] ~^ image[23][21] + signed_kernel[1][3] ~^ image[23][22] + signed_kernel[1][4] ~^ image[23][23] + signed_kernel[2][0] ~^ image[24][19] + signed_kernel[2][1] ~^ image[24][20] + signed_kernel[2][2] ~^ image[24][21] + signed_kernel[2][3] ~^ image[24][22] + signed_kernel[2][4] ~^ image[24][23] + signed_kernel[3][0] ~^ image[25][19] + signed_kernel[3][1] ~^ image[25][20] + signed_kernel[3][2] ~^ image[25][21] + signed_kernel[3][3] ~^ image[25][22] + signed_kernel[3][4] ~^ image[25][23] + signed_kernel[4][0] ~^ image[26][19] + signed_kernel[4][1] ~^ image[26][20] + signed_kernel[4][2] ~^ image[26][21] + signed_kernel[4][3] ~^ image[26][22] + signed_kernel[4][4] ~^ image[26][23];
assign xor_sum[22][20] = signed_kernel[0][0] ~^ image[22][20] + signed_kernel[0][1] ~^ image[22][21] + signed_kernel[0][2] ~^ image[22][22] + signed_kernel[0][3] ~^ image[22][23] + signed_kernel[0][4] ~^ image[22][24] + signed_kernel[1][0] ~^ image[23][20] + signed_kernel[1][1] ~^ image[23][21] + signed_kernel[1][2] ~^ image[23][22] + signed_kernel[1][3] ~^ image[23][23] + signed_kernel[1][4] ~^ image[23][24] + signed_kernel[2][0] ~^ image[24][20] + signed_kernel[2][1] ~^ image[24][21] + signed_kernel[2][2] ~^ image[24][22] + signed_kernel[2][3] ~^ image[24][23] + signed_kernel[2][4] ~^ image[24][24] + signed_kernel[3][0] ~^ image[25][20] + signed_kernel[3][1] ~^ image[25][21] + signed_kernel[3][2] ~^ image[25][22] + signed_kernel[3][3] ~^ image[25][23] + signed_kernel[3][4] ~^ image[25][24] + signed_kernel[4][0] ~^ image[26][20] + signed_kernel[4][1] ~^ image[26][21] + signed_kernel[4][2] ~^ image[26][22] + signed_kernel[4][3] ~^ image[26][23] + signed_kernel[4][4] ~^ image[26][24];
assign xor_sum[22][21] = signed_kernel[0][0] ~^ image[22][21] + signed_kernel[0][1] ~^ image[22][22] + signed_kernel[0][2] ~^ image[22][23] + signed_kernel[0][3] ~^ image[22][24] + signed_kernel[0][4] ~^ image[22][25] + signed_kernel[1][0] ~^ image[23][21] + signed_kernel[1][1] ~^ image[23][22] + signed_kernel[1][2] ~^ image[23][23] + signed_kernel[1][3] ~^ image[23][24] + signed_kernel[1][4] ~^ image[23][25] + signed_kernel[2][0] ~^ image[24][21] + signed_kernel[2][1] ~^ image[24][22] + signed_kernel[2][2] ~^ image[24][23] + signed_kernel[2][3] ~^ image[24][24] + signed_kernel[2][4] ~^ image[24][25] + signed_kernel[3][0] ~^ image[25][21] + signed_kernel[3][1] ~^ image[25][22] + signed_kernel[3][2] ~^ image[25][23] + signed_kernel[3][3] ~^ image[25][24] + signed_kernel[3][4] ~^ image[25][25] + signed_kernel[4][0] ~^ image[26][21] + signed_kernel[4][1] ~^ image[26][22] + signed_kernel[4][2] ~^ image[26][23] + signed_kernel[4][3] ~^ image[26][24] + signed_kernel[4][4] ~^ image[26][25];
assign xor_sum[22][22] = signed_kernel[0][0] ~^ image[22][22] + signed_kernel[0][1] ~^ image[22][23] + signed_kernel[0][2] ~^ image[22][24] + signed_kernel[0][3] ~^ image[22][25] + signed_kernel[0][4] ~^ image[22][26] + signed_kernel[1][0] ~^ image[23][22] + signed_kernel[1][1] ~^ image[23][23] + signed_kernel[1][2] ~^ image[23][24] + signed_kernel[1][3] ~^ image[23][25] + signed_kernel[1][4] ~^ image[23][26] + signed_kernel[2][0] ~^ image[24][22] + signed_kernel[2][1] ~^ image[24][23] + signed_kernel[2][2] ~^ image[24][24] + signed_kernel[2][3] ~^ image[24][25] + signed_kernel[2][4] ~^ image[24][26] + signed_kernel[3][0] ~^ image[25][22] + signed_kernel[3][1] ~^ image[25][23] + signed_kernel[3][2] ~^ image[25][24] + signed_kernel[3][3] ~^ image[25][25] + signed_kernel[3][4] ~^ image[25][26] + signed_kernel[4][0] ~^ image[26][22] + signed_kernel[4][1] ~^ image[26][23] + signed_kernel[4][2] ~^ image[26][24] + signed_kernel[4][3] ~^ image[26][25] + signed_kernel[4][4] ~^ image[26][26];
assign xor_sum[22][23] = signed_kernel[0][0] ~^ image[22][23] + signed_kernel[0][1] ~^ image[22][24] + signed_kernel[0][2] ~^ image[22][25] + signed_kernel[0][3] ~^ image[22][26] + signed_kernel[0][4] ~^ image[22][27] + signed_kernel[1][0] ~^ image[23][23] + signed_kernel[1][1] ~^ image[23][24] + signed_kernel[1][2] ~^ image[23][25] + signed_kernel[1][3] ~^ image[23][26] + signed_kernel[1][4] ~^ image[23][27] + signed_kernel[2][0] ~^ image[24][23] + signed_kernel[2][1] ~^ image[24][24] + signed_kernel[2][2] ~^ image[24][25] + signed_kernel[2][3] ~^ image[24][26] + signed_kernel[2][4] ~^ image[24][27] + signed_kernel[3][0] ~^ image[25][23] + signed_kernel[3][1] ~^ image[25][24] + signed_kernel[3][2] ~^ image[25][25] + signed_kernel[3][3] ~^ image[25][26] + signed_kernel[3][4] ~^ image[25][27] + signed_kernel[4][0] ~^ image[26][23] + signed_kernel[4][1] ~^ image[26][24] + signed_kernel[4][2] ~^ image[26][25] + signed_kernel[4][3] ~^ image[26][26] + signed_kernel[4][4] ~^ image[26][27];
assign xor_sum[23][0] = signed_kernel[0][0] ~^ image[23][0] + signed_kernel[0][1] ~^ image[23][1] + signed_kernel[0][2] ~^ image[23][2] + signed_kernel[0][3] ~^ image[23][3] + signed_kernel[0][4] ~^ image[23][4] + signed_kernel[1][0] ~^ image[24][0] + signed_kernel[1][1] ~^ image[24][1] + signed_kernel[1][2] ~^ image[24][2] + signed_kernel[1][3] ~^ image[24][3] + signed_kernel[1][4] ~^ image[24][4] + signed_kernel[2][0] ~^ image[25][0] + signed_kernel[2][1] ~^ image[25][1] + signed_kernel[2][2] ~^ image[25][2] + signed_kernel[2][3] ~^ image[25][3] + signed_kernel[2][4] ~^ image[25][4] + signed_kernel[3][0] ~^ image[26][0] + signed_kernel[3][1] ~^ image[26][1] + signed_kernel[3][2] ~^ image[26][2] + signed_kernel[3][3] ~^ image[26][3] + signed_kernel[3][4] ~^ image[26][4] + signed_kernel[4][0] ~^ image[27][0] + signed_kernel[4][1] ~^ image[27][1] + signed_kernel[4][2] ~^ image[27][2] + signed_kernel[4][3] ~^ image[27][3] + signed_kernel[4][4] ~^ image[27][4];
assign xor_sum[23][1] = signed_kernel[0][0] ~^ image[23][1] + signed_kernel[0][1] ~^ image[23][2] + signed_kernel[0][2] ~^ image[23][3] + signed_kernel[0][3] ~^ image[23][4] + signed_kernel[0][4] ~^ image[23][5] + signed_kernel[1][0] ~^ image[24][1] + signed_kernel[1][1] ~^ image[24][2] + signed_kernel[1][2] ~^ image[24][3] + signed_kernel[1][3] ~^ image[24][4] + signed_kernel[1][4] ~^ image[24][5] + signed_kernel[2][0] ~^ image[25][1] + signed_kernel[2][1] ~^ image[25][2] + signed_kernel[2][2] ~^ image[25][3] + signed_kernel[2][3] ~^ image[25][4] + signed_kernel[2][4] ~^ image[25][5] + signed_kernel[3][0] ~^ image[26][1] + signed_kernel[3][1] ~^ image[26][2] + signed_kernel[3][2] ~^ image[26][3] + signed_kernel[3][3] ~^ image[26][4] + signed_kernel[3][4] ~^ image[26][5] + signed_kernel[4][0] ~^ image[27][1] + signed_kernel[4][1] ~^ image[27][2] + signed_kernel[4][2] ~^ image[27][3] + signed_kernel[4][3] ~^ image[27][4] + signed_kernel[4][4] ~^ image[27][5];
assign xor_sum[23][2] = signed_kernel[0][0] ~^ image[23][2] + signed_kernel[0][1] ~^ image[23][3] + signed_kernel[0][2] ~^ image[23][4] + signed_kernel[0][3] ~^ image[23][5] + signed_kernel[0][4] ~^ image[23][6] + signed_kernel[1][0] ~^ image[24][2] + signed_kernel[1][1] ~^ image[24][3] + signed_kernel[1][2] ~^ image[24][4] + signed_kernel[1][3] ~^ image[24][5] + signed_kernel[1][4] ~^ image[24][6] + signed_kernel[2][0] ~^ image[25][2] + signed_kernel[2][1] ~^ image[25][3] + signed_kernel[2][2] ~^ image[25][4] + signed_kernel[2][3] ~^ image[25][5] + signed_kernel[2][4] ~^ image[25][6] + signed_kernel[3][0] ~^ image[26][2] + signed_kernel[3][1] ~^ image[26][3] + signed_kernel[3][2] ~^ image[26][4] + signed_kernel[3][3] ~^ image[26][5] + signed_kernel[3][4] ~^ image[26][6] + signed_kernel[4][0] ~^ image[27][2] + signed_kernel[4][1] ~^ image[27][3] + signed_kernel[4][2] ~^ image[27][4] + signed_kernel[4][3] ~^ image[27][5] + signed_kernel[4][4] ~^ image[27][6];
assign xor_sum[23][3] = signed_kernel[0][0] ~^ image[23][3] + signed_kernel[0][1] ~^ image[23][4] + signed_kernel[0][2] ~^ image[23][5] + signed_kernel[0][3] ~^ image[23][6] + signed_kernel[0][4] ~^ image[23][7] + signed_kernel[1][0] ~^ image[24][3] + signed_kernel[1][1] ~^ image[24][4] + signed_kernel[1][2] ~^ image[24][5] + signed_kernel[1][3] ~^ image[24][6] + signed_kernel[1][4] ~^ image[24][7] + signed_kernel[2][0] ~^ image[25][3] + signed_kernel[2][1] ~^ image[25][4] + signed_kernel[2][2] ~^ image[25][5] + signed_kernel[2][3] ~^ image[25][6] + signed_kernel[2][4] ~^ image[25][7] + signed_kernel[3][0] ~^ image[26][3] + signed_kernel[3][1] ~^ image[26][4] + signed_kernel[3][2] ~^ image[26][5] + signed_kernel[3][3] ~^ image[26][6] + signed_kernel[3][4] ~^ image[26][7] + signed_kernel[4][0] ~^ image[27][3] + signed_kernel[4][1] ~^ image[27][4] + signed_kernel[4][2] ~^ image[27][5] + signed_kernel[4][3] ~^ image[27][6] + signed_kernel[4][4] ~^ image[27][7];
assign xor_sum[23][4] = signed_kernel[0][0] ~^ image[23][4] + signed_kernel[0][1] ~^ image[23][5] + signed_kernel[0][2] ~^ image[23][6] + signed_kernel[0][3] ~^ image[23][7] + signed_kernel[0][4] ~^ image[23][8] + signed_kernel[1][0] ~^ image[24][4] + signed_kernel[1][1] ~^ image[24][5] + signed_kernel[1][2] ~^ image[24][6] + signed_kernel[1][3] ~^ image[24][7] + signed_kernel[1][4] ~^ image[24][8] + signed_kernel[2][0] ~^ image[25][4] + signed_kernel[2][1] ~^ image[25][5] + signed_kernel[2][2] ~^ image[25][6] + signed_kernel[2][3] ~^ image[25][7] + signed_kernel[2][4] ~^ image[25][8] + signed_kernel[3][0] ~^ image[26][4] + signed_kernel[3][1] ~^ image[26][5] + signed_kernel[3][2] ~^ image[26][6] + signed_kernel[3][3] ~^ image[26][7] + signed_kernel[3][4] ~^ image[26][8] + signed_kernel[4][0] ~^ image[27][4] + signed_kernel[4][1] ~^ image[27][5] + signed_kernel[4][2] ~^ image[27][6] + signed_kernel[4][3] ~^ image[27][7] + signed_kernel[4][4] ~^ image[27][8];
assign xor_sum[23][5] = signed_kernel[0][0] ~^ image[23][5] + signed_kernel[0][1] ~^ image[23][6] + signed_kernel[0][2] ~^ image[23][7] + signed_kernel[0][3] ~^ image[23][8] + signed_kernel[0][4] ~^ image[23][9] + signed_kernel[1][0] ~^ image[24][5] + signed_kernel[1][1] ~^ image[24][6] + signed_kernel[1][2] ~^ image[24][7] + signed_kernel[1][3] ~^ image[24][8] + signed_kernel[1][4] ~^ image[24][9] + signed_kernel[2][0] ~^ image[25][5] + signed_kernel[2][1] ~^ image[25][6] + signed_kernel[2][2] ~^ image[25][7] + signed_kernel[2][3] ~^ image[25][8] + signed_kernel[2][4] ~^ image[25][9] + signed_kernel[3][0] ~^ image[26][5] + signed_kernel[3][1] ~^ image[26][6] + signed_kernel[3][2] ~^ image[26][7] + signed_kernel[3][3] ~^ image[26][8] + signed_kernel[3][4] ~^ image[26][9] + signed_kernel[4][0] ~^ image[27][5] + signed_kernel[4][1] ~^ image[27][6] + signed_kernel[4][2] ~^ image[27][7] + signed_kernel[4][3] ~^ image[27][8] + signed_kernel[4][4] ~^ image[27][9];
assign xor_sum[23][6] = signed_kernel[0][0] ~^ image[23][6] + signed_kernel[0][1] ~^ image[23][7] + signed_kernel[0][2] ~^ image[23][8] + signed_kernel[0][3] ~^ image[23][9] + signed_kernel[0][4] ~^ image[23][10] + signed_kernel[1][0] ~^ image[24][6] + signed_kernel[1][1] ~^ image[24][7] + signed_kernel[1][2] ~^ image[24][8] + signed_kernel[1][3] ~^ image[24][9] + signed_kernel[1][4] ~^ image[24][10] + signed_kernel[2][0] ~^ image[25][6] + signed_kernel[2][1] ~^ image[25][7] + signed_kernel[2][2] ~^ image[25][8] + signed_kernel[2][3] ~^ image[25][9] + signed_kernel[2][4] ~^ image[25][10] + signed_kernel[3][0] ~^ image[26][6] + signed_kernel[3][1] ~^ image[26][7] + signed_kernel[3][2] ~^ image[26][8] + signed_kernel[3][3] ~^ image[26][9] + signed_kernel[3][4] ~^ image[26][10] + signed_kernel[4][0] ~^ image[27][6] + signed_kernel[4][1] ~^ image[27][7] + signed_kernel[4][2] ~^ image[27][8] + signed_kernel[4][3] ~^ image[27][9] + signed_kernel[4][4] ~^ image[27][10];
assign xor_sum[23][7] = signed_kernel[0][0] ~^ image[23][7] + signed_kernel[0][1] ~^ image[23][8] + signed_kernel[0][2] ~^ image[23][9] + signed_kernel[0][3] ~^ image[23][10] + signed_kernel[0][4] ~^ image[23][11] + signed_kernel[1][0] ~^ image[24][7] + signed_kernel[1][1] ~^ image[24][8] + signed_kernel[1][2] ~^ image[24][9] + signed_kernel[1][3] ~^ image[24][10] + signed_kernel[1][4] ~^ image[24][11] + signed_kernel[2][0] ~^ image[25][7] + signed_kernel[2][1] ~^ image[25][8] + signed_kernel[2][2] ~^ image[25][9] + signed_kernel[2][3] ~^ image[25][10] + signed_kernel[2][4] ~^ image[25][11] + signed_kernel[3][0] ~^ image[26][7] + signed_kernel[3][1] ~^ image[26][8] + signed_kernel[3][2] ~^ image[26][9] + signed_kernel[3][3] ~^ image[26][10] + signed_kernel[3][4] ~^ image[26][11] + signed_kernel[4][0] ~^ image[27][7] + signed_kernel[4][1] ~^ image[27][8] + signed_kernel[4][2] ~^ image[27][9] + signed_kernel[4][3] ~^ image[27][10] + signed_kernel[4][4] ~^ image[27][11];
assign xor_sum[23][8] = signed_kernel[0][0] ~^ image[23][8] + signed_kernel[0][1] ~^ image[23][9] + signed_kernel[0][2] ~^ image[23][10] + signed_kernel[0][3] ~^ image[23][11] + signed_kernel[0][4] ~^ image[23][12] + signed_kernel[1][0] ~^ image[24][8] + signed_kernel[1][1] ~^ image[24][9] + signed_kernel[1][2] ~^ image[24][10] + signed_kernel[1][3] ~^ image[24][11] + signed_kernel[1][4] ~^ image[24][12] + signed_kernel[2][0] ~^ image[25][8] + signed_kernel[2][1] ~^ image[25][9] + signed_kernel[2][2] ~^ image[25][10] + signed_kernel[2][3] ~^ image[25][11] + signed_kernel[2][4] ~^ image[25][12] + signed_kernel[3][0] ~^ image[26][8] + signed_kernel[3][1] ~^ image[26][9] + signed_kernel[3][2] ~^ image[26][10] + signed_kernel[3][3] ~^ image[26][11] + signed_kernel[3][4] ~^ image[26][12] + signed_kernel[4][0] ~^ image[27][8] + signed_kernel[4][1] ~^ image[27][9] + signed_kernel[4][2] ~^ image[27][10] + signed_kernel[4][3] ~^ image[27][11] + signed_kernel[4][4] ~^ image[27][12];
assign xor_sum[23][9] = signed_kernel[0][0] ~^ image[23][9] + signed_kernel[0][1] ~^ image[23][10] + signed_kernel[0][2] ~^ image[23][11] + signed_kernel[0][3] ~^ image[23][12] + signed_kernel[0][4] ~^ image[23][13] + signed_kernel[1][0] ~^ image[24][9] + signed_kernel[1][1] ~^ image[24][10] + signed_kernel[1][2] ~^ image[24][11] + signed_kernel[1][3] ~^ image[24][12] + signed_kernel[1][4] ~^ image[24][13] + signed_kernel[2][0] ~^ image[25][9] + signed_kernel[2][1] ~^ image[25][10] + signed_kernel[2][2] ~^ image[25][11] + signed_kernel[2][3] ~^ image[25][12] + signed_kernel[2][4] ~^ image[25][13] + signed_kernel[3][0] ~^ image[26][9] + signed_kernel[3][1] ~^ image[26][10] + signed_kernel[3][2] ~^ image[26][11] + signed_kernel[3][3] ~^ image[26][12] + signed_kernel[3][4] ~^ image[26][13] + signed_kernel[4][0] ~^ image[27][9] + signed_kernel[4][1] ~^ image[27][10] + signed_kernel[4][2] ~^ image[27][11] + signed_kernel[4][3] ~^ image[27][12] + signed_kernel[4][4] ~^ image[27][13];
assign xor_sum[23][10] = signed_kernel[0][0] ~^ image[23][10] + signed_kernel[0][1] ~^ image[23][11] + signed_kernel[0][2] ~^ image[23][12] + signed_kernel[0][3] ~^ image[23][13] + signed_kernel[0][4] ~^ image[23][14] + signed_kernel[1][0] ~^ image[24][10] + signed_kernel[1][1] ~^ image[24][11] + signed_kernel[1][2] ~^ image[24][12] + signed_kernel[1][3] ~^ image[24][13] + signed_kernel[1][4] ~^ image[24][14] + signed_kernel[2][0] ~^ image[25][10] + signed_kernel[2][1] ~^ image[25][11] + signed_kernel[2][2] ~^ image[25][12] + signed_kernel[2][3] ~^ image[25][13] + signed_kernel[2][4] ~^ image[25][14] + signed_kernel[3][0] ~^ image[26][10] + signed_kernel[3][1] ~^ image[26][11] + signed_kernel[3][2] ~^ image[26][12] + signed_kernel[3][3] ~^ image[26][13] + signed_kernel[3][4] ~^ image[26][14] + signed_kernel[4][0] ~^ image[27][10] + signed_kernel[4][1] ~^ image[27][11] + signed_kernel[4][2] ~^ image[27][12] + signed_kernel[4][3] ~^ image[27][13] + signed_kernel[4][4] ~^ image[27][14];
assign xor_sum[23][11] = signed_kernel[0][0] ~^ image[23][11] + signed_kernel[0][1] ~^ image[23][12] + signed_kernel[0][2] ~^ image[23][13] + signed_kernel[0][3] ~^ image[23][14] + signed_kernel[0][4] ~^ image[23][15] + signed_kernel[1][0] ~^ image[24][11] + signed_kernel[1][1] ~^ image[24][12] + signed_kernel[1][2] ~^ image[24][13] + signed_kernel[1][3] ~^ image[24][14] + signed_kernel[1][4] ~^ image[24][15] + signed_kernel[2][0] ~^ image[25][11] + signed_kernel[2][1] ~^ image[25][12] + signed_kernel[2][2] ~^ image[25][13] + signed_kernel[2][3] ~^ image[25][14] + signed_kernel[2][4] ~^ image[25][15] + signed_kernel[3][0] ~^ image[26][11] + signed_kernel[3][1] ~^ image[26][12] + signed_kernel[3][2] ~^ image[26][13] + signed_kernel[3][3] ~^ image[26][14] + signed_kernel[3][4] ~^ image[26][15] + signed_kernel[4][0] ~^ image[27][11] + signed_kernel[4][1] ~^ image[27][12] + signed_kernel[4][2] ~^ image[27][13] + signed_kernel[4][3] ~^ image[27][14] + signed_kernel[4][4] ~^ image[27][15];
assign xor_sum[23][12] = signed_kernel[0][0] ~^ image[23][12] + signed_kernel[0][1] ~^ image[23][13] + signed_kernel[0][2] ~^ image[23][14] + signed_kernel[0][3] ~^ image[23][15] + signed_kernel[0][4] ~^ image[23][16] + signed_kernel[1][0] ~^ image[24][12] + signed_kernel[1][1] ~^ image[24][13] + signed_kernel[1][2] ~^ image[24][14] + signed_kernel[1][3] ~^ image[24][15] + signed_kernel[1][4] ~^ image[24][16] + signed_kernel[2][0] ~^ image[25][12] + signed_kernel[2][1] ~^ image[25][13] + signed_kernel[2][2] ~^ image[25][14] + signed_kernel[2][3] ~^ image[25][15] + signed_kernel[2][4] ~^ image[25][16] + signed_kernel[3][0] ~^ image[26][12] + signed_kernel[3][1] ~^ image[26][13] + signed_kernel[3][2] ~^ image[26][14] + signed_kernel[3][3] ~^ image[26][15] + signed_kernel[3][4] ~^ image[26][16] + signed_kernel[4][0] ~^ image[27][12] + signed_kernel[4][1] ~^ image[27][13] + signed_kernel[4][2] ~^ image[27][14] + signed_kernel[4][3] ~^ image[27][15] + signed_kernel[4][4] ~^ image[27][16];
assign xor_sum[23][13] = signed_kernel[0][0] ~^ image[23][13] + signed_kernel[0][1] ~^ image[23][14] + signed_kernel[0][2] ~^ image[23][15] + signed_kernel[0][3] ~^ image[23][16] + signed_kernel[0][4] ~^ image[23][17] + signed_kernel[1][0] ~^ image[24][13] + signed_kernel[1][1] ~^ image[24][14] + signed_kernel[1][2] ~^ image[24][15] + signed_kernel[1][3] ~^ image[24][16] + signed_kernel[1][4] ~^ image[24][17] + signed_kernel[2][0] ~^ image[25][13] + signed_kernel[2][1] ~^ image[25][14] + signed_kernel[2][2] ~^ image[25][15] + signed_kernel[2][3] ~^ image[25][16] + signed_kernel[2][4] ~^ image[25][17] + signed_kernel[3][0] ~^ image[26][13] + signed_kernel[3][1] ~^ image[26][14] + signed_kernel[3][2] ~^ image[26][15] + signed_kernel[3][3] ~^ image[26][16] + signed_kernel[3][4] ~^ image[26][17] + signed_kernel[4][0] ~^ image[27][13] + signed_kernel[4][1] ~^ image[27][14] + signed_kernel[4][2] ~^ image[27][15] + signed_kernel[4][3] ~^ image[27][16] + signed_kernel[4][4] ~^ image[27][17];
assign xor_sum[23][14] = signed_kernel[0][0] ~^ image[23][14] + signed_kernel[0][1] ~^ image[23][15] + signed_kernel[0][2] ~^ image[23][16] + signed_kernel[0][3] ~^ image[23][17] + signed_kernel[0][4] ~^ image[23][18] + signed_kernel[1][0] ~^ image[24][14] + signed_kernel[1][1] ~^ image[24][15] + signed_kernel[1][2] ~^ image[24][16] + signed_kernel[1][3] ~^ image[24][17] + signed_kernel[1][4] ~^ image[24][18] + signed_kernel[2][0] ~^ image[25][14] + signed_kernel[2][1] ~^ image[25][15] + signed_kernel[2][2] ~^ image[25][16] + signed_kernel[2][3] ~^ image[25][17] + signed_kernel[2][4] ~^ image[25][18] + signed_kernel[3][0] ~^ image[26][14] + signed_kernel[3][1] ~^ image[26][15] + signed_kernel[3][2] ~^ image[26][16] + signed_kernel[3][3] ~^ image[26][17] + signed_kernel[3][4] ~^ image[26][18] + signed_kernel[4][0] ~^ image[27][14] + signed_kernel[4][1] ~^ image[27][15] + signed_kernel[4][2] ~^ image[27][16] + signed_kernel[4][3] ~^ image[27][17] + signed_kernel[4][4] ~^ image[27][18];
assign xor_sum[23][15] = signed_kernel[0][0] ~^ image[23][15] + signed_kernel[0][1] ~^ image[23][16] + signed_kernel[0][2] ~^ image[23][17] + signed_kernel[0][3] ~^ image[23][18] + signed_kernel[0][4] ~^ image[23][19] + signed_kernel[1][0] ~^ image[24][15] + signed_kernel[1][1] ~^ image[24][16] + signed_kernel[1][2] ~^ image[24][17] + signed_kernel[1][3] ~^ image[24][18] + signed_kernel[1][4] ~^ image[24][19] + signed_kernel[2][0] ~^ image[25][15] + signed_kernel[2][1] ~^ image[25][16] + signed_kernel[2][2] ~^ image[25][17] + signed_kernel[2][3] ~^ image[25][18] + signed_kernel[2][4] ~^ image[25][19] + signed_kernel[3][0] ~^ image[26][15] + signed_kernel[3][1] ~^ image[26][16] + signed_kernel[3][2] ~^ image[26][17] + signed_kernel[3][3] ~^ image[26][18] + signed_kernel[3][4] ~^ image[26][19] + signed_kernel[4][0] ~^ image[27][15] + signed_kernel[4][1] ~^ image[27][16] + signed_kernel[4][2] ~^ image[27][17] + signed_kernel[4][3] ~^ image[27][18] + signed_kernel[4][4] ~^ image[27][19];
assign xor_sum[23][16] = signed_kernel[0][0] ~^ image[23][16] + signed_kernel[0][1] ~^ image[23][17] + signed_kernel[0][2] ~^ image[23][18] + signed_kernel[0][3] ~^ image[23][19] + signed_kernel[0][4] ~^ image[23][20] + signed_kernel[1][0] ~^ image[24][16] + signed_kernel[1][1] ~^ image[24][17] + signed_kernel[1][2] ~^ image[24][18] + signed_kernel[1][3] ~^ image[24][19] + signed_kernel[1][4] ~^ image[24][20] + signed_kernel[2][0] ~^ image[25][16] + signed_kernel[2][1] ~^ image[25][17] + signed_kernel[2][2] ~^ image[25][18] + signed_kernel[2][3] ~^ image[25][19] + signed_kernel[2][4] ~^ image[25][20] + signed_kernel[3][0] ~^ image[26][16] + signed_kernel[3][1] ~^ image[26][17] + signed_kernel[3][2] ~^ image[26][18] + signed_kernel[3][3] ~^ image[26][19] + signed_kernel[3][4] ~^ image[26][20] + signed_kernel[4][0] ~^ image[27][16] + signed_kernel[4][1] ~^ image[27][17] + signed_kernel[4][2] ~^ image[27][18] + signed_kernel[4][3] ~^ image[27][19] + signed_kernel[4][4] ~^ image[27][20];
assign xor_sum[23][17] = signed_kernel[0][0] ~^ image[23][17] + signed_kernel[0][1] ~^ image[23][18] + signed_kernel[0][2] ~^ image[23][19] + signed_kernel[0][3] ~^ image[23][20] + signed_kernel[0][4] ~^ image[23][21] + signed_kernel[1][0] ~^ image[24][17] + signed_kernel[1][1] ~^ image[24][18] + signed_kernel[1][2] ~^ image[24][19] + signed_kernel[1][3] ~^ image[24][20] + signed_kernel[1][4] ~^ image[24][21] + signed_kernel[2][0] ~^ image[25][17] + signed_kernel[2][1] ~^ image[25][18] + signed_kernel[2][2] ~^ image[25][19] + signed_kernel[2][3] ~^ image[25][20] + signed_kernel[2][4] ~^ image[25][21] + signed_kernel[3][0] ~^ image[26][17] + signed_kernel[3][1] ~^ image[26][18] + signed_kernel[3][2] ~^ image[26][19] + signed_kernel[3][3] ~^ image[26][20] + signed_kernel[3][4] ~^ image[26][21] + signed_kernel[4][0] ~^ image[27][17] + signed_kernel[4][1] ~^ image[27][18] + signed_kernel[4][2] ~^ image[27][19] + signed_kernel[4][3] ~^ image[27][20] + signed_kernel[4][4] ~^ image[27][21];
assign xor_sum[23][18] = signed_kernel[0][0] ~^ image[23][18] + signed_kernel[0][1] ~^ image[23][19] + signed_kernel[0][2] ~^ image[23][20] + signed_kernel[0][3] ~^ image[23][21] + signed_kernel[0][4] ~^ image[23][22] + signed_kernel[1][0] ~^ image[24][18] + signed_kernel[1][1] ~^ image[24][19] + signed_kernel[1][2] ~^ image[24][20] + signed_kernel[1][3] ~^ image[24][21] + signed_kernel[1][4] ~^ image[24][22] + signed_kernel[2][0] ~^ image[25][18] + signed_kernel[2][1] ~^ image[25][19] + signed_kernel[2][2] ~^ image[25][20] + signed_kernel[2][3] ~^ image[25][21] + signed_kernel[2][4] ~^ image[25][22] + signed_kernel[3][0] ~^ image[26][18] + signed_kernel[3][1] ~^ image[26][19] + signed_kernel[3][2] ~^ image[26][20] + signed_kernel[3][3] ~^ image[26][21] + signed_kernel[3][4] ~^ image[26][22] + signed_kernel[4][0] ~^ image[27][18] + signed_kernel[4][1] ~^ image[27][19] + signed_kernel[4][2] ~^ image[27][20] + signed_kernel[4][3] ~^ image[27][21] + signed_kernel[4][4] ~^ image[27][22];
assign xor_sum[23][19] = signed_kernel[0][0] ~^ image[23][19] + signed_kernel[0][1] ~^ image[23][20] + signed_kernel[0][2] ~^ image[23][21] + signed_kernel[0][3] ~^ image[23][22] + signed_kernel[0][4] ~^ image[23][23] + signed_kernel[1][0] ~^ image[24][19] + signed_kernel[1][1] ~^ image[24][20] + signed_kernel[1][2] ~^ image[24][21] + signed_kernel[1][3] ~^ image[24][22] + signed_kernel[1][4] ~^ image[24][23] + signed_kernel[2][0] ~^ image[25][19] + signed_kernel[2][1] ~^ image[25][20] + signed_kernel[2][2] ~^ image[25][21] + signed_kernel[2][3] ~^ image[25][22] + signed_kernel[2][4] ~^ image[25][23] + signed_kernel[3][0] ~^ image[26][19] + signed_kernel[3][1] ~^ image[26][20] + signed_kernel[3][2] ~^ image[26][21] + signed_kernel[3][3] ~^ image[26][22] + signed_kernel[3][4] ~^ image[26][23] + signed_kernel[4][0] ~^ image[27][19] + signed_kernel[4][1] ~^ image[27][20] + signed_kernel[4][2] ~^ image[27][21] + signed_kernel[4][3] ~^ image[27][22] + signed_kernel[4][4] ~^ image[27][23];
assign xor_sum[23][20] = signed_kernel[0][0] ~^ image[23][20] + signed_kernel[0][1] ~^ image[23][21] + signed_kernel[0][2] ~^ image[23][22] + signed_kernel[0][3] ~^ image[23][23] + signed_kernel[0][4] ~^ image[23][24] + signed_kernel[1][0] ~^ image[24][20] + signed_kernel[1][1] ~^ image[24][21] + signed_kernel[1][2] ~^ image[24][22] + signed_kernel[1][3] ~^ image[24][23] + signed_kernel[1][4] ~^ image[24][24] + signed_kernel[2][0] ~^ image[25][20] + signed_kernel[2][1] ~^ image[25][21] + signed_kernel[2][2] ~^ image[25][22] + signed_kernel[2][3] ~^ image[25][23] + signed_kernel[2][4] ~^ image[25][24] + signed_kernel[3][0] ~^ image[26][20] + signed_kernel[3][1] ~^ image[26][21] + signed_kernel[3][2] ~^ image[26][22] + signed_kernel[3][3] ~^ image[26][23] + signed_kernel[3][4] ~^ image[26][24] + signed_kernel[4][0] ~^ image[27][20] + signed_kernel[4][1] ~^ image[27][21] + signed_kernel[4][2] ~^ image[27][22] + signed_kernel[4][3] ~^ image[27][23] + signed_kernel[4][4] ~^ image[27][24];
assign xor_sum[23][21] = signed_kernel[0][0] ~^ image[23][21] + signed_kernel[0][1] ~^ image[23][22] + signed_kernel[0][2] ~^ image[23][23] + signed_kernel[0][3] ~^ image[23][24] + signed_kernel[0][4] ~^ image[23][25] + signed_kernel[1][0] ~^ image[24][21] + signed_kernel[1][1] ~^ image[24][22] + signed_kernel[1][2] ~^ image[24][23] + signed_kernel[1][3] ~^ image[24][24] + signed_kernel[1][4] ~^ image[24][25] + signed_kernel[2][0] ~^ image[25][21] + signed_kernel[2][1] ~^ image[25][22] + signed_kernel[2][2] ~^ image[25][23] + signed_kernel[2][3] ~^ image[25][24] + signed_kernel[2][4] ~^ image[25][25] + signed_kernel[3][0] ~^ image[26][21] + signed_kernel[3][1] ~^ image[26][22] + signed_kernel[3][2] ~^ image[26][23] + signed_kernel[3][3] ~^ image[26][24] + signed_kernel[3][4] ~^ image[26][25] + signed_kernel[4][0] ~^ image[27][21] + signed_kernel[4][1] ~^ image[27][22] + signed_kernel[4][2] ~^ image[27][23] + signed_kernel[4][3] ~^ image[27][24] + signed_kernel[4][4] ~^ image[27][25];
assign xor_sum[23][22] = signed_kernel[0][0] ~^ image[23][22] + signed_kernel[0][1] ~^ image[23][23] + signed_kernel[0][2] ~^ image[23][24] + signed_kernel[0][3] ~^ image[23][25] + signed_kernel[0][4] ~^ image[23][26] + signed_kernel[1][0] ~^ image[24][22] + signed_kernel[1][1] ~^ image[24][23] + signed_kernel[1][2] ~^ image[24][24] + signed_kernel[1][3] ~^ image[24][25] + signed_kernel[1][4] ~^ image[24][26] + signed_kernel[2][0] ~^ image[25][22] + signed_kernel[2][1] ~^ image[25][23] + signed_kernel[2][2] ~^ image[25][24] + signed_kernel[2][3] ~^ image[25][25] + signed_kernel[2][4] ~^ image[25][26] + signed_kernel[3][0] ~^ image[26][22] + signed_kernel[3][1] ~^ image[26][23] + signed_kernel[3][2] ~^ image[26][24] + signed_kernel[3][3] ~^ image[26][25] + signed_kernel[3][4] ~^ image[26][26] + signed_kernel[4][0] ~^ image[27][22] + signed_kernel[4][1] ~^ image[27][23] + signed_kernel[4][2] ~^ image[27][24] + signed_kernel[4][3] ~^ image[27][25] + signed_kernel[4][4] ~^ image[27][26];
assign xor_sum[23][23] = signed_kernel[0][0] ~^ image[23][23] + signed_kernel[0][1] ~^ image[23][24] + signed_kernel[0][2] ~^ image[23][25] + signed_kernel[0][3] ~^ image[23][26] + signed_kernel[0][4] ~^ image[23][27] + signed_kernel[1][0] ~^ image[24][23] + signed_kernel[1][1] ~^ image[24][24] + signed_kernel[1][2] ~^ image[24][25] + signed_kernel[1][3] ~^ image[24][26] + signed_kernel[1][4] ~^ image[24][27] + signed_kernel[2][0] ~^ image[25][23] + signed_kernel[2][1] ~^ image[25][24] + signed_kernel[2][2] ~^ image[25][25] + signed_kernel[2][3] ~^ image[25][26] + signed_kernel[2][4] ~^ image[25][27] + signed_kernel[3][0] ~^ image[26][23] + signed_kernel[3][1] ~^ image[26][24] + signed_kernel[3][2] ~^ image[26][25] + signed_kernel[3][3] ~^ image[26][26] + signed_kernel[3][4] ~^ image[26][27] + signed_kernel[4][0] ~^ image[27][23] + signed_kernel[4][1] ~^ image[27][24] + signed_kernel[4][2] ~^ image[27][25] + signed_kernel[4][3] ~^ image[27][26] + signed_kernel[4][4] ~^ image[27][27];


 // output just the sign bit 

assign out_fmap[0][0] = xor_sum[0][0][0];
assign out_fmap[0][1] = xor_sum[0][1][0];
assign out_fmap[0][2] = xor_sum[0][2][0];
assign out_fmap[0][3] = xor_sum[0][3][0];
assign out_fmap[0][4] = xor_sum[0][4][0];
assign out_fmap[0][5] = xor_sum[0][5][0];
assign out_fmap[0][6] = xor_sum[0][6][0];
assign out_fmap[0][7] = xor_sum[0][7][0];
assign out_fmap[0][8] = xor_sum[0][8][0];
assign out_fmap[0][9] = xor_sum[0][9][0];
assign out_fmap[0][10] = xor_sum[0][10][0];
assign out_fmap[0][11] = xor_sum[0][11][0];
assign out_fmap[0][12] = xor_sum[0][12][0];
assign out_fmap[0][13] = xor_sum[0][13][0];
assign out_fmap[0][14] = xor_sum[0][14][0];
assign out_fmap[0][15] = xor_sum[0][15][0];
assign out_fmap[0][16] = xor_sum[0][16][0];
assign out_fmap[0][17] = xor_sum[0][17][0];
assign out_fmap[0][18] = xor_sum[0][18][0];
assign out_fmap[0][19] = xor_sum[0][19][0];
assign out_fmap[0][20] = xor_sum[0][20][0];
assign out_fmap[0][21] = xor_sum[0][21][0];
assign out_fmap[0][22] = xor_sum[0][22][0];
assign out_fmap[0][23] = xor_sum[0][23][0];
assign out_fmap[1][0] = xor_sum[1][0][0];
assign out_fmap[1][1] = xor_sum[1][1][0];
assign out_fmap[1][2] = xor_sum[1][2][0];
assign out_fmap[1][3] = xor_sum[1][3][0];
assign out_fmap[1][4] = xor_sum[1][4][0];
assign out_fmap[1][5] = xor_sum[1][5][0];
assign out_fmap[1][6] = xor_sum[1][6][0];
assign out_fmap[1][7] = xor_sum[1][7][0];
assign out_fmap[1][8] = xor_sum[1][8][0];
assign out_fmap[1][9] = xor_sum[1][9][0];
assign out_fmap[1][10] = xor_sum[1][10][0];
assign out_fmap[1][11] = xor_sum[1][11][0];
assign out_fmap[1][12] = xor_sum[1][12][0];
assign out_fmap[1][13] = xor_sum[1][13][0];
assign out_fmap[1][14] = xor_sum[1][14][0];
assign out_fmap[1][15] = xor_sum[1][15][0];
assign out_fmap[1][16] = xor_sum[1][16][0];
assign out_fmap[1][17] = xor_sum[1][17][0];
assign out_fmap[1][18] = xor_sum[1][18][0];
assign out_fmap[1][19] = xor_sum[1][19][0];
assign out_fmap[1][20] = xor_sum[1][20][0];
assign out_fmap[1][21] = xor_sum[1][21][0];
assign out_fmap[1][22] = xor_sum[1][22][0];
assign out_fmap[1][23] = xor_sum[1][23][0];
assign out_fmap[2][0] = xor_sum[2][0][0];
assign out_fmap[2][1] = xor_sum[2][1][0];
assign out_fmap[2][2] = xor_sum[2][2][0];
assign out_fmap[2][3] = xor_sum[2][3][0];
assign out_fmap[2][4] = xor_sum[2][4][0];
assign out_fmap[2][5] = xor_sum[2][5][0];
assign out_fmap[2][6] = xor_sum[2][6][0];
assign out_fmap[2][7] = xor_sum[2][7][0];
assign out_fmap[2][8] = xor_sum[2][8][0];
assign out_fmap[2][9] = xor_sum[2][9][0];
assign out_fmap[2][10] = xor_sum[2][10][0];
assign out_fmap[2][11] = xor_sum[2][11][0];
assign out_fmap[2][12] = xor_sum[2][12][0];
assign out_fmap[2][13] = xor_sum[2][13][0];
assign out_fmap[2][14] = xor_sum[2][14][0];
assign out_fmap[2][15] = xor_sum[2][15][0];
assign out_fmap[2][16] = xor_sum[2][16][0];
assign out_fmap[2][17] = xor_sum[2][17][0];
assign out_fmap[2][18] = xor_sum[2][18][0];
assign out_fmap[2][19] = xor_sum[2][19][0];
assign out_fmap[2][20] = xor_sum[2][20][0];
assign out_fmap[2][21] = xor_sum[2][21][0];
assign out_fmap[2][22] = xor_sum[2][22][0];
assign out_fmap[2][23] = xor_sum[2][23][0];
assign out_fmap[3][0] = xor_sum[3][0][0];
assign out_fmap[3][1] = xor_sum[3][1][0];
assign out_fmap[3][2] = xor_sum[3][2][0];
assign out_fmap[3][3] = xor_sum[3][3][0];
assign out_fmap[3][4] = xor_sum[3][4][0];
assign out_fmap[3][5] = xor_sum[3][5][0];
assign out_fmap[3][6] = xor_sum[3][6][0];
assign out_fmap[3][7] = xor_sum[3][7][0];
assign out_fmap[3][8] = xor_sum[3][8][0];
assign out_fmap[3][9] = xor_sum[3][9][0];
assign out_fmap[3][10] = xor_sum[3][10][0];
assign out_fmap[3][11] = xor_sum[3][11][0];
assign out_fmap[3][12] = xor_sum[3][12][0];
assign out_fmap[3][13] = xor_sum[3][13][0];
assign out_fmap[3][14] = xor_sum[3][14][0];
assign out_fmap[3][15] = xor_sum[3][15][0];
assign out_fmap[3][16] = xor_sum[3][16][0];
assign out_fmap[3][17] = xor_sum[3][17][0];
assign out_fmap[3][18] = xor_sum[3][18][0];
assign out_fmap[3][19] = xor_sum[3][19][0];
assign out_fmap[3][20] = xor_sum[3][20][0];
assign out_fmap[3][21] = xor_sum[3][21][0];
assign out_fmap[3][22] = xor_sum[3][22][0];
assign out_fmap[3][23] = xor_sum[3][23][0];
assign out_fmap[4][0] = xor_sum[4][0][0];
assign out_fmap[4][1] = xor_sum[4][1][0];
assign out_fmap[4][2] = xor_sum[4][2][0];
assign out_fmap[4][3] = xor_sum[4][3][0];
assign out_fmap[4][4] = xor_sum[4][4][0];
assign out_fmap[4][5] = xor_sum[4][5][0];
assign out_fmap[4][6] = xor_sum[4][6][0];
assign out_fmap[4][7] = xor_sum[4][7][0];
assign out_fmap[4][8] = xor_sum[4][8][0];
assign out_fmap[4][9] = xor_sum[4][9][0];
assign out_fmap[4][10] = xor_sum[4][10][0];
assign out_fmap[4][11] = xor_sum[4][11][0];
assign out_fmap[4][12] = xor_sum[4][12][0];
assign out_fmap[4][13] = xor_sum[4][13][0];
assign out_fmap[4][14] = xor_sum[4][14][0];
assign out_fmap[4][15] = xor_sum[4][15][0];
assign out_fmap[4][16] = xor_sum[4][16][0];
assign out_fmap[4][17] = xor_sum[4][17][0];
assign out_fmap[4][18] = xor_sum[4][18][0];
assign out_fmap[4][19] = xor_sum[4][19][0];
assign out_fmap[4][20] = xor_sum[4][20][0];
assign out_fmap[4][21] = xor_sum[4][21][0];
assign out_fmap[4][22] = xor_sum[4][22][0];
assign out_fmap[4][23] = xor_sum[4][23][0];
assign out_fmap[5][0] = xor_sum[5][0][0];
assign out_fmap[5][1] = xor_sum[5][1][0];
assign out_fmap[5][2] = xor_sum[5][2][0];
assign out_fmap[5][3] = xor_sum[5][3][0];
assign out_fmap[5][4] = xor_sum[5][4][0];
assign out_fmap[5][5] = xor_sum[5][5][0];
assign out_fmap[5][6] = xor_sum[5][6][0];
assign out_fmap[5][7] = xor_sum[5][7][0];
assign out_fmap[5][8] = xor_sum[5][8][0];
assign out_fmap[5][9] = xor_sum[5][9][0];
assign out_fmap[5][10] = xor_sum[5][10][0];
assign out_fmap[5][11] = xor_sum[5][11][0];
assign out_fmap[5][12] = xor_sum[5][12][0];
assign out_fmap[5][13] = xor_sum[5][13][0];
assign out_fmap[5][14] = xor_sum[5][14][0];
assign out_fmap[5][15] = xor_sum[5][15][0];
assign out_fmap[5][16] = xor_sum[5][16][0];
assign out_fmap[5][17] = xor_sum[5][17][0];
assign out_fmap[5][18] = xor_sum[5][18][0];
assign out_fmap[5][19] = xor_sum[5][19][0];
assign out_fmap[5][20] = xor_sum[5][20][0];
assign out_fmap[5][21] = xor_sum[5][21][0];
assign out_fmap[5][22] = xor_sum[5][22][0];
assign out_fmap[5][23] = xor_sum[5][23][0];
assign out_fmap[6][0] = xor_sum[6][0][0];
assign out_fmap[6][1] = xor_sum[6][1][0];
assign out_fmap[6][2] = xor_sum[6][2][0];
assign out_fmap[6][3] = xor_sum[6][3][0];
assign out_fmap[6][4] = xor_sum[6][4][0];
assign out_fmap[6][5] = xor_sum[6][5][0];
assign out_fmap[6][6] = xor_sum[6][6][0];
assign out_fmap[6][7] = xor_sum[6][7][0];
assign out_fmap[6][8] = xor_sum[6][8][0];
assign out_fmap[6][9] = xor_sum[6][9][0];
assign out_fmap[6][10] = xor_sum[6][10][0];
assign out_fmap[6][11] = xor_sum[6][11][0];
assign out_fmap[6][12] = xor_sum[6][12][0];
assign out_fmap[6][13] = xor_sum[6][13][0];
assign out_fmap[6][14] = xor_sum[6][14][0];
assign out_fmap[6][15] = xor_sum[6][15][0];
assign out_fmap[6][16] = xor_sum[6][16][0];
assign out_fmap[6][17] = xor_sum[6][17][0];
assign out_fmap[6][18] = xor_sum[6][18][0];
assign out_fmap[6][19] = xor_sum[6][19][0];
assign out_fmap[6][20] = xor_sum[6][20][0];
assign out_fmap[6][21] = xor_sum[6][21][0];
assign out_fmap[6][22] = xor_sum[6][22][0];
assign out_fmap[6][23] = xor_sum[6][23][0];
assign out_fmap[7][0] = xor_sum[7][0][0];
assign out_fmap[7][1] = xor_sum[7][1][0];
assign out_fmap[7][2] = xor_sum[7][2][0];
assign out_fmap[7][3] = xor_sum[7][3][0];
assign out_fmap[7][4] = xor_sum[7][4][0];
assign out_fmap[7][5] = xor_sum[7][5][0];
assign out_fmap[7][6] = xor_sum[7][6][0];
assign out_fmap[7][7] = xor_sum[7][7][0];
assign out_fmap[7][8] = xor_sum[7][8][0];
assign out_fmap[7][9] = xor_sum[7][9][0];
assign out_fmap[7][10] = xor_sum[7][10][0];
assign out_fmap[7][11] = xor_sum[7][11][0];
assign out_fmap[7][12] = xor_sum[7][12][0];
assign out_fmap[7][13] = xor_sum[7][13][0];
assign out_fmap[7][14] = xor_sum[7][14][0];
assign out_fmap[7][15] = xor_sum[7][15][0];
assign out_fmap[7][16] = xor_sum[7][16][0];
assign out_fmap[7][17] = xor_sum[7][17][0];
assign out_fmap[7][18] = xor_sum[7][18][0];
assign out_fmap[7][19] = xor_sum[7][19][0];
assign out_fmap[7][20] = xor_sum[7][20][0];
assign out_fmap[7][21] = xor_sum[7][21][0];
assign out_fmap[7][22] = xor_sum[7][22][0];
assign out_fmap[7][23] = xor_sum[7][23][0];
assign out_fmap[8][0] = xor_sum[8][0][0];
assign out_fmap[8][1] = xor_sum[8][1][0];
assign out_fmap[8][2] = xor_sum[8][2][0];
assign out_fmap[8][3] = xor_sum[8][3][0];
assign out_fmap[8][4] = xor_sum[8][4][0];
assign out_fmap[8][5] = xor_sum[8][5][0];
assign out_fmap[8][6] = xor_sum[8][6][0];
assign out_fmap[8][7] = xor_sum[8][7][0];
assign out_fmap[8][8] = xor_sum[8][8][0];
assign out_fmap[8][9] = xor_sum[8][9][0];
assign out_fmap[8][10] = xor_sum[8][10][0];
assign out_fmap[8][11] = xor_sum[8][11][0];
assign out_fmap[8][12] = xor_sum[8][12][0];
assign out_fmap[8][13] = xor_sum[8][13][0];
assign out_fmap[8][14] = xor_sum[8][14][0];
assign out_fmap[8][15] = xor_sum[8][15][0];
assign out_fmap[8][16] = xor_sum[8][16][0];
assign out_fmap[8][17] = xor_sum[8][17][0];
assign out_fmap[8][18] = xor_sum[8][18][0];
assign out_fmap[8][19] = xor_sum[8][19][0];
assign out_fmap[8][20] = xor_sum[8][20][0];
assign out_fmap[8][21] = xor_sum[8][21][0];
assign out_fmap[8][22] = xor_sum[8][22][0];
assign out_fmap[8][23] = xor_sum[8][23][0];
assign out_fmap[9][0] = xor_sum[9][0][0];
assign out_fmap[9][1] = xor_sum[9][1][0];
assign out_fmap[9][2] = xor_sum[9][2][0];
assign out_fmap[9][3] = xor_sum[9][3][0];
assign out_fmap[9][4] = xor_sum[9][4][0];
assign out_fmap[9][5] = xor_sum[9][5][0];
assign out_fmap[9][6] = xor_sum[9][6][0];
assign out_fmap[9][7] = xor_sum[9][7][0];
assign out_fmap[9][8] = xor_sum[9][8][0];
assign out_fmap[9][9] = xor_sum[9][9][0];
assign out_fmap[9][10] = xor_sum[9][10][0];
assign out_fmap[9][11] = xor_sum[9][11][0];
assign out_fmap[9][12] = xor_sum[9][12][0];
assign out_fmap[9][13] = xor_sum[9][13][0];
assign out_fmap[9][14] = xor_sum[9][14][0];
assign out_fmap[9][15] = xor_sum[9][15][0];
assign out_fmap[9][16] = xor_sum[9][16][0];
assign out_fmap[9][17] = xor_sum[9][17][0];
assign out_fmap[9][18] = xor_sum[9][18][0];
assign out_fmap[9][19] = xor_sum[9][19][0];
assign out_fmap[9][20] = xor_sum[9][20][0];
assign out_fmap[9][21] = xor_sum[9][21][0];
assign out_fmap[9][22] = xor_sum[9][22][0];
assign out_fmap[9][23] = xor_sum[9][23][0];
assign out_fmap[10][0] = xor_sum[10][0][0];
assign out_fmap[10][1] = xor_sum[10][1][0];
assign out_fmap[10][2] = xor_sum[10][2][0];
assign out_fmap[10][3] = xor_sum[10][3][0];
assign out_fmap[10][4] = xor_sum[10][4][0];
assign out_fmap[10][5] = xor_sum[10][5][0];
assign out_fmap[10][6] = xor_sum[10][6][0];
assign out_fmap[10][7] = xor_sum[10][7][0];
assign out_fmap[10][8] = xor_sum[10][8][0];
assign out_fmap[10][9] = xor_sum[10][9][0];
assign out_fmap[10][10] = xor_sum[10][10][0];
assign out_fmap[10][11] = xor_sum[10][11][0];
assign out_fmap[10][12] = xor_sum[10][12][0];
assign out_fmap[10][13] = xor_sum[10][13][0];
assign out_fmap[10][14] = xor_sum[10][14][0];
assign out_fmap[10][15] = xor_sum[10][15][0];
assign out_fmap[10][16] = xor_sum[10][16][0];
assign out_fmap[10][17] = xor_sum[10][17][0];
assign out_fmap[10][18] = xor_sum[10][18][0];
assign out_fmap[10][19] = xor_sum[10][19][0];
assign out_fmap[10][20] = xor_sum[10][20][0];
assign out_fmap[10][21] = xor_sum[10][21][0];
assign out_fmap[10][22] = xor_sum[10][22][0];
assign out_fmap[10][23] = xor_sum[10][23][0];
assign out_fmap[11][0] = xor_sum[11][0][0];
assign out_fmap[11][1] = xor_sum[11][1][0];
assign out_fmap[11][2] = xor_sum[11][2][0];
assign out_fmap[11][3] = xor_sum[11][3][0];
assign out_fmap[11][4] = xor_sum[11][4][0];
assign out_fmap[11][5] = xor_sum[11][5][0];
assign out_fmap[11][6] = xor_sum[11][6][0];
assign out_fmap[11][7] = xor_sum[11][7][0];
assign out_fmap[11][8] = xor_sum[11][8][0];
assign out_fmap[11][9] = xor_sum[11][9][0];
assign out_fmap[11][10] = xor_sum[11][10][0];
assign out_fmap[11][11] = xor_sum[11][11][0];
assign out_fmap[11][12] = xor_sum[11][12][0];
assign out_fmap[11][13] = xor_sum[11][13][0];
assign out_fmap[11][14] = xor_sum[11][14][0];
assign out_fmap[11][15] = xor_sum[11][15][0];
assign out_fmap[11][16] = xor_sum[11][16][0];
assign out_fmap[11][17] = xor_sum[11][17][0];
assign out_fmap[11][18] = xor_sum[11][18][0];
assign out_fmap[11][19] = xor_sum[11][19][0];
assign out_fmap[11][20] = xor_sum[11][20][0];
assign out_fmap[11][21] = xor_sum[11][21][0];
assign out_fmap[11][22] = xor_sum[11][22][0];
assign out_fmap[11][23] = xor_sum[11][23][0];
assign out_fmap[12][0] = xor_sum[12][0][0];
assign out_fmap[12][1] = xor_sum[12][1][0];
assign out_fmap[12][2] = xor_sum[12][2][0];
assign out_fmap[12][3] = xor_sum[12][3][0];
assign out_fmap[12][4] = xor_sum[12][4][0];
assign out_fmap[12][5] = xor_sum[12][5][0];
assign out_fmap[12][6] = xor_sum[12][6][0];
assign out_fmap[12][7] = xor_sum[12][7][0];
assign out_fmap[12][8] = xor_sum[12][8][0];
assign out_fmap[12][9] = xor_sum[12][9][0];
assign out_fmap[12][10] = xor_sum[12][10][0];
assign out_fmap[12][11] = xor_sum[12][11][0];
assign out_fmap[12][12] = xor_sum[12][12][0];
assign out_fmap[12][13] = xor_sum[12][13][0];
assign out_fmap[12][14] = xor_sum[12][14][0];
assign out_fmap[12][15] = xor_sum[12][15][0];
assign out_fmap[12][16] = xor_sum[12][16][0];
assign out_fmap[12][17] = xor_sum[12][17][0];
assign out_fmap[12][18] = xor_sum[12][18][0];
assign out_fmap[12][19] = xor_sum[12][19][0];
assign out_fmap[12][20] = xor_sum[12][20][0];
assign out_fmap[12][21] = xor_sum[12][21][0];
assign out_fmap[12][22] = xor_sum[12][22][0];
assign out_fmap[12][23] = xor_sum[12][23][0];
assign out_fmap[13][0] = xor_sum[13][0][0];
assign out_fmap[13][1] = xor_sum[13][1][0];
assign out_fmap[13][2] = xor_sum[13][2][0];
assign out_fmap[13][3] = xor_sum[13][3][0];
assign out_fmap[13][4] = xor_sum[13][4][0];
assign out_fmap[13][5] = xor_sum[13][5][0];
assign out_fmap[13][6] = xor_sum[13][6][0];
assign out_fmap[13][7] = xor_sum[13][7][0];
assign out_fmap[13][8] = xor_sum[13][8][0];
assign out_fmap[13][9] = xor_sum[13][9][0];
assign out_fmap[13][10] = xor_sum[13][10][0];
assign out_fmap[13][11] = xor_sum[13][11][0];
assign out_fmap[13][12] = xor_sum[13][12][0];
assign out_fmap[13][13] = xor_sum[13][13][0];
assign out_fmap[13][14] = xor_sum[13][14][0];
assign out_fmap[13][15] = xor_sum[13][15][0];
assign out_fmap[13][16] = xor_sum[13][16][0];
assign out_fmap[13][17] = xor_sum[13][17][0];
assign out_fmap[13][18] = xor_sum[13][18][0];
assign out_fmap[13][19] = xor_sum[13][19][0];
assign out_fmap[13][20] = xor_sum[13][20][0];
assign out_fmap[13][21] = xor_sum[13][21][0];
assign out_fmap[13][22] = xor_sum[13][22][0];
assign out_fmap[13][23] = xor_sum[13][23][0];
assign out_fmap[14][0] = xor_sum[14][0][0];
assign out_fmap[14][1] = xor_sum[14][1][0];
assign out_fmap[14][2] = xor_sum[14][2][0];
assign out_fmap[14][3] = xor_sum[14][3][0];
assign out_fmap[14][4] = xor_sum[14][4][0];
assign out_fmap[14][5] = xor_sum[14][5][0];
assign out_fmap[14][6] = xor_sum[14][6][0];
assign out_fmap[14][7] = xor_sum[14][7][0];
assign out_fmap[14][8] = xor_sum[14][8][0];
assign out_fmap[14][9] = xor_sum[14][9][0];
assign out_fmap[14][10] = xor_sum[14][10][0];
assign out_fmap[14][11] = xor_sum[14][11][0];
assign out_fmap[14][12] = xor_sum[14][12][0];
assign out_fmap[14][13] = xor_sum[14][13][0];
assign out_fmap[14][14] = xor_sum[14][14][0];
assign out_fmap[14][15] = xor_sum[14][15][0];
assign out_fmap[14][16] = xor_sum[14][16][0];
assign out_fmap[14][17] = xor_sum[14][17][0];
assign out_fmap[14][18] = xor_sum[14][18][0];
assign out_fmap[14][19] = xor_sum[14][19][0];
assign out_fmap[14][20] = xor_sum[14][20][0];
assign out_fmap[14][21] = xor_sum[14][21][0];
assign out_fmap[14][22] = xor_sum[14][22][0];
assign out_fmap[14][23] = xor_sum[14][23][0];
assign out_fmap[15][0] = xor_sum[15][0][0];
assign out_fmap[15][1] = xor_sum[15][1][0];
assign out_fmap[15][2] = xor_sum[15][2][0];
assign out_fmap[15][3] = xor_sum[15][3][0];
assign out_fmap[15][4] = xor_sum[15][4][0];
assign out_fmap[15][5] = xor_sum[15][5][0];
assign out_fmap[15][6] = xor_sum[15][6][0];
assign out_fmap[15][7] = xor_sum[15][7][0];
assign out_fmap[15][8] = xor_sum[15][8][0];
assign out_fmap[15][9] = xor_sum[15][9][0];
assign out_fmap[15][10] = xor_sum[15][10][0];
assign out_fmap[15][11] = xor_sum[15][11][0];
assign out_fmap[15][12] = xor_sum[15][12][0];
assign out_fmap[15][13] = xor_sum[15][13][0];
assign out_fmap[15][14] = xor_sum[15][14][0];
assign out_fmap[15][15] = xor_sum[15][15][0];
assign out_fmap[15][16] = xor_sum[15][16][0];
assign out_fmap[15][17] = xor_sum[15][17][0];
assign out_fmap[15][18] = xor_sum[15][18][0];
assign out_fmap[15][19] = xor_sum[15][19][0];
assign out_fmap[15][20] = xor_sum[15][20][0];
assign out_fmap[15][21] = xor_sum[15][21][0];
assign out_fmap[15][22] = xor_sum[15][22][0];
assign out_fmap[15][23] = xor_sum[15][23][0];
assign out_fmap[16][0] = xor_sum[16][0][0];
assign out_fmap[16][1] = xor_sum[16][1][0];
assign out_fmap[16][2] = xor_sum[16][2][0];
assign out_fmap[16][3] = xor_sum[16][3][0];
assign out_fmap[16][4] = xor_sum[16][4][0];
assign out_fmap[16][5] = xor_sum[16][5][0];
assign out_fmap[16][6] = xor_sum[16][6][0];
assign out_fmap[16][7] = xor_sum[16][7][0];
assign out_fmap[16][8] = xor_sum[16][8][0];
assign out_fmap[16][9] = xor_sum[16][9][0];
assign out_fmap[16][10] = xor_sum[16][10][0];
assign out_fmap[16][11] = xor_sum[16][11][0];
assign out_fmap[16][12] = xor_sum[16][12][0];
assign out_fmap[16][13] = xor_sum[16][13][0];
assign out_fmap[16][14] = xor_sum[16][14][0];
assign out_fmap[16][15] = xor_sum[16][15][0];
assign out_fmap[16][16] = xor_sum[16][16][0];
assign out_fmap[16][17] = xor_sum[16][17][0];
assign out_fmap[16][18] = xor_sum[16][18][0];
assign out_fmap[16][19] = xor_sum[16][19][0];
assign out_fmap[16][20] = xor_sum[16][20][0];
assign out_fmap[16][21] = xor_sum[16][21][0];
assign out_fmap[16][22] = xor_sum[16][22][0];
assign out_fmap[16][23] = xor_sum[16][23][0];
assign out_fmap[17][0] = xor_sum[17][0][0];
assign out_fmap[17][1] = xor_sum[17][1][0];
assign out_fmap[17][2] = xor_sum[17][2][0];
assign out_fmap[17][3] = xor_sum[17][3][0];
assign out_fmap[17][4] = xor_sum[17][4][0];
assign out_fmap[17][5] = xor_sum[17][5][0];
assign out_fmap[17][6] = xor_sum[17][6][0];
assign out_fmap[17][7] = xor_sum[17][7][0];
assign out_fmap[17][8] = xor_sum[17][8][0];
assign out_fmap[17][9] = xor_sum[17][9][0];
assign out_fmap[17][10] = xor_sum[17][10][0];
assign out_fmap[17][11] = xor_sum[17][11][0];
assign out_fmap[17][12] = xor_sum[17][12][0];
assign out_fmap[17][13] = xor_sum[17][13][0];
assign out_fmap[17][14] = xor_sum[17][14][0];
assign out_fmap[17][15] = xor_sum[17][15][0];
assign out_fmap[17][16] = xor_sum[17][16][0];
assign out_fmap[17][17] = xor_sum[17][17][0];
assign out_fmap[17][18] = xor_sum[17][18][0];
assign out_fmap[17][19] = xor_sum[17][19][0];
assign out_fmap[17][20] = xor_sum[17][20][0];
assign out_fmap[17][21] = xor_sum[17][21][0];
assign out_fmap[17][22] = xor_sum[17][22][0];
assign out_fmap[17][23] = xor_sum[17][23][0];
assign out_fmap[18][0] = xor_sum[18][0][0];
assign out_fmap[18][1] = xor_sum[18][1][0];
assign out_fmap[18][2] = xor_sum[18][2][0];
assign out_fmap[18][3] = xor_sum[18][3][0];
assign out_fmap[18][4] = xor_sum[18][4][0];
assign out_fmap[18][5] = xor_sum[18][5][0];
assign out_fmap[18][6] = xor_sum[18][6][0];
assign out_fmap[18][7] = xor_sum[18][7][0];
assign out_fmap[18][8] = xor_sum[18][8][0];
assign out_fmap[18][9] = xor_sum[18][9][0];
assign out_fmap[18][10] = xor_sum[18][10][0];
assign out_fmap[18][11] = xor_sum[18][11][0];
assign out_fmap[18][12] = xor_sum[18][12][0];
assign out_fmap[18][13] = xor_sum[18][13][0];
assign out_fmap[18][14] = xor_sum[18][14][0];
assign out_fmap[18][15] = xor_sum[18][15][0];
assign out_fmap[18][16] = xor_sum[18][16][0];
assign out_fmap[18][17] = xor_sum[18][17][0];
assign out_fmap[18][18] = xor_sum[18][18][0];
assign out_fmap[18][19] = xor_sum[18][19][0];
assign out_fmap[18][20] = xor_sum[18][20][0];
assign out_fmap[18][21] = xor_sum[18][21][0];
assign out_fmap[18][22] = xor_sum[18][22][0];
assign out_fmap[18][23] = xor_sum[18][23][0];
assign out_fmap[19][0] = xor_sum[19][0][0];
assign out_fmap[19][1] = xor_sum[19][1][0];
assign out_fmap[19][2] = xor_sum[19][2][0];
assign out_fmap[19][3] = xor_sum[19][3][0];
assign out_fmap[19][4] = xor_sum[19][4][0];
assign out_fmap[19][5] = xor_sum[19][5][0];
assign out_fmap[19][6] = xor_sum[19][6][0];
assign out_fmap[19][7] = xor_sum[19][7][0];
assign out_fmap[19][8] = xor_sum[19][8][0];
assign out_fmap[19][9] = xor_sum[19][9][0];
assign out_fmap[19][10] = xor_sum[19][10][0];
assign out_fmap[19][11] = xor_sum[19][11][0];
assign out_fmap[19][12] = xor_sum[19][12][0];
assign out_fmap[19][13] = xor_sum[19][13][0];
assign out_fmap[19][14] = xor_sum[19][14][0];
assign out_fmap[19][15] = xor_sum[19][15][0];
assign out_fmap[19][16] = xor_sum[19][16][0];
assign out_fmap[19][17] = xor_sum[19][17][0];
assign out_fmap[19][18] = xor_sum[19][18][0];
assign out_fmap[19][19] = xor_sum[19][19][0];
assign out_fmap[19][20] = xor_sum[19][20][0];
assign out_fmap[19][21] = xor_sum[19][21][0];
assign out_fmap[19][22] = xor_sum[19][22][0];
assign out_fmap[19][23] = xor_sum[19][23][0];
assign out_fmap[20][0] = xor_sum[20][0][0];
assign out_fmap[20][1] = xor_sum[20][1][0];
assign out_fmap[20][2] = xor_sum[20][2][0];
assign out_fmap[20][3] = xor_sum[20][3][0];
assign out_fmap[20][4] = xor_sum[20][4][0];
assign out_fmap[20][5] = xor_sum[20][5][0];
assign out_fmap[20][6] = xor_sum[20][6][0];
assign out_fmap[20][7] = xor_sum[20][7][0];
assign out_fmap[20][8] = xor_sum[20][8][0];
assign out_fmap[20][9] = xor_sum[20][9][0];
assign out_fmap[20][10] = xor_sum[20][10][0];
assign out_fmap[20][11] = xor_sum[20][11][0];
assign out_fmap[20][12] = xor_sum[20][12][0];
assign out_fmap[20][13] = xor_sum[20][13][0];
assign out_fmap[20][14] = xor_sum[20][14][0];
assign out_fmap[20][15] = xor_sum[20][15][0];
assign out_fmap[20][16] = xor_sum[20][16][0];
assign out_fmap[20][17] = xor_sum[20][17][0];
assign out_fmap[20][18] = xor_sum[20][18][0];
assign out_fmap[20][19] = xor_sum[20][19][0];
assign out_fmap[20][20] = xor_sum[20][20][0];
assign out_fmap[20][21] = xor_sum[20][21][0];
assign out_fmap[20][22] = xor_sum[20][22][0];
assign out_fmap[20][23] = xor_sum[20][23][0];
assign out_fmap[21][0] = xor_sum[21][0][0];
assign out_fmap[21][1] = xor_sum[21][1][0];
assign out_fmap[21][2] = xor_sum[21][2][0];
assign out_fmap[21][3] = xor_sum[21][3][0];
assign out_fmap[21][4] = xor_sum[21][4][0];
assign out_fmap[21][5] = xor_sum[21][5][0];
assign out_fmap[21][6] = xor_sum[21][6][0];
assign out_fmap[21][7] = xor_sum[21][7][0];
assign out_fmap[21][8] = xor_sum[21][8][0];
assign out_fmap[21][9] = xor_sum[21][9][0];
assign out_fmap[21][10] = xor_sum[21][10][0];
assign out_fmap[21][11] = xor_sum[21][11][0];
assign out_fmap[21][12] = xor_sum[21][12][0];
assign out_fmap[21][13] = xor_sum[21][13][0];
assign out_fmap[21][14] = xor_sum[21][14][0];
assign out_fmap[21][15] = xor_sum[21][15][0];
assign out_fmap[21][16] = xor_sum[21][16][0];
assign out_fmap[21][17] = xor_sum[21][17][0];
assign out_fmap[21][18] = xor_sum[21][18][0];
assign out_fmap[21][19] = xor_sum[21][19][0];
assign out_fmap[21][20] = xor_sum[21][20][0];
assign out_fmap[21][21] = xor_sum[21][21][0];
assign out_fmap[21][22] = xor_sum[21][22][0];
assign out_fmap[21][23] = xor_sum[21][23][0];
assign out_fmap[22][0] = xor_sum[22][0][0];
assign out_fmap[22][1] = xor_sum[22][1][0];
assign out_fmap[22][2] = xor_sum[22][2][0];
assign out_fmap[22][3] = xor_sum[22][3][0];
assign out_fmap[22][4] = xor_sum[22][4][0];
assign out_fmap[22][5] = xor_sum[22][5][0];
assign out_fmap[22][6] = xor_sum[22][6][0];
assign out_fmap[22][7] = xor_sum[22][7][0];
assign out_fmap[22][8] = xor_sum[22][8][0];
assign out_fmap[22][9] = xor_sum[22][9][0];
assign out_fmap[22][10] = xor_sum[22][10][0];
assign out_fmap[22][11] = xor_sum[22][11][0];
assign out_fmap[22][12] = xor_sum[22][12][0];
assign out_fmap[22][13] = xor_sum[22][13][0];
assign out_fmap[22][14] = xor_sum[22][14][0];
assign out_fmap[22][15] = xor_sum[22][15][0];
assign out_fmap[22][16] = xor_sum[22][16][0];
assign out_fmap[22][17] = xor_sum[22][17][0];
assign out_fmap[22][18] = xor_sum[22][18][0];
assign out_fmap[22][19] = xor_sum[22][19][0];
assign out_fmap[22][20] = xor_sum[22][20][0];
assign out_fmap[22][21] = xor_sum[22][21][0];
assign out_fmap[22][22] = xor_sum[22][22][0];
assign out_fmap[22][23] = xor_sum[22][23][0];
assign out_fmap[23][0] = xor_sum[23][0][0];
assign out_fmap[23][1] = xor_sum[23][1][0];
assign out_fmap[23][2] = xor_sum[23][2][0];
assign out_fmap[23][3] = xor_sum[23][3][0];
assign out_fmap[23][4] = xor_sum[23][4][0];
assign out_fmap[23][5] = xor_sum[23][5][0];
assign out_fmap[23][6] = xor_sum[23][6][0];
assign out_fmap[23][7] = xor_sum[23][7][0];
assign out_fmap[23][8] = xor_sum[23][8][0];
assign out_fmap[23][9] = xor_sum[23][9][0];
assign out_fmap[23][10] = xor_sum[23][10][0];
assign out_fmap[23][11] = xor_sum[23][11][0];
assign out_fmap[23][12] = xor_sum[23][12][0];
assign out_fmap[23][13] = xor_sum[23][13][0];
assign out_fmap[23][14] = xor_sum[23][14][0];
assign out_fmap[23][15] = xor_sum[23][15][0];
assign out_fmap[23][16] = xor_sum[23][16][0];
assign out_fmap[23][17] = xor_sum[23][17][0];
assign out_fmap[23][18] = xor_sum[23][18][0];
assign out_fmap[23][19] = xor_sum[23][19][0];
assign out_fmap[23][20] = xor_sum[23][20][0];
assign out_fmap[23][21] = xor_sum[23][21][0];
assign out_fmap[23][22] = xor_sum[23][22][0];
assign out_fmap[23][23] = xor_sum[23][23][0];

endmodule